/*
  Warren Getlin
  wgetlin@gmail.com

  hazard unit
*/

module hazard_unit(

);