// Copyright (C) 1991-2013 Altera Corporation
// Your use of Altera Corporation's design tools, logic functions 
// and other software and tools, and its AMPP partner logic 
// functions, and any output files from any of the foregoing 
// (including device programming or simulation files), and any 
// associated documentation or information are expressly subject 
// to the terms and conditions of the Altera Program License 
// Subscription Agreement, Altera MegaCore Function License 
// Agreement, or other applicable license agreement, including, 
// without limitation, that your use is for the sole purpose of 
// programming logic devices manufactured by Altera and sold by 
// Altera or its authorized distributors.  Please refer to the 
// applicable agreement for further details.

// VENDOR "Altera"
// PROGRAM "Quartus II 32-bit"
// VERSION "Version 13.0.1 Build 232 06/12/2013 Service Pack 1 SJ Full Version"

// DATE "10/10/2014 15:02:21"

// 
// Device: Altera EP4CE115F29C8 Package FBGA780
// 

// 
// This Verilog file should be used for ModelSim (Verilog) only
// 

`timescale 1 ps/ 1 ps

module system (
	altera_reserved_tms,
	altera_reserved_tck,
	altera_reserved_tdi,
	altera_reserved_tdo,
	CLK,
	nRST,
	\syif.halt ,
	\syif.load ,
	\syif.addr ,
	\syif.store ,
	\syif.REN ,
	\syif.WEN ,
	\syif.tbCTRL );
input 	altera_reserved_tms;
input 	altera_reserved_tck;
input 	altera_reserved_tdi;
output 	altera_reserved_tdo;
input 	CLK;
input 	nRST;
output 	\syif.halt ;
output 	[31:0] \syif.load ;
input 	[31:0] \syif.addr ;
input 	[31:0] \syif.store ;
input 	\syif.REN ;
input 	\syif.WEN ;
input 	\syif.tbCTRL ;

// Design Ports Information
// syif.halt	=>  Location: PIN_AD11,	 I/O Standard: 2.5 V,	 Current Strength: Default
// syif.load[0]	=>  Location: PIN_T3,	 I/O Standard: 2.5 V,	 Current Strength: Default
// syif.load[1]	=>  Location: PIN_AA16,	 I/O Standard: 2.5 V,	 Current Strength: Default
// syif.load[2]	=>  Location: PIN_AC15,	 I/O Standard: 2.5 V,	 Current Strength: Default
// syif.load[3]	=>  Location: PIN_AD14,	 I/O Standard: 2.5 V,	 Current Strength: Default
// syif.load[4]	=>  Location: PIN_AA15,	 I/O Standard: 2.5 V,	 Current Strength: Default
// syif.load[5]	=>  Location: PIN_AF15,	 I/O Standard: 2.5 V,	 Current Strength: Default
// syif.load[6]	=>  Location: PIN_AC14,	 I/O Standard: 2.5 V,	 Current Strength: Default
// syif.load[7]	=>  Location: PIN_U2,	 I/O Standard: 2.5 V,	 Current Strength: Default
// syif.load[8]	=>  Location: PIN_R5,	 I/O Standard: 2.5 V,	 Current Strength: Default
// syif.load[9]	=>  Location: PIN_AB16,	 I/O Standard: 2.5 V,	 Current Strength: Default
// syif.load[10]	=>  Location: PIN_H15,	 I/O Standard: 2.5 V,	 Current Strength: Default
// syif.load[11]	=>  Location: PIN_AD15,	 I/O Standard: 2.5 V,	 Current Strength: Default
// syif.load[12]	=>  Location: PIN_Y15,	 I/O Standard: 2.5 V,	 Current Strength: Default
// syif.load[13]	=>  Location: PIN_AB13,	 I/O Standard: 2.5 V,	 Current Strength: Default
// syif.load[14]	=>  Location: PIN_AH17,	 I/O Standard: 2.5 V,	 Current Strength: Default
// syif.load[15]	=>  Location: PIN_D16,	 I/O Standard: 2.5 V,	 Current Strength: Default
// syif.load[16]	=>  Location: PIN_R1,	 I/O Standard: 2.5 V,	 Current Strength: Default
// syif.load[17]	=>  Location: PIN_AH18,	 I/O Standard: 2.5 V,	 Current Strength: Default
// syif.load[18]	=>  Location: PIN_C16,	 I/O Standard: 2.5 V,	 Current Strength: Default
// syif.load[19]	=>  Location: PIN_H16,	 I/O Standard: 2.5 V,	 Current Strength: Default
// syif.load[20]	=>  Location: PIN_AE16,	 I/O Standard: 2.5 V,	 Current Strength: Default
// syif.load[21]	=>  Location: PIN_E15,	 I/O Standard: 2.5 V,	 Current Strength: Default
// syif.load[22]	=>  Location: PIN_AH19,	 I/O Standard: 2.5 V,	 Current Strength: Default
// syif.load[23]	=>  Location: PIN_AB15,	 I/O Standard: 2.5 V,	 Current Strength: Default
// syif.load[24]	=>  Location: PIN_J15,	 I/O Standard: 2.5 V,	 Current Strength: Default
// syif.load[25]	=>  Location: PIN_R24,	 I/O Standard: 2.5 V,	 Current Strength: Default
// syif.load[26]	=>  Location: PIN_C15,	 I/O Standard: 2.5 V,	 Current Strength: Default
// syif.load[27]	=>  Location: PIN_AC17,	 I/O Standard: 2.5 V,	 Current Strength: Default
// syif.load[28]	=>  Location: PIN_AF16,	 I/O Standard: 2.5 V,	 Current Strength: Default
// syif.load[29]	=>  Location: PIN_AE15,	 I/O Standard: 2.5 V,	 Current Strength: Default
// syif.load[30]	=>  Location: PIN_AG17,	 I/O Standard: 2.5 V,	 Current Strength: Default
// syif.load[31]	=>  Location: PIN_T7,	 I/O Standard: 2.5 V,	 Current Strength: Default
// syif.tbCTRL	=>  Location: PIN_AG15,	 I/O Standard: 2.5 V,	 Current Strength: Default
// syif.addr[1]	=>  Location: PIN_AH15,	 I/O Standard: 2.5 V,	 Current Strength: Default
// syif.addr[0]	=>  Location: PIN_J13,	 I/O Standard: 2.5 V,	 Current Strength: Default
// syif.addr[3]	=>  Location: PIN_AF13,	 I/O Standard: 2.5 V,	 Current Strength: Default
// syif.addr[2]	=>  Location: PIN_H14,	 I/O Standard: 2.5 V,	 Current Strength: Default
// syif.addr[5]	=>  Location: PIN_AC11,	 I/O Standard: 2.5 V,	 Current Strength: Default
// syif.addr[4]	=>  Location: PIN_AG11,	 I/O Standard: 2.5 V,	 Current Strength: Default
// syif.addr[7]	=>  Location: PIN_R23,	 I/O Standard: 2.5 V,	 Current Strength: Default
// syif.addr[6]	=>  Location: PIN_D12,	 I/O Standard: 2.5 V,	 Current Strength: Default
// syif.addr[9]	=>  Location: PIN_T4,	 I/O Standard: 2.5 V,	 Current Strength: Default
// syif.addr[8]	=>  Location: PIN_AD12,	 I/O Standard: 2.5 V,	 Current Strength: Default
// syif.addr[11]	=>  Location: PIN_C13,	 I/O Standard: 2.5 V,	 Current Strength: Default
// syif.addr[10]	=>  Location: PIN_P21,	 I/O Standard: 2.5 V,	 Current Strength: Default
// syif.addr[13]	=>  Location: PIN_T21,	 I/O Standard: 2.5 V,	 Current Strength: Default
// syif.addr[12]	=>  Location: PIN_G14,	 I/O Standard: 2.5 V,	 Current Strength: Default
// syif.addr[15]	=>  Location: PIN_AA12,	 I/O Standard: 2.5 V,	 Current Strength: Default
// syif.addr[14]	=>  Location: PIN_J12,	 I/O Standard: 2.5 V,	 Current Strength: Default
// syif.addr[17]	=>  Location: PIN_AE14,	 I/O Standard: 2.5 V,	 Current Strength: Default
// syif.addr[16]	=>  Location: PIN_AE13,	 I/O Standard: 2.5 V,	 Current Strength: Default
// syif.addr[19]	=>  Location: PIN_AG12,	 I/O Standard: 2.5 V,	 Current Strength: Default
// syif.addr[18]	=>  Location: PIN_AG21,	 I/O Standard: 2.5 V,	 Current Strength: Default
// syif.addr[21]	=>  Location: PIN_C12,	 I/O Standard: 2.5 V,	 Current Strength: Default
// syif.addr[20]	=>  Location: PIN_B11,	 I/O Standard: 2.5 V,	 Current Strength: Default
// syif.addr[23]	=>  Location: PIN_E14,	 I/O Standard: 2.5 V,	 Current Strength: Default
// syif.addr[22]	=>  Location: PIN_C14,	 I/O Standard: 2.5 V,	 Current Strength: Default
// syif.addr[25]	=>  Location: PIN_AB12,	 I/O Standard: 2.5 V,	 Current Strength: Default
// syif.addr[24]	=>  Location: PIN_A12,	 I/O Standard: 2.5 V,	 Current Strength: Default
// syif.addr[27]	=>  Location: PIN_R27,	 I/O Standard: 2.5 V,	 Current Strength: Default
// syif.addr[26]	=>  Location: PIN_AF14,	 I/O Standard: 2.5 V,	 Current Strength: Default
// syif.addr[29]	=>  Location: PIN_U4,	 I/O Standard: 2.5 V,	 Current Strength: Default
// syif.addr[28]	=>  Location: PIN_F14,	 I/O Standard: 2.5 V,	 Current Strength: Default
// syif.addr[31]	=>  Location: PIN_D14,	 I/O Standard: 2.5 V,	 Current Strength: Default
// syif.addr[30]	=>  Location: PIN_J14,	 I/O Standard: 2.5 V,	 Current Strength: Default
// syif.WEN	=>  Location: PIN_R3,	 I/O Standard: 2.5 V,	 Current Strength: Default
// syif.REN	=>  Location: PIN_R28,	 I/O Standard: 2.5 V,	 Current Strength: Default
// nRST	=>  Location: PIN_Y2,	 I/O Standard: 2.5 V,	 Current Strength: Default
// CLK	=>  Location: PIN_J1,	 I/O Standard: 2.5 V,	 Current Strength: Default
// syif.store[0]	=>  Location: PIN_F17,	 I/O Standard: 2.5 V,	 Current Strength: Default
// syif.store[1]	=>  Location: PIN_AA14,	 I/O Standard: 2.5 V,	 Current Strength: Default
// syif.store[2]	=>  Location: PIN_B17,	 I/O Standard: 2.5 V,	 Current Strength: Default
// syif.store[3]	=>  Location: PIN_AA13,	 I/O Standard: 2.5 V,	 Current Strength: Default
// syif.store[4]	=>  Location: PIN_R6,	 I/O Standard: 2.5 V,	 Current Strength: Default
// syif.store[5]	=>  Location: PIN_G16,	 I/O Standard: 2.5 V,	 Current Strength: Default
// syif.store[6]	=>  Location: PIN_AB14,	 I/O Standard: 2.5 V,	 Current Strength: Default
// syif.store[7]	=>  Location: PIN_D15,	 I/O Standard: 2.5 V,	 Current Strength: Default
// syif.store[8]	=>  Location: PIN_U3,	 I/O Standard: 2.5 V,	 Current Strength: Default
// syif.store[9]	=>  Location: PIN_G18,	 I/O Standard: 2.5 V,	 Current Strength: Default
// syif.store[10]	=>  Location: PIN_Y12,	 I/O Standard: 2.5 V,	 Current Strength: Default
// syif.store[11]	=>  Location: PIN_AG19,	 I/O Standard: 2.5 V,	 Current Strength: Default
// syif.store[12]	=>  Location: PIN_F15,	 I/O Standard: 2.5 V,	 Current Strength: Default
// syif.store[13]	=>  Location: PIN_M23,	 I/O Standard: 2.5 V,	 Current Strength: Default
// syif.store[14]	=>  Location: PIN_D13,	 I/O Standard: 2.5 V,	 Current Strength: Default
// syif.store[15]	=>  Location: PIN_R7,	 I/O Standard: 2.5 V,	 Current Strength: Default
// syif.store[16]	=>  Location: PIN_U1,	 I/O Standard: 2.5 V,	 Current Strength: Default
// syif.store[17]	=>  Location: PIN_H17,	 I/O Standard: 2.5 V,	 Current Strength: Default
// syif.store[18]	=>  Location: PIN_Y14,	 I/O Standard: 2.5 V,	 Current Strength: Default
// syif.store[19]	=>  Location: PIN_AE17,	 I/O Standard: 2.5 V,	 Current Strength: Default
// syif.store[20]	=>  Location: PIN_B10,	 I/O Standard: 2.5 V,	 Current Strength: Default
// syif.store[21]	=>  Location: PIN_T22,	 I/O Standard: 2.5 V,	 Current Strength: Default
// syif.store[22]	=>  Location: PIN_A17,	 I/O Standard: 2.5 V,	 Current Strength: Default
// syif.store[23]	=>  Location: PIN_Y13,	 I/O Standard: 2.5 V,	 Current Strength: Default
// syif.store[24]	=>  Location: PIN_V4,	 I/O Standard: 2.5 V,	 Current Strength: Default
// syif.store[25]	=>  Location: PIN_AH12,	 I/O Standard: 2.5 V,	 Current Strength: Default
// syif.store[26]	=>  Location: PIN_AC12,	 I/O Standard: 2.5 V,	 Current Strength: Default
// syif.store[27]	=>  Location: PIN_A11,	 I/O Standard: 2.5 V,	 Current Strength: Default
// syif.store[28]	=>  Location: PIN_G15,	 I/O Standard: 2.5 V,	 Current Strength: Default
// syif.store[29]	=>  Location: PIN_J16,	 I/O Standard: 2.5 V,	 Current Strength: Default
// syif.store[30]	=>  Location: PIN_AG18,	 I/O Standard: 2.5 V,	 Current Strength: Default
// syif.store[31]	=>  Location: PIN_AF17,	 I/O Standard: 2.5 V,	 Current Strength: Default
// altera_reserved_tms	=>  Location: PIN_P8,	 I/O Standard: 2.5 V,	 Current Strength: Default
// altera_reserved_tck	=>  Location: PIN_P5,	 I/O Standard: 2.5 V,	 Current Strength: Default
// altera_reserved_tdi	=>  Location: PIN_P7,	 I/O Standard: 2.5 V,	 Current Strength: Default
// altera_reserved_tdo	=>  Location: PIN_P6,	 I/O Standard: 2.5 V,	 Current Strength: Default


wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
assign unknown = 1'bx;

tri1 devclrn;
tri1 devpor;
tri1 devoe;
// synopsys translate_off
initial $sdf_annotate("mapped/system_v.sdo");
// synopsys translate_on

wire \RAM|altsyncram_component|auto_generated|mgl_prim2|is_in_use_reg~q ;
wire \CPU|DP|EXMEM|plif_exmem.hlt_l~q ;
wire \CPU|DP|EXMEM|plif_exmem.dmemWEN_l~q ;
wire \CPU|DP|EXMEM|plif_exmem.dmemREN_l~q ;
wire \ramaddr~0_combout ;
wire \ramaddr~1_combout ;
wire \ramaddr~2_combout ;
wire \ramaddr~3_combout ;
wire \ramaddr~4_combout ;
wire \ramaddr~5_combout ;
wire \ramaddr~6_combout ;
wire \ramaddr~7_combout ;
wire \ramaddr~8_combout ;
wire \ramaddr~9_combout ;
wire \ramaddr~10_combout ;
wire \ramaddr~11_combout ;
wire \ramaddr~12_combout ;
wire \ramaddr~13_combout ;
wire \ramaddr~14_combout ;
wire \ramaddr~15_combout ;
wire \ramaddr~16_combout ;
wire \ramaddr~17_combout ;
wire \ramaddr~18_combout ;
wire \ramaddr~19_combout ;
wire \ramaddr~20_combout ;
wire \ramaddr~21_combout ;
wire \ramaddr~22_combout ;
wire \ramaddr~23_combout ;
wire \ramaddr~24_combout ;
wire \ramaddr~25_combout ;
wire \ramaddr~26_combout ;
wire \ramaddr~27_combout ;
wire \ramaddr~28_combout ;
wire \ramaddr~29_combout ;
wire \ramaddr~30_combout ;
wire \ramaddr~31_combout ;
wire \ramaddr~32_combout ;
wire \ramaddr~33_combout ;
wire \ramaddr~34_combout ;
wire \ramaddr~35_combout ;
wire \ramaddr~36_combout ;
wire \ramaddr~37_combout ;
wire \ramaddr~38_combout ;
wire \ramaddr~39_combout ;
wire \ramaddr~40_combout ;
wire \ramaddr~41_combout ;
wire \ramaddr~42_combout ;
wire \ramaddr~43_combout ;
wire \ramaddr~44_combout ;
wire \ramaddr~45_combout ;
wire \ramaddr~46_combout ;
wire \ramaddr~47_combout ;
wire \ramaddr~48_combout ;
wire \ramaddr~49_combout ;
wire \ramaddr~50_combout ;
wire \ramaddr~51_combout ;
wire \ramaddr~52_combout ;
wire \ramaddr~53_combout ;
wire \ramaddr~54_combout ;
wire \ramaddr~55_combout ;
wire \ramaddr~56_combout ;
wire \ramaddr~57_combout ;
wire \ramaddr~58_combout ;
wire \ramaddr~59_combout ;
wire \ramaddr~60_combout ;
wire \ramaddr~61_combout ;
wire \ramWEN~0_combout ;
wire \CPU|DP|dpif.imemREN~q ;
wire \ramREN~0_combout ;
wire \ramREN~1_combout ;
wire \RAM|always1~0_combout ;
wire \RAM|ramif.ramload[0]~0_combout ;
wire \RAM|ramif.ramload[1]~1_combout ;
wire \RAM|ramif.ramload[2]~2_combout ;
wire \RAM|ramif.ramload[3]~3_combout ;
wire \RAM|ramif.ramload[4]~4_combout ;
wire \RAM|ramif.ramload[5]~5_combout ;
wire \RAM|ramif.ramload[6]~6_combout ;
wire \RAM|ramif.ramload[7]~7_combout ;
wire \RAM|ramif.ramload[8]~8_combout ;
wire \RAM|ramif.ramload[9]~9_combout ;
wire \RAM|ramif.ramload[10]~10_combout ;
wire \RAM|ramif.ramload[11]~11_combout ;
wire \RAM|ramif.ramload[12]~12_combout ;
wire \RAM|ramif.ramload[13]~13_combout ;
wire \RAM|ramif.ramload[14]~14_combout ;
wire \RAM|ramif.ramload[15]~15_combout ;
wire \RAM|ramif.ramload[16]~16_combout ;
wire \RAM|ramif.ramload[17]~17_combout ;
wire \RAM|ramif.ramload[18]~18_combout ;
wire \RAM|ramif.ramload[19]~19_combout ;
wire \RAM|ramif.ramload[20]~20_combout ;
wire \RAM|ramif.ramload[21]~21_combout ;
wire \RAM|ramif.ramload[22]~22_combout ;
wire \RAM|ramif.ramload[23]~23_combout ;
wire \RAM|ramif.ramload[24]~24_combout ;
wire \RAM|ramif.ramload[25]~25_combout ;
wire \RAM|ramif.ramload[26]~26_combout ;
wire \RAM|ramif.ramload[27]~27_combout ;
wire \RAM|ramif.ramload[28]~28_combout ;
wire \RAM|ramif.ramload[29]~29_combout ;
wire \RAM|ramif.ramload[30]~30_combout ;
wire \RAM|ramif.ramload[31]~31_combout ;
wire \RAM|altsyncram_component|auto_generated|mgl_prim2|tdo~1_combout ;
wire \CPUCLK~q ;
wire \ramstore~0_combout ;
wire \ramaddr~62_combout ;
wire \ramaddr~63_combout ;
wire \ramstore~1_combout ;
wire \ramstore~2_combout ;
wire \ramstore~3_combout ;
wire \ramstore~4_combout ;
wire \ramstore~5_combout ;
wire \ramstore~6_combout ;
wire \ramstore~7_combout ;
wire \ramstore~8_combout ;
wire \ramstore~9_combout ;
wire \ramstore~10_combout ;
wire \ramstore~11_combout ;
wire \ramstore~12_combout ;
wire \ramstore~13_combout ;
wire \ramstore~14_combout ;
wire \ramstore~15_combout ;
wire \ramstore~16_combout ;
wire \ramstore~17_combout ;
wire \ramstore~18_combout ;
wire \ramstore~19_combout ;
wire \ramstore~20_combout ;
wire \ramstore~21_combout ;
wire \ramstore~22_combout ;
wire \ramstore~23_combout ;
wire \ramstore~24_combout ;
wire \ramstore~25_combout ;
wire \ramstore~26_combout ;
wire \ramstore~27_combout ;
wire \ramstore~28_combout ;
wire \ramstore~29_combout ;
wire \ramstore~30_combout ;
wire \ramstore~31_combout ;
wire \Equal0~0_combout ;
wire \CPUCLK~0_combout ;
wire \count[3]~0_combout ;
wire \count[2]~1_combout ;
wire \count[1]~2_combout ;
wire \count~3_combout ;
wire \ramaddr~27_wirecell_combout ;
wire \altera_internal_jtag~TCKUTAP ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter[0]~12 ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter[0]~11_combout ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter[1]~14 ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter[1]~13_combout ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter[2]~16 ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter[2]~15_combout ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter[3]~19 ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter[3]~18_combout ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter[4]~20_combout ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irf_reg[1][0]~q ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irf_reg[1][1]~q ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irf_reg[1][2]~q ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irf_reg[1][3]~q ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irf_reg[1][4]~q ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|node_ena[1]~reg0_q ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|tdo~0_combout ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|reset_ena_reg_proc~0_combout ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irf_reg[1][0]~0_combout ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|node_ena~0_combout ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|node_ena~1_combout ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|node_ena_proc~0_combout ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|node_ena~2_combout ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|node_ena~3_combout ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|Equal0~0_combout ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg[3]~13_combout ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_minor_ver_reg~0_combout ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|WORD_SR~6_combout ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|WORD_SR~7_combout ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|WORD_SR~8_combout ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg~7_combout ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|reset_ena_reg~q ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg~15_combout ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|Equal3~0_combout ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_mode_reg[0]~4_combout ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_minor_ver_reg~1_combout ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter[1]~17_combout ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|WORD_SR~9_combout ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|tms_cnt~2_combout ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg~16_combout ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg~17_combout ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg~18_combout ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_minor_ver_reg~2_combout ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|WORD_SR~10_combout ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|WORD_SR~11_combout ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|WORD_SR~12_combout ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_minor_ver_reg~3_combout ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|WORD_SR~13_combout ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|WORD_SR~14_combout ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|WORD_SR[1]~15_combout ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter[1]~22_combout ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter[1]~23_combout ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|WORD_SR~16_combout ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg~20_combout ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg~21_combout ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg~22_combout ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg~23_combout ;
wire \auto_hub|~GND~combout ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|clr_reg~_wirecell_combout ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state[0]~_wirecell_combout ;
wire \syif.tbCTRL~input_o ;
wire \syif.addr[1]~input_o ;
wire \syif.addr[0]~input_o ;
wire \syif.addr[3]~input_o ;
wire \syif.addr[2]~input_o ;
wire \syif.addr[5]~input_o ;
wire \syif.addr[4]~input_o ;
wire \syif.addr[7]~input_o ;
wire \syif.addr[6]~input_o ;
wire \syif.addr[9]~input_o ;
wire \syif.addr[8]~input_o ;
wire \syif.addr[11]~input_o ;
wire \syif.addr[10]~input_o ;
wire \syif.addr[13]~input_o ;
wire \syif.addr[12]~input_o ;
wire \syif.addr[15]~input_o ;
wire \syif.addr[14]~input_o ;
wire \syif.addr[17]~input_o ;
wire \syif.addr[16]~input_o ;
wire \syif.addr[19]~input_o ;
wire \syif.addr[18]~input_o ;
wire \syif.addr[21]~input_o ;
wire \syif.addr[20]~input_o ;
wire \syif.addr[23]~input_o ;
wire \syif.addr[22]~input_o ;
wire \syif.addr[25]~input_o ;
wire \syif.addr[24]~input_o ;
wire \syif.addr[27]~input_o ;
wire \syif.addr[26]~input_o ;
wire \syif.addr[29]~input_o ;
wire \syif.addr[28]~input_o ;
wire \syif.addr[31]~input_o ;
wire \syif.addr[30]~input_o ;
wire \syif.WEN~input_o ;
wire \syif.REN~input_o ;
wire \nRST~input_o ;
wire \CLK~input_o ;
wire \syif.store[0]~input_o ;
wire \syif.store[1]~input_o ;
wire \syif.store[2]~input_o ;
wire \syif.store[3]~input_o ;
wire \syif.store[4]~input_o ;
wire \syif.store[5]~input_o ;
wire \syif.store[6]~input_o ;
wire \syif.store[7]~input_o ;
wire \syif.store[8]~input_o ;
wire \syif.store[9]~input_o ;
wire \syif.store[10]~input_o ;
wire \syif.store[11]~input_o ;
wire \syif.store[12]~input_o ;
wire \syif.store[13]~input_o ;
wire \syif.store[14]~input_o ;
wire \syif.store[15]~input_o ;
wire \syif.store[16]~input_o ;
wire \syif.store[17]~input_o ;
wire \syif.store[18]~input_o ;
wire \syif.store[19]~input_o ;
wire \syif.store[20]~input_o ;
wire \syif.store[21]~input_o ;
wire \syif.store[22]~input_o ;
wire \syif.store[23]~input_o ;
wire \syif.store[24]~input_o ;
wire \syif.store[25]~input_o ;
wire \syif.store[26]~input_o ;
wire \syif.store[27]~input_o ;
wire \syif.store[28]~input_o ;
wire \syif.store[29]~input_o ;
wire \syif.store[30]~input_o ;
wire \syif.store[31]~input_o ;
wire \altera_internal_jtag~TCKUTAPclkctrl_outclk ;
wire \CPUCLK~clkctrl_outclk ;
wire \nRST~inputclkctrl_outclk ;
wire \CLK~inputclkctrl_outclk ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irf_reg[1][3]~feeder_combout ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irf_reg[1][0]~feeder_combout ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irf_reg[1][2]~feeder_combout ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irf_reg[1][1]~feeder_combout ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|identity_contrib_update_reg[1]~feeder_combout ;
wire \altera_reserved_tms~input_o ;
wire \altera_reserved_tck~input_o ;
wire \altera_reserved_tdi~input_o ;
wire \altera_internal_jtag~TDIUTAP ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg[5]~0_combout ;
wire \~QIC_CREATED_GND~I_combout ;
wire \altera_internal_jtag~TMSUTAP ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state~6_combout ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state~7_combout ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state~4_combout ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state~5_combout ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irf_proc~0_combout ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|tms_cnt~1_combout ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|tms_cnt~0_combout ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state~0_combout ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state~1_combout ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|node_ena_proc~1_combout ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state[9]~feeder_combout ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state~8_combout ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state~11_combout ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state~12_combout ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state~9_combout ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state~10_combout ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|virtual_ir_dr_scan_proc~0_combout ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state~2_combout ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state~3_combout ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg~5_combout ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg[9]~feeder_combout ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg[8]~feeder_combout ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg[7]~feeder_combout ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg[6]~feeder_combout ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg[4]~feeder_combout ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg[3]~feeder_combout ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg[2]~0_combout ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg[1]~feeder_combout ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg[0]~1_combout ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|Equal0~1_combout ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|Equal1~0_combout ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|virtual_ir_scan_reg~q ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg[3]~1_combout ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg~9_combout ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg~8_combout ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg[2]~3_combout ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg[0]~4_combout ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg~6_combout ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg~2_combout ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_mode_reg[1]~0_combout ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_mode_reg[1]~1_combout ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_mode_reg[2]~2_combout ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_mode_reg[2]~3_combout ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|clr_reg_proc~0_combout ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|clr_reg~q ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|tdo_bypass_reg~0_combout ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|tdo_bypass_reg~q ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|tdo~1_combout ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|tdo~2_combout ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg[0]~5_combout ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|clear_signal~combout ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg[2]~9_combout ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|Equal0~2_combout ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|virtual_dr_scan_reg~q ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg[4]~12_combout ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg[3]~13_combout ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg~12_combout ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg[4]~11_combout ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg[0]~6 ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg[1]~7_combout ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg[1]~8 ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg[2]~10 ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg[3]~14 ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg[4]~15_combout ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg[3]~14_combout ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|identity_contrib_shift_reg[3]~feeder_combout ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|identity_contrib_shift_reg[0]~0_combout ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|identity_contrib_shift_reg[0]~1_combout ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|identity_contrib_shift_reg[1]~feeder_combout ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|identity_contrib_shift_reg[0]~feeder_combout ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|identity_contrib_update_reg[0]~feeder_combout ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|identity_contrib_update_reg[0]~0_combout ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg[0]~0_combout ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg~11_combout ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg~10_combout ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg~19_combout ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg[1]~1_combout ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|identity_contrib_update_reg[2]~feeder_combout ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg[2]~2_combout ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg[3]~3_combout ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_proc~0_combout ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg_ena~combout ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|tdo~3_combout ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|tdo~4_combout ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|tdo~5_combout ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg_ena~0_combout ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|tdo~q ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|tdo~_wirecell_combout ;
wire \altera_internal_jtag~TDO ;
wire [4:0] \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg ;
wire [9:0] \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg ;
wire [5:0] \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg ;
wire [3:0] \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|identity_contrib_update_reg ;
wire [3:0] \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|identity_contrib_shift_reg ;
wire [2:0] \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_mode_reg ;
wire [3:0] \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_minor_ver_reg ;
wire [3:0] \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg ;
wire [2:0] \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|tms_cnt ;
wire [15:0] \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state ;
wire [4:0] \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter ;
wire [3:0] \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|WORD_SR ;
wire [3:0] count;
wire [31:0] \CPU|DP|PC|PCreg ;
wire [3:0] \RAM|altsyncram_component|auto_generated|mgl_prim2|ir_loaded_address_reg ;
wire [31:0] \CPU|DP|EXMEM|plif_exmem.rdat2_l ;
wire [31:0] \CPU|DP|EXMEM|plif_exmem.porto_l ;


ram RAM(
	.is_in_use_reg(\RAM|altsyncram_component|auto_generated|mgl_prim2|is_in_use_reg~q ),
	.ramaddr(\ramaddr~0_combout ),
	.ramaddr1(\ramaddr~1_combout ),
	.ramaddr2(\ramaddr~3_combout ),
	.ramaddr3(\ramaddr~5_combout ),
	.ramaddr4(\ramaddr~7_combout ),
	.ramaddr5(\ramaddr~9_combout ),
	.ramaddr6(\ramaddr~11_combout ),
	.ramaddr7(\ramaddr~13_combout ),
	.ramaddr8(\ramaddr~15_combout ),
	.ramaddr9(\ramaddr~17_combout ),
	.ramaddr10(\ramaddr~19_combout ),
	.ramaddr11(\ramaddr~21_combout ),
	.ramaddr12(\ramaddr~23_combout ),
	.ramaddr13(\ramaddr~25_combout ),
	.ramaddr14(\ramaddr~27_combout ),
	.ramaddr15(\ramaddr~29_combout ),
	.\ramif.ramaddr ({\ramaddr~59_combout ,\ramaddr~61_combout ,\ramaddr~55_combout ,gnd,\ramaddr~51_combout ,\ramaddr~53_combout ,gnd,gnd,\ramaddr~43_combout ,\ramaddr~45_combout ,\ramaddr~39_combout ,\ramaddr~41_combout ,\ramaddr~35_combout ,gnd,\ramaddr~31_combout ,\ramaddr~33_combout ,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,\ramaddr~62_combout ,\ramaddr~63_combout }),
	.ramaddr16(\ramaddr~37_combout ),
	.ramaddr17(\ramaddr~47_combout ),
	.ramaddr18(\ramaddr~49_combout ),
	.ramaddr19(\ramaddr~57_combout ),
	.\ramif.ramWEN (\ramWEN~0_combout ),
	.\ramif.ramREN (\ramREN~1_combout ),
	.always1(\RAM|always1~0_combout ),
	.ramiframload_0(\RAM|ramif.ramload[0]~0_combout ),
	.ramiframload_1(\RAM|ramif.ramload[1]~1_combout ),
	.ramiframload_2(\RAM|ramif.ramload[2]~2_combout ),
	.ramiframload_3(\RAM|ramif.ramload[3]~3_combout ),
	.ramiframload_4(\RAM|ramif.ramload[4]~4_combout ),
	.ramiframload_5(\RAM|ramif.ramload[5]~5_combout ),
	.ramiframload_6(\RAM|ramif.ramload[6]~6_combout ),
	.ramiframload_7(\RAM|ramif.ramload[7]~7_combout ),
	.ramiframload_8(\RAM|ramif.ramload[8]~8_combout ),
	.ramiframload_9(\RAM|ramif.ramload[9]~9_combout ),
	.ramiframload_10(\RAM|ramif.ramload[10]~10_combout ),
	.ramiframload_11(\RAM|ramif.ramload[11]~11_combout ),
	.ramiframload_12(\RAM|ramif.ramload[12]~12_combout ),
	.ramiframload_13(\RAM|ramif.ramload[13]~13_combout ),
	.ramiframload_14(\RAM|ramif.ramload[14]~14_combout ),
	.ramiframload_15(\RAM|ramif.ramload[15]~15_combout ),
	.ramiframload_16(\RAM|ramif.ramload[16]~16_combout ),
	.ramiframload_17(\RAM|ramif.ramload[17]~17_combout ),
	.ramiframload_18(\RAM|ramif.ramload[18]~18_combout ),
	.ramiframload_19(\RAM|ramif.ramload[19]~19_combout ),
	.ramiframload_20(\RAM|ramif.ramload[20]~20_combout ),
	.ramiframload_21(\RAM|ramif.ramload[21]~21_combout ),
	.ramiframload_22(\RAM|ramif.ramload[22]~22_combout ),
	.ramiframload_23(\RAM|ramif.ramload[23]~23_combout ),
	.ramiframload_24(\RAM|ramif.ramload[24]~24_combout ),
	.ramiframload_25(\RAM|ramif.ramload[25]~25_combout ),
	.ramiframload_26(\RAM|ramif.ramload[26]~26_combout ),
	.ramiframload_27(\RAM|ramif.ramload[27]~27_combout ),
	.ramiframload_28(\RAM|ramif.ramload[28]~28_combout ),
	.ramiframload_29(\RAM|ramif.ramload[29]~29_combout ),
	.ramiframload_30(\RAM|ramif.ramload[30]~30_combout ),
	.ramiframload_31(\RAM|ramif.ramload[31]~31_combout ),
	.ir_loaded_address_reg_0(\RAM|altsyncram_component|auto_generated|mgl_prim2|ir_loaded_address_reg [0]),
	.ir_loaded_address_reg_1(\RAM|altsyncram_component|auto_generated|mgl_prim2|ir_loaded_address_reg [1]),
	.ir_loaded_address_reg_2(\RAM|altsyncram_component|auto_generated|mgl_prim2|ir_loaded_address_reg [2]),
	.ir_loaded_address_reg_3(\RAM|altsyncram_component|auto_generated|mgl_prim2|ir_loaded_address_reg [3]),
	.tdo(\RAM|altsyncram_component|auto_generated|mgl_prim2|tdo~1_combout ),
	.ramstore(\ramstore~0_combout ),
	.ramstore1(\ramstore~1_combout ),
	.ramstore2(\ramstore~2_combout ),
	.ramstore3(\ramstore~3_combout ),
	.ramstore4(\ramstore~4_combout ),
	.ramstore5(\ramstore~5_combout ),
	.ramstore6(\ramstore~6_combout ),
	.ramstore7(\ramstore~7_combout ),
	.ramstore8(\ramstore~8_combout ),
	.ramstore9(\ramstore~9_combout ),
	.ramstore10(\ramstore~10_combout ),
	.ramstore11(\ramstore~11_combout ),
	.ramstore12(\ramstore~12_combout ),
	.ramstore13(\ramstore~13_combout ),
	.ramstore14(\ramstore~14_combout ),
	.ramstore15(\ramstore~15_combout ),
	.ramstore16(\ramstore~16_combout ),
	.ramstore17(\ramstore~17_combout ),
	.ramstore18(\ramstore~18_combout ),
	.ramstore19(\ramstore~19_combout ),
	.ramstore20(\ramstore~20_combout ),
	.ramstore21(\ramstore~21_combout ),
	.ramstore22(\ramstore~22_combout ),
	.ramstore23(\ramstore~23_combout ),
	.ramstore24(\ramstore~24_combout ),
	.ramstore25(\ramstore~25_combout ),
	.ramstore26(\ramstore~26_combout ),
	.ramstore27(\ramstore~27_combout ),
	.ramstore28(\ramstore~28_combout ),
	.ramstore29(\ramstore~29_combout ),
	.ramstore30(\ramstore~30_combout ),
	.ramstore31(\ramstore~31_combout ),
	.ramaddr20(\ramaddr~27_wirecell_combout ),
	.altera_internal_jtag(\altera_internal_jtag~TDIUTAP ),
	.state_4(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [4]),
	.irf_reg_0_1(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irf_reg[1][0]~q ),
	.irf_reg_1_1(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irf_reg[1][1]~q ),
	.irf_reg_2_1(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irf_reg[1][2]~q ),
	.irf_reg_3_1(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irf_reg[1][3]~q ),
	.irf_reg_4_1(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irf_reg[1][4]~q ),
	.node_ena_1(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|node_ena[1]~reg0_q ),
	.clr_reg(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|clr_reg~q ),
	.virtual_ir_scan_reg(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|virtual_ir_scan_reg~q ),
	.state_3(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [3]),
	.state_5(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [5]),
	.state_8(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [8]),
	.syiftbCTRL(\syif.tbCTRL~input_o ),
	.syifaddr_1(\syif.addr[1]~input_o ),
	.syifaddr_0(\syif.addr[0]~input_o ),
	.nRST(\nRST~input_o ),
	.altera_internal_jtag1(\altera_internal_jtag~TCKUTAPclkctrl_outclk ),
	.nRST1(\nRST~inputclkctrl_outclk ),
	.CLK(\CLK~inputclkctrl_outclk ),
	.devpor(devpor),
	.devclrn(devclrn),
	.devoe(devoe));

pipeline CPU(
	.PCreg_1(\CPU|DP|PC|PCreg [1]),
	.PCreg_0(\CPU|DP|PC|PCreg [0]),
	.plif_exmemhlt_l(\CPU|DP|EXMEM|plif_exmem.hlt_l~q ),
	.plif_exmemporto_l_1(\CPU|DP|EXMEM|plif_exmem.porto_l [1]),
	.plif_exmemdmemWEN_l(\CPU|DP|EXMEM|plif_exmem.dmemWEN_l~q ),
	.plif_exmemdmemREN_l(\CPU|DP|EXMEM|plif_exmem.dmemREN_l~q ),
	.plif_exmemporto_l_0(\CPU|DP|EXMEM|plif_exmem.porto_l [0]),
	.plif_exmemporto_l_3(\CPU|DP|EXMEM|plif_exmem.porto_l [3]),
	.PCreg_3(\CPU|DP|PC|PCreg [3]),
	.plif_exmemporto_l_2(\CPU|DP|EXMEM|plif_exmem.porto_l [2]),
	.PCreg_2(\CPU|DP|PC|PCreg [2]),
	.plif_exmemporto_l_5(\CPU|DP|EXMEM|plif_exmem.porto_l [5]),
	.PCreg_5(\CPU|DP|PC|PCreg [5]),
	.plif_exmemporto_l_4(\CPU|DP|EXMEM|plif_exmem.porto_l [4]),
	.PCreg_4(\CPU|DP|PC|PCreg [4]),
	.plif_exmemporto_l_7(\CPU|DP|EXMEM|plif_exmem.porto_l [7]),
	.PCreg_7(\CPU|DP|PC|PCreg [7]),
	.plif_exmemporto_l_6(\CPU|DP|EXMEM|plif_exmem.porto_l [6]),
	.PCreg_6(\CPU|DP|PC|PCreg [6]),
	.plif_exmemporto_l_9(\CPU|DP|EXMEM|plif_exmem.porto_l [9]),
	.PCreg_9(\CPU|DP|PC|PCreg [9]),
	.plif_exmemporto_l_8(\CPU|DP|EXMEM|plif_exmem.porto_l [8]),
	.PCreg_8(\CPU|DP|PC|PCreg [8]),
	.plif_exmemporto_l_11(\CPU|DP|EXMEM|plif_exmem.porto_l [11]),
	.PCreg_11(\CPU|DP|PC|PCreg [11]),
	.plif_exmemporto_l_10(\CPU|DP|EXMEM|plif_exmem.porto_l [10]),
	.PCreg_10(\CPU|DP|PC|PCreg [10]),
	.plif_exmemporto_l_13(\CPU|DP|EXMEM|plif_exmem.porto_l [13]),
	.PCreg_13(\CPU|DP|PC|PCreg [13]),
	.plif_exmemporto_l_12(\CPU|DP|EXMEM|plif_exmem.porto_l [12]),
	.PCreg_12(\CPU|DP|PC|PCreg [12]),
	.plif_exmemporto_l_15(\CPU|DP|EXMEM|plif_exmem.porto_l [15]),
	.PCreg_15(\CPU|DP|PC|PCreg [15]),
	.plif_exmemporto_l_14(\CPU|DP|EXMEM|plif_exmem.porto_l [14]),
	.PCreg_14(\CPU|DP|PC|PCreg [14]),
	.plif_exmemporto_l_17(\CPU|DP|EXMEM|plif_exmem.porto_l [17]),
	.PCreg_17(\CPU|DP|PC|PCreg [17]),
	.plif_exmemporto_l_16(\CPU|DP|EXMEM|plif_exmem.porto_l [16]),
	.PCreg_16(\CPU|DP|PC|PCreg [16]),
	.plif_exmemporto_l_19(\CPU|DP|EXMEM|plif_exmem.porto_l [19]),
	.PCreg_19(\CPU|DP|PC|PCreg [19]),
	.plif_exmemporto_l_18(\CPU|DP|EXMEM|plif_exmem.porto_l [18]),
	.PCreg_18(\CPU|DP|PC|PCreg [18]),
	.plif_exmemporto_l_21(\CPU|DP|EXMEM|plif_exmem.porto_l [21]),
	.PCreg_21(\CPU|DP|PC|PCreg [21]),
	.plif_exmemporto_l_20(\CPU|DP|EXMEM|plif_exmem.porto_l [20]),
	.PCreg_20(\CPU|DP|PC|PCreg [20]),
	.plif_exmemporto_l_23(\CPU|DP|EXMEM|plif_exmem.porto_l [23]),
	.PCreg_23(\CPU|DP|PC|PCreg [23]),
	.plif_exmemporto_l_22(\CPU|DP|EXMEM|plif_exmem.porto_l [22]),
	.PCreg_22(\CPU|DP|PC|PCreg [22]),
	.plif_exmemporto_l_25(\CPU|DP|EXMEM|plif_exmem.porto_l [25]),
	.PCreg_25(\CPU|DP|PC|PCreg [25]),
	.plif_exmemporto_l_24(\CPU|DP|EXMEM|plif_exmem.porto_l [24]),
	.PCreg_24(\CPU|DP|PC|PCreg [24]),
	.plif_exmemporto_l_27(\CPU|DP|EXMEM|plif_exmem.porto_l [27]),
	.PCreg_27(\CPU|DP|PC|PCreg [27]),
	.plif_exmemporto_l_26(\CPU|DP|EXMEM|plif_exmem.porto_l [26]),
	.PCreg_26(\CPU|DP|PC|PCreg [26]),
	.plif_exmemporto_l_29(\CPU|DP|EXMEM|plif_exmem.porto_l [29]),
	.PCreg_29(\CPU|DP|PC|PCreg [29]),
	.plif_exmemporto_l_28(\CPU|DP|EXMEM|plif_exmem.porto_l [28]),
	.PCreg_28(\CPU|DP|PC|PCreg [28]),
	.plif_exmemporto_l_31(\CPU|DP|EXMEM|plif_exmem.porto_l [31]),
	.PCreg_31(\CPU|DP|PC|PCreg [31]),
	.plif_exmemporto_l_30(\CPU|DP|EXMEM|plif_exmem.porto_l [30]),
	.PCreg_30(\CPU|DP|PC|PCreg [30]),
	.dpifimemREN(\CPU|DP|dpif.imemREN~q ),
	.always1(\RAM|always1~0_combout ),
	.ramiframload_0(\RAM|ramif.ramload[0]~0_combout ),
	.ramiframload_1(\RAM|ramif.ramload[1]~1_combout ),
	.ramiframload_2(\RAM|ramif.ramload[2]~2_combout ),
	.ramiframload_3(\RAM|ramif.ramload[3]~3_combout ),
	.ramiframload_4(\RAM|ramif.ramload[4]~4_combout ),
	.ramiframload_5(\RAM|ramif.ramload[5]~5_combout ),
	.ramiframload_6(\RAM|ramif.ramload[6]~6_combout ),
	.ramiframload_7(\RAM|ramif.ramload[7]~7_combout ),
	.ramiframload_8(\RAM|ramif.ramload[8]~8_combout ),
	.ramiframload_9(\RAM|ramif.ramload[9]~9_combout ),
	.ramiframload_10(\RAM|ramif.ramload[10]~10_combout ),
	.ramiframload_11(\RAM|ramif.ramload[11]~11_combout ),
	.ramiframload_12(\RAM|ramif.ramload[12]~12_combout ),
	.ramiframload_13(\RAM|ramif.ramload[13]~13_combout ),
	.ramiframload_14(\RAM|ramif.ramload[14]~14_combout ),
	.ramiframload_15(\RAM|ramif.ramload[15]~15_combout ),
	.ramiframload_16(\RAM|ramif.ramload[16]~16_combout ),
	.ramiframload_17(\RAM|ramif.ramload[17]~17_combout ),
	.ramiframload_18(\RAM|ramif.ramload[18]~18_combout ),
	.ramiframload_19(\RAM|ramif.ramload[19]~19_combout ),
	.ramiframload_20(\RAM|ramif.ramload[20]~20_combout ),
	.ramiframload_21(\RAM|ramif.ramload[21]~21_combout ),
	.ramiframload_22(\RAM|ramif.ramload[22]~22_combout ),
	.ramiframload_23(\RAM|ramif.ramload[23]~23_combout ),
	.ramiframload_24(\RAM|ramif.ramload[24]~24_combout ),
	.ramiframload_25(\RAM|ramif.ramload[25]~25_combout ),
	.ramiframload_26(\RAM|ramif.ramload[26]~26_combout ),
	.ramiframload_27(\RAM|ramif.ramload[27]~27_combout ),
	.ramiframload_28(\RAM|ramif.ramload[28]~28_combout ),
	.ramiframload_29(\RAM|ramif.ramload[29]~29_combout ),
	.ramiframload_30(\RAM|ramif.ramload[30]~30_combout ),
	.ramiframload_31(\RAM|ramif.ramload[31]~31_combout ),
	.plif_exmemrdat2_l_0(\CPU|DP|EXMEM|plif_exmem.rdat2_l [0]),
	.plif_exmemrdat2_l_1(\CPU|DP|EXMEM|plif_exmem.rdat2_l [1]),
	.plif_exmemrdat2_l_2(\CPU|DP|EXMEM|plif_exmem.rdat2_l [2]),
	.plif_exmemrdat2_l_3(\CPU|DP|EXMEM|plif_exmem.rdat2_l [3]),
	.plif_exmemrdat2_l_4(\CPU|DP|EXMEM|plif_exmem.rdat2_l [4]),
	.plif_exmemrdat2_l_5(\CPU|DP|EXMEM|plif_exmem.rdat2_l [5]),
	.plif_exmemrdat2_l_6(\CPU|DP|EXMEM|plif_exmem.rdat2_l [6]),
	.plif_exmemrdat2_l_7(\CPU|DP|EXMEM|plif_exmem.rdat2_l [7]),
	.plif_exmemrdat2_l_8(\CPU|DP|EXMEM|plif_exmem.rdat2_l [8]),
	.plif_exmemrdat2_l_9(\CPU|DP|EXMEM|plif_exmem.rdat2_l [9]),
	.plif_exmemrdat2_l_10(\CPU|DP|EXMEM|plif_exmem.rdat2_l [10]),
	.plif_exmemrdat2_l_11(\CPU|DP|EXMEM|plif_exmem.rdat2_l [11]),
	.plif_exmemrdat2_l_12(\CPU|DP|EXMEM|plif_exmem.rdat2_l [12]),
	.plif_exmemrdat2_l_13(\CPU|DP|EXMEM|plif_exmem.rdat2_l [13]),
	.plif_exmemrdat2_l_14(\CPU|DP|EXMEM|plif_exmem.rdat2_l [14]),
	.plif_exmemrdat2_l_15(\CPU|DP|EXMEM|plif_exmem.rdat2_l [15]),
	.plif_exmemrdat2_l_16(\CPU|DP|EXMEM|plif_exmem.rdat2_l [16]),
	.plif_exmemrdat2_l_17(\CPU|DP|EXMEM|plif_exmem.rdat2_l [17]),
	.plif_exmemrdat2_l_18(\CPU|DP|EXMEM|plif_exmem.rdat2_l [18]),
	.plif_exmemrdat2_l_19(\CPU|DP|EXMEM|plif_exmem.rdat2_l [19]),
	.plif_exmemrdat2_l_20(\CPU|DP|EXMEM|plif_exmem.rdat2_l [20]),
	.plif_exmemrdat2_l_21(\CPU|DP|EXMEM|plif_exmem.rdat2_l [21]),
	.plif_exmemrdat2_l_22(\CPU|DP|EXMEM|plif_exmem.rdat2_l [22]),
	.plif_exmemrdat2_l_23(\CPU|DP|EXMEM|plif_exmem.rdat2_l [23]),
	.plif_exmemrdat2_l_24(\CPU|DP|EXMEM|plif_exmem.rdat2_l [24]),
	.plif_exmemrdat2_l_25(\CPU|DP|EXMEM|plif_exmem.rdat2_l [25]),
	.plif_exmemrdat2_l_26(\CPU|DP|EXMEM|plif_exmem.rdat2_l [26]),
	.plif_exmemrdat2_l_27(\CPU|DP|EXMEM|plif_exmem.rdat2_l [27]),
	.plif_exmemrdat2_l_28(\CPU|DP|EXMEM|plif_exmem.rdat2_l [28]),
	.plif_exmemrdat2_l_29(\CPU|DP|EXMEM|plif_exmem.rdat2_l [29]),
	.plif_exmemrdat2_l_30(\CPU|DP|EXMEM|plif_exmem.rdat2_l [30]),
	.plif_exmemrdat2_l_31(\CPU|DP|EXMEM|plif_exmem.rdat2_l [31]),
	.nRST(\nRST~input_o ),
	.CLK(\CPUCLK~clkctrl_outclk ),
	.nRST1(\nRST~inputclkctrl_outclk ),
	.devpor(devpor),
	.devclrn(devclrn),
	.devoe(devoe));

// Location: LCCOMB_X49_Y34_N20
cycloneive_lcell_comb \ramaddr~0 (
// Equation(s):
// \ramaddr~0_combout  = (plif_exmemdmemREN_l & (((plif_exmemporto_l_1)))) # (!plif_exmemdmemREN_l & ((plif_exmemdmemWEN_l & ((plif_exmemporto_l_1))) # (!plif_exmemdmemWEN_l & (PCreg_1))))

	.dataa(\CPU|DP|PC|PCreg [1]),
	.datab(\CPU|DP|EXMEM|plif_exmem.dmemREN_l~q ),
	.datac(\CPU|DP|EXMEM|plif_exmem.dmemWEN_l~q ),
	.datad(\CPU|DP|EXMEM|plif_exmem.porto_l [1]),
	.cin(gnd),
	.combout(\ramaddr~0_combout ),
	.cout());
// synopsys translate_off
defparam \ramaddr~0 .lut_mask = 16'hFE02;
defparam \ramaddr~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X49_Y34_N0
cycloneive_lcell_comb \ramaddr~1 (
// Equation(s):
// \ramaddr~1_combout  = (plif_exmemdmemWEN_l & (((plif_exmemporto_l_0)))) # (!plif_exmemdmemWEN_l & ((plif_exmemdmemREN_l & (plif_exmemporto_l_0)) # (!plif_exmemdmemREN_l & ((PCreg_0)))))

	.dataa(\CPU|DP|EXMEM|plif_exmem.dmemWEN_l~q ),
	.datab(\CPU|DP|EXMEM|plif_exmem.dmemREN_l~q ),
	.datac(\CPU|DP|EXMEM|plif_exmem.porto_l [0]),
	.datad(\CPU|DP|PC|PCreg [0]),
	.cin(gnd),
	.combout(\ramaddr~1_combout ),
	.cout());
// synopsys translate_off
defparam \ramaddr~1 .lut_mask = 16'hF1E0;
defparam \ramaddr~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y35_N6
cycloneive_lcell_comb \ramaddr~2 (
// Equation(s):
// \ramaddr~2_combout  = (plif_exmemdmemREN_l & (((plif_exmemporto_l_3)))) # (!plif_exmemdmemREN_l & ((plif_exmemdmemWEN_l & ((plif_exmemporto_l_3))) # (!plif_exmemdmemWEN_l & (PCreg_3))))

	.dataa(\CPU|DP|EXMEM|plif_exmem.dmemREN_l~q ),
	.datab(\CPU|DP|PC|PCreg [3]),
	.datac(\CPU|DP|EXMEM|plif_exmem.dmemWEN_l~q ),
	.datad(\CPU|DP|EXMEM|plif_exmem.porto_l [3]),
	.cin(gnd),
	.combout(\ramaddr~2_combout ),
	.cout());
// synopsys translate_off
defparam \ramaddr~2 .lut_mask = 16'hFE04;
defparam \ramaddr~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y35_N20
cycloneive_lcell_comb \ramaddr~3 (
// Equation(s):
// \ramaddr~3_combout  = (\syif.tbCTRL~input_o  & (\syif.addr[3]~input_o )) # (!\syif.tbCTRL~input_o  & ((\ramaddr~2_combout )))

	.dataa(\syif.tbCTRL~input_o ),
	.datab(gnd),
	.datac(\syif.addr[3]~input_o ),
	.datad(\ramaddr~2_combout ),
	.cin(gnd),
	.combout(\ramaddr~3_combout ),
	.cout());
// synopsys translate_off
defparam \ramaddr~3 .lut_mask = 16'hF5A0;
defparam \ramaddr~3 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y35_N28
cycloneive_lcell_comb \ramaddr~4 (
// Equation(s):
// \ramaddr~4_combout  = (plif_exmemdmemREN_l & (((plif_exmemporto_l_2)))) # (!plif_exmemdmemREN_l & ((plif_exmemdmemWEN_l & ((plif_exmemporto_l_2))) # (!plif_exmemdmemWEN_l & (PCreg_2))))

	.dataa(\CPU|DP|EXMEM|plif_exmem.dmemREN_l~q ),
	.datab(\CPU|DP|PC|PCreg [2]),
	.datac(\CPU|DP|EXMEM|plif_exmem.porto_l [2]),
	.datad(\CPU|DP|EXMEM|plif_exmem.dmemWEN_l~q ),
	.cin(gnd),
	.combout(\ramaddr~4_combout ),
	.cout());
// synopsys translate_off
defparam \ramaddr~4 .lut_mask = 16'hF0E4;
defparam \ramaddr~4 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y35_N14
cycloneive_lcell_comb \ramaddr~5 (
// Equation(s):
// \ramaddr~5_combout  = (\syif.tbCTRL~input_o  & (\syif.addr[2]~input_o )) # (!\syif.tbCTRL~input_o  & ((\ramaddr~4_combout )))

	.dataa(\syif.tbCTRL~input_o ),
	.datab(gnd),
	.datac(\syif.addr[2]~input_o ),
	.datad(\ramaddr~4_combout ),
	.cin(gnd),
	.combout(\ramaddr~5_combout ),
	.cout());
// synopsys translate_off
defparam \ramaddr~5 .lut_mask = 16'hF5A0;
defparam \ramaddr~5 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X49_Y34_N24
cycloneive_lcell_comb \ramaddr~6 (
// Equation(s):
// \ramaddr~6_combout  = (plif_exmemdmemWEN_l & (((plif_exmemporto_l_5)))) # (!plif_exmemdmemWEN_l & ((plif_exmemdmemREN_l & ((plif_exmemporto_l_5))) # (!plif_exmemdmemREN_l & (PCreg_5))))

	.dataa(\CPU|DP|PC|PCreg [5]),
	.datab(\CPU|DP|EXMEM|plif_exmem.dmemWEN_l~q ),
	.datac(\CPU|DP|EXMEM|plif_exmem.dmemREN_l~q ),
	.datad(\CPU|DP|EXMEM|plif_exmem.porto_l [5]),
	.cin(gnd),
	.combout(\ramaddr~6_combout ),
	.cout());
// synopsys translate_off
defparam \ramaddr~6 .lut_mask = 16'hFE02;
defparam \ramaddr~6 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X49_Y34_N6
cycloneive_lcell_comb \ramaddr~7 (
// Equation(s):
// \ramaddr~7_combout  = (\syif.tbCTRL~input_o  & (\syif.addr[5]~input_o )) # (!\syif.tbCTRL~input_o  & ((\ramaddr~6_combout )))

	.dataa(\syif.tbCTRL~input_o ),
	.datab(\syif.addr[5]~input_o ),
	.datac(gnd),
	.datad(\ramaddr~6_combout ),
	.cin(gnd),
	.combout(\ramaddr~7_combout ),
	.cout());
// synopsys translate_off
defparam \ramaddr~7 .lut_mask = 16'hDD88;
defparam \ramaddr~7 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X49_Y34_N18
cycloneive_lcell_comb \ramaddr~8 (
// Equation(s):
// \ramaddr~8_combout  = (plif_exmemdmemWEN_l & (((plif_exmemporto_l_4)))) # (!plif_exmemdmemWEN_l & ((plif_exmemdmemREN_l & ((plif_exmemporto_l_4))) # (!plif_exmemdmemREN_l & (PCreg_4))))

	.dataa(\CPU|DP|EXMEM|plif_exmem.dmemWEN_l~q ),
	.datab(\CPU|DP|PC|PCreg [4]),
	.datac(\CPU|DP|EXMEM|plif_exmem.dmemREN_l~q ),
	.datad(\CPU|DP|EXMEM|plif_exmem.porto_l [4]),
	.cin(gnd),
	.combout(\ramaddr~8_combout ),
	.cout());
// synopsys translate_off
defparam \ramaddr~8 .lut_mask = 16'hFE04;
defparam \ramaddr~8 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X49_Y34_N16
cycloneive_lcell_comb \ramaddr~9 (
// Equation(s):
// \ramaddr~9_combout  = (\syif.tbCTRL~input_o  & (\syif.addr[4]~input_o )) # (!\syif.tbCTRL~input_o  & ((\ramaddr~8_combout )))

	.dataa(\syif.tbCTRL~input_o ),
	.datab(\syif.addr[4]~input_o ),
	.datac(gnd),
	.datad(\ramaddr~8_combout ),
	.cin(gnd),
	.combout(\ramaddr~9_combout ),
	.cout());
// synopsys translate_off
defparam \ramaddr~9 .lut_mask = 16'hDD88;
defparam \ramaddr~9 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y34_N10
cycloneive_lcell_comb \ramaddr~10 (
// Equation(s):
// \ramaddr~10_combout  = (plif_exmemdmemREN_l & (((plif_exmemporto_l_7)))) # (!plif_exmemdmemREN_l & ((plif_exmemdmemWEN_l & ((plif_exmemporto_l_7))) # (!plif_exmemdmemWEN_l & (PCreg_7))))

	.dataa(\CPU|DP|EXMEM|plif_exmem.dmemREN_l~q ),
	.datab(\CPU|DP|PC|PCreg [7]),
	.datac(\CPU|DP|EXMEM|plif_exmem.dmemWEN_l~q ),
	.datad(\CPU|DP|EXMEM|plif_exmem.porto_l [7]),
	.cin(gnd),
	.combout(\ramaddr~10_combout ),
	.cout());
// synopsys translate_off
defparam \ramaddr~10 .lut_mask = 16'hFE04;
defparam \ramaddr~10 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y34_N16
cycloneive_lcell_comb \ramaddr~11 (
// Equation(s):
// \ramaddr~11_combout  = (\syif.tbCTRL~input_o  & (\syif.addr[7]~input_o )) # (!\syif.tbCTRL~input_o  & ((\ramaddr~10_combout )))

	.dataa(gnd),
	.datab(\syif.addr[7]~input_o ),
	.datac(\syif.tbCTRL~input_o ),
	.datad(\ramaddr~10_combout ),
	.cin(gnd),
	.combout(\ramaddr~11_combout ),
	.cout());
// synopsys translate_off
defparam \ramaddr~11 .lut_mask = 16'hCFC0;
defparam \ramaddr~11 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y34_N24
cycloneive_lcell_comb \ramaddr~12 (
// Equation(s):
// \ramaddr~12_combout  = (plif_exmemdmemREN_l & (((plif_exmemporto_l_6)))) # (!plif_exmemdmemREN_l & ((plif_exmemdmemWEN_l & ((plif_exmemporto_l_6))) # (!plif_exmemdmemWEN_l & (PCreg_6))))

	.dataa(\CPU|DP|PC|PCreg [6]),
	.datab(\CPU|DP|EXMEM|plif_exmem.dmemREN_l~q ),
	.datac(\CPU|DP|EXMEM|plif_exmem.dmemWEN_l~q ),
	.datad(\CPU|DP|EXMEM|plif_exmem.porto_l [6]),
	.cin(gnd),
	.combout(\ramaddr~12_combout ),
	.cout());
// synopsys translate_off
defparam \ramaddr~12 .lut_mask = 16'hFE02;
defparam \ramaddr~12 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y34_N6
cycloneive_lcell_comb \ramaddr~13 (
// Equation(s):
// \ramaddr~13_combout  = (\syif.tbCTRL~input_o  & (\syif.addr[6]~input_o )) # (!\syif.tbCTRL~input_o  & ((\ramaddr~12_combout )))

	.dataa(\syif.tbCTRL~input_o ),
	.datab(gnd),
	.datac(\syif.addr[6]~input_o ),
	.datad(\ramaddr~12_combout ),
	.cin(gnd),
	.combout(\ramaddr~13_combout ),
	.cout());
// synopsys translate_off
defparam \ramaddr~13 .lut_mask = 16'hF5A0;
defparam \ramaddr~13 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y33_N20
cycloneive_lcell_comb \ramaddr~14 (
// Equation(s):
// \ramaddr~14_combout  = (plif_exmemdmemWEN_l & (((plif_exmemporto_l_9)))) # (!plif_exmemdmemWEN_l & ((plif_exmemdmemREN_l & ((plif_exmemporto_l_9))) # (!plif_exmemdmemREN_l & (PCreg_9))))

	.dataa(\CPU|DP|PC|PCreg [9]),
	.datab(\CPU|DP|EXMEM|plif_exmem.dmemWEN_l~q ),
	.datac(\CPU|DP|EXMEM|plif_exmem.dmemREN_l~q ),
	.datad(\CPU|DP|EXMEM|plif_exmem.porto_l [9]),
	.cin(gnd),
	.combout(\ramaddr~14_combout ),
	.cout());
// synopsys translate_off
defparam \ramaddr~14 .lut_mask = 16'hFE02;
defparam \ramaddr~14 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y33_N10
cycloneive_lcell_comb \ramaddr~15 (
// Equation(s):
// \ramaddr~15_combout  = (\syif.tbCTRL~input_o  & (\syif.addr[9]~input_o )) # (!\syif.tbCTRL~input_o  & ((\ramaddr~14_combout )))

	.dataa(\syif.tbCTRL~input_o ),
	.datab(gnd),
	.datac(\syif.addr[9]~input_o ),
	.datad(\ramaddr~14_combout ),
	.cin(gnd),
	.combout(\ramaddr~15_combout ),
	.cout());
// synopsys translate_off
defparam \ramaddr~15 .lut_mask = 16'hF5A0;
defparam \ramaddr~15 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y33_N24
cycloneive_lcell_comb \ramaddr~16 (
// Equation(s):
// \ramaddr~16_combout  = (plif_exmemdmemWEN_l & (((plif_exmemporto_l_8)))) # (!plif_exmemdmemWEN_l & ((plif_exmemdmemREN_l & ((plif_exmemporto_l_8))) # (!plif_exmemdmemREN_l & (PCreg_8))))

	.dataa(\CPU|DP|PC|PCreg [8]),
	.datab(\CPU|DP|EXMEM|plif_exmem.dmemWEN_l~q ),
	.datac(\CPU|DP|EXMEM|plif_exmem.dmemREN_l~q ),
	.datad(\CPU|DP|EXMEM|plif_exmem.porto_l [8]),
	.cin(gnd),
	.combout(\ramaddr~16_combout ),
	.cout());
// synopsys translate_off
defparam \ramaddr~16 .lut_mask = 16'hFE02;
defparam \ramaddr~16 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y33_N8
cycloneive_lcell_comb \ramaddr~17 (
// Equation(s):
// \ramaddr~17_combout  = (\syif.tbCTRL~input_o  & (\syif.addr[8]~input_o )) # (!\syif.tbCTRL~input_o  & ((\ramaddr~16_combout )))

	.dataa(gnd),
	.datab(\syif.addr[8]~input_o ),
	.datac(\syif.tbCTRL~input_o ),
	.datad(\ramaddr~16_combout ),
	.cin(gnd),
	.combout(\ramaddr~17_combout ),
	.cout());
// synopsys translate_off
defparam \ramaddr~17 .lut_mask = 16'hCFC0;
defparam \ramaddr~17 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y37_N6
cycloneive_lcell_comb \ramaddr~18 (
// Equation(s):
// \ramaddr~18_combout  = (plif_exmemdmemREN_l & (plif_exmemporto_l_11)) # (!plif_exmemdmemREN_l & ((plif_exmemdmemWEN_l & (plif_exmemporto_l_11)) # (!plif_exmemdmemWEN_l & ((PCreg_11)))))

	.dataa(\CPU|DP|EXMEM|plif_exmem.porto_l [11]),
	.datab(\CPU|DP|EXMEM|plif_exmem.dmemREN_l~q ),
	.datac(\CPU|DP|PC|PCreg [11]),
	.datad(\CPU|DP|EXMEM|plif_exmem.dmemWEN_l~q ),
	.cin(gnd),
	.combout(\ramaddr~18_combout ),
	.cout());
// synopsys translate_off
defparam \ramaddr~18 .lut_mask = 16'hAAB8;
defparam \ramaddr~18 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y37_N22
cycloneive_lcell_comb \ramaddr~19 (
// Equation(s):
// \ramaddr~19_combout  = (\syif.tbCTRL~input_o  & (\syif.addr[11]~input_o )) # (!\syif.tbCTRL~input_o  & ((\ramaddr~18_combout )))

	.dataa(gnd),
	.datab(\syif.tbCTRL~input_o ),
	.datac(\syif.addr[11]~input_o ),
	.datad(\ramaddr~18_combout ),
	.cin(gnd),
	.combout(\ramaddr~19_combout ),
	.cout());
// synopsys translate_off
defparam \ramaddr~19 .lut_mask = 16'hF3C0;
defparam \ramaddr~19 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y37_N10
cycloneive_lcell_comb \ramaddr~20 (
// Equation(s):
// \ramaddr~20_combout  = (plif_exmemdmemREN_l & (((plif_exmemporto_l_10)))) # (!plif_exmemdmemREN_l & ((plif_exmemdmemWEN_l & ((plif_exmemporto_l_10))) # (!plif_exmemdmemWEN_l & (PCreg_10))))

	.dataa(\CPU|DP|PC|PCreg [10]),
	.datab(\CPU|DP|EXMEM|plif_exmem.porto_l [10]),
	.datac(\CPU|DP|EXMEM|plif_exmem.dmemREN_l~q ),
	.datad(\CPU|DP|EXMEM|plif_exmem.dmemWEN_l~q ),
	.cin(gnd),
	.combout(\ramaddr~20_combout ),
	.cout());
// synopsys translate_off
defparam \ramaddr~20 .lut_mask = 16'hCCCA;
defparam \ramaddr~20 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y37_N12
cycloneive_lcell_comb \ramaddr~21 (
// Equation(s):
// \ramaddr~21_combout  = (\syif.tbCTRL~input_o  & (\syif.addr[10]~input_o )) # (!\syif.tbCTRL~input_o  & ((\ramaddr~20_combout )))

	.dataa(\syif.tbCTRL~input_o ),
	.datab(\syif.addr[10]~input_o ),
	.datac(gnd),
	.datad(\ramaddr~20_combout ),
	.cin(gnd),
	.combout(\ramaddr~21_combout ),
	.cout());
// synopsys translate_off
defparam \ramaddr~21 .lut_mask = 16'hDD88;
defparam \ramaddr~21 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y32_N6
cycloneive_lcell_comb \ramaddr~22 (
// Equation(s):
// \ramaddr~22_combout  = (plif_exmemdmemREN_l & (((plif_exmemporto_l_13)))) # (!plif_exmemdmemREN_l & ((plif_exmemdmemWEN_l & ((plif_exmemporto_l_13))) # (!plif_exmemdmemWEN_l & (PCreg_13))))

	.dataa(\CPU|DP|EXMEM|plif_exmem.dmemREN_l~q ),
	.datab(\CPU|DP|EXMEM|plif_exmem.dmemWEN_l~q ),
	.datac(\CPU|DP|PC|PCreg [13]),
	.datad(\CPU|DP|EXMEM|plif_exmem.porto_l [13]),
	.cin(gnd),
	.combout(\ramaddr~22_combout ),
	.cout());
// synopsys translate_off
defparam \ramaddr~22 .lut_mask = 16'hFE10;
defparam \ramaddr~22 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y32_N24
cycloneive_lcell_comb \ramaddr~23 (
// Equation(s):
// \ramaddr~23_combout  = (\syif.tbCTRL~input_o  & (\syif.addr[13]~input_o )) # (!\syif.tbCTRL~input_o  & ((\ramaddr~22_combout )))

	.dataa(\syif.tbCTRL~input_o ),
	.datab(gnd),
	.datac(\syif.addr[13]~input_o ),
	.datad(\ramaddr~22_combout ),
	.cin(gnd),
	.combout(\ramaddr~23_combout ),
	.cout());
// synopsys translate_off
defparam \ramaddr~23 .lut_mask = 16'hF5A0;
defparam \ramaddr~23 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y32_N28
cycloneive_lcell_comb \ramaddr~24 (
// Equation(s):
// \ramaddr~24_combout  = (plif_exmemdmemREN_l & (((plif_exmemporto_l_12)))) # (!plif_exmemdmemREN_l & ((plif_exmemdmemWEN_l & ((plif_exmemporto_l_12))) # (!plif_exmemdmemWEN_l & (PCreg_12))))

	.dataa(\CPU|DP|EXMEM|plif_exmem.dmemREN_l~q ),
	.datab(\CPU|DP|PC|PCreg [12]),
	.datac(\CPU|DP|EXMEM|plif_exmem.porto_l [12]),
	.datad(\CPU|DP|EXMEM|plif_exmem.dmemWEN_l~q ),
	.cin(gnd),
	.combout(\ramaddr~24_combout ),
	.cout());
// synopsys translate_off
defparam \ramaddr~24 .lut_mask = 16'hF0E4;
defparam \ramaddr~24 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y32_N2
cycloneive_lcell_comb \ramaddr~25 (
// Equation(s):
// \ramaddr~25_combout  = (\syif.tbCTRL~input_o  & (\syif.addr[12]~input_o )) # (!\syif.tbCTRL~input_o  & ((\ramaddr~24_combout )))

	.dataa(\syif.tbCTRL~input_o ),
	.datab(gnd),
	.datac(\syif.addr[12]~input_o ),
	.datad(\ramaddr~24_combout ),
	.cin(gnd),
	.combout(\ramaddr~25_combout ),
	.cout());
// synopsys translate_off
defparam \ramaddr~25 .lut_mask = 16'hF5A0;
defparam \ramaddr~25 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X52_Y34_N2
cycloneive_lcell_comb \ramaddr~26 (
// Equation(s):
// \ramaddr~26_combout  = (plif_exmemdmemWEN_l & (((plif_exmemporto_l_15)))) # (!plif_exmemdmemWEN_l & ((plif_exmemdmemREN_l & ((plif_exmemporto_l_15))) # (!plif_exmemdmemREN_l & (PCreg_15))))

	.dataa(\CPU|DP|EXMEM|plif_exmem.dmemWEN_l~q ),
	.datab(\CPU|DP|PC|PCreg [15]),
	.datac(\CPU|DP|EXMEM|plif_exmem.porto_l [15]),
	.datad(\CPU|DP|EXMEM|plif_exmem.dmemREN_l~q ),
	.cin(gnd),
	.combout(\ramaddr~26_combout ),
	.cout());
// synopsys translate_off
defparam \ramaddr~26 .lut_mask = 16'hF0E4;
defparam \ramaddr~26 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X52_Y34_N12
cycloneive_lcell_comb \ramaddr~27 (
// Equation(s):
// \ramaddr~27_combout  = (\syif.tbCTRL~input_o  & (!\syif.addr[15]~input_o )) # (!\syif.tbCTRL~input_o  & ((!\ramaddr~26_combout )))

	.dataa(gnd),
	.datab(\syif.addr[15]~input_o ),
	.datac(\syif.tbCTRL~input_o ),
	.datad(\ramaddr~26_combout ),
	.cin(gnd),
	.combout(\ramaddr~27_combout ),
	.cout());
// synopsys translate_off
defparam \ramaddr~27 .lut_mask = 16'h303F;
defparam \ramaddr~27 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X52_Y34_N24
cycloneive_lcell_comb \ramaddr~28 (
// Equation(s):
// \ramaddr~28_combout  = (plif_exmemdmemREN_l & (((plif_exmemporto_l_14)))) # (!plif_exmemdmemREN_l & ((plif_exmemdmemWEN_l & ((plif_exmemporto_l_14))) # (!plif_exmemdmemWEN_l & (PCreg_14))))

	.dataa(\CPU|DP|EXMEM|plif_exmem.dmemREN_l~q ),
	.datab(\CPU|DP|PC|PCreg [14]),
	.datac(\CPU|DP|EXMEM|plif_exmem.dmemWEN_l~q ),
	.datad(\CPU|DP|EXMEM|plif_exmem.porto_l [14]),
	.cin(gnd),
	.combout(\ramaddr~28_combout ),
	.cout());
// synopsys translate_off
defparam \ramaddr~28 .lut_mask = 16'hFE04;
defparam \ramaddr~28 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X52_Y34_N6
cycloneive_lcell_comb \ramaddr~29 (
// Equation(s):
// \ramaddr~29_combout  = (\syif.tbCTRL~input_o  & (\syif.addr[14]~input_o )) # (!\syif.tbCTRL~input_o  & ((\ramaddr~28_combout )))

	.dataa(\syif.addr[14]~input_o ),
	.datab(gnd),
	.datac(\syif.tbCTRL~input_o ),
	.datad(\ramaddr~28_combout ),
	.cin(gnd),
	.combout(\ramaddr~29_combout ),
	.cout());
// synopsys translate_off
defparam \ramaddr~29 .lut_mask = 16'hAFA0;
defparam \ramaddr~29 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X50_Y34_N2
cycloneive_lcell_comb \ramaddr~30 (
// Equation(s):
// \ramaddr~30_combout  = (plif_exmemdmemWEN_l & (((plif_exmemporto_l_17)))) # (!plif_exmemdmemWEN_l & ((plif_exmemdmemREN_l & ((plif_exmemporto_l_17))) # (!plif_exmemdmemREN_l & (PCreg_17))))

	.dataa(\CPU|DP|EXMEM|plif_exmem.dmemWEN_l~q ),
	.datab(\CPU|DP|EXMEM|plif_exmem.dmemREN_l~q ),
	.datac(\CPU|DP|PC|PCreg [17]),
	.datad(\CPU|DP|EXMEM|plif_exmem.porto_l [17]),
	.cin(gnd),
	.combout(\ramaddr~30_combout ),
	.cout());
// synopsys translate_off
defparam \ramaddr~30 .lut_mask = 16'hFE10;
defparam \ramaddr~30 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X50_Y34_N10
cycloneive_lcell_comb \ramaddr~31 (
// Equation(s):
// \ramaddr~31_combout  = (\syif.tbCTRL~input_o  & (\syif.addr[17]~input_o )) # (!\syif.tbCTRL~input_o  & ((\ramaddr~30_combout )))

	.dataa(\syif.tbCTRL~input_o ),
	.datab(gnd),
	.datac(\syif.addr[17]~input_o ),
	.datad(\ramaddr~30_combout ),
	.cin(gnd),
	.combout(\ramaddr~31_combout ),
	.cout());
// synopsys translate_off
defparam \ramaddr~31 .lut_mask = 16'hF5A0;
defparam \ramaddr~31 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X50_Y34_N18
cycloneive_lcell_comb \ramaddr~32 (
// Equation(s):
// \ramaddr~32_combout  = (plif_exmemdmemWEN_l & (((plif_exmemporto_l_16)))) # (!plif_exmemdmemWEN_l & ((plif_exmemdmemREN_l & ((plif_exmemporto_l_16))) # (!plif_exmemdmemREN_l & (PCreg_16))))

	.dataa(\CPU|DP|EXMEM|plif_exmem.dmemWEN_l~q ),
	.datab(\CPU|DP|PC|PCreg [16]),
	.datac(\CPU|DP|EXMEM|plif_exmem.porto_l [16]),
	.datad(\CPU|DP|EXMEM|plif_exmem.dmemREN_l~q ),
	.cin(gnd),
	.combout(\ramaddr~32_combout ),
	.cout());
// synopsys translate_off
defparam \ramaddr~32 .lut_mask = 16'hF0E4;
defparam \ramaddr~32 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X50_Y34_N8
cycloneive_lcell_comb \ramaddr~33 (
// Equation(s):
// \ramaddr~33_combout  = (\syif.tbCTRL~input_o  & (\syif.addr[16]~input_o )) # (!\syif.tbCTRL~input_o  & ((\ramaddr~32_combout )))

	.dataa(gnd),
	.datab(\syif.addr[16]~input_o ),
	.datac(\syif.tbCTRL~input_o ),
	.datad(\ramaddr~32_combout ),
	.cin(gnd),
	.combout(\ramaddr~33_combout ),
	.cout());
// synopsys translate_off
defparam \ramaddr~33 .lut_mask = 16'hCFC0;
defparam \ramaddr~33 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y33_N18
cycloneive_lcell_comb \ramaddr~34 (
// Equation(s):
// \ramaddr~34_combout  = (plif_exmemdmemREN_l & (((plif_exmemporto_l_19)))) # (!plif_exmemdmemREN_l & ((plif_exmemdmemWEN_l & ((plif_exmemporto_l_19))) # (!plif_exmemdmemWEN_l & (PCreg_19))))

	.dataa(\CPU|DP|EXMEM|plif_exmem.dmemREN_l~q ),
	.datab(\CPU|DP|PC|PCreg [19]),
	.datac(\CPU|DP|EXMEM|plif_exmem.dmemWEN_l~q ),
	.datad(\CPU|DP|EXMEM|plif_exmem.porto_l [19]),
	.cin(gnd),
	.combout(\ramaddr~34_combout ),
	.cout());
// synopsys translate_off
defparam \ramaddr~34 .lut_mask = 16'hFE04;
defparam \ramaddr~34 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y33_N2
cycloneive_lcell_comb \ramaddr~35 (
// Equation(s):
// \ramaddr~35_combout  = (\syif.tbCTRL~input_o  & (\syif.addr[19]~input_o )) # (!\syif.tbCTRL~input_o  & ((\ramaddr~34_combout )))

	.dataa(\syif.tbCTRL~input_o ),
	.datab(gnd),
	.datac(\syif.addr[19]~input_o ),
	.datad(\ramaddr~34_combout ),
	.cin(gnd),
	.combout(\ramaddr~35_combout ),
	.cout());
// synopsys translate_off
defparam \ramaddr~35 .lut_mask = 16'hF5A0;
defparam \ramaddr~35 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y33_N6
cycloneive_lcell_comb \ramaddr~36 (
// Equation(s):
// \ramaddr~36_combout  = (plif_exmemdmemREN_l & (((plif_exmemporto_l_18)))) # (!plif_exmemdmemREN_l & ((plif_exmemdmemWEN_l & ((plif_exmemporto_l_18))) # (!plif_exmemdmemWEN_l & (PCreg_18))))

	.dataa(\CPU|DP|EXMEM|plif_exmem.dmemREN_l~q ),
	.datab(\CPU|DP|PC|PCreg [18]),
	.datac(\CPU|DP|EXMEM|plif_exmem.dmemWEN_l~q ),
	.datad(\CPU|DP|EXMEM|plif_exmem.porto_l [18]),
	.cin(gnd),
	.combout(\ramaddr~36_combout ),
	.cout());
// synopsys translate_off
defparam \ramaddr~36 .lut_mask = 16'hFE04;
defparam \ramaddr~36 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y33_N16
cycloneive_lcell_comb \ramaddr~37 (
// Equation(s):
// \ramaddr~37_combout  = (\syif.tbCTRL~input_o  & (\syif.addr[18]~input_o )) # (!\syif.tbCTRL~input_o  & ((\ramaddr~36_combout )))

	.dataa(\syif.tbCTRL~input_o ),
	.datab(gnd),
	.datac(\syif.addr[18]~input_o ),
	.datad(\ramaddr~36_combout ),
	.cin(gnd),
	.combout(\ramaddr~37_combout ),
	.cout());
// synopsys translate_off
defparam \ramaddr~37 .lut_mask = 16'hF5A0;
defparam \ramaddr~37 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y34_N20
cycloneive_lcell_comb \ramaddr~38 (
// Equation(s):
// \ramaddr~38_combout  = (\syif.tbCTRL~input_o  & (\syif.addr[21]~input_o )) # (!\syif.tbCTRL~input_o  & (((plif_exmemdmemREN_l) # (plif_exmemdmemWEN_l))))

	.dataa(\syif.addr[21]~input_o ),
	.datab(\CPU|DP|EXMEM|plif_exmem.dmemREN_l~q ),
	.datac(\CPU|DP|EXMEM|plif_exmem.dmemWEN_l~q ),
	.datad(\syif.tbCTRL~input_o ),
	.cin(gnd),
	.combout(\ramaddr~38_combout ),
	.cout());
// synopsys translate_off
defparam \ramaddr~38 .lut_mask = 16'hAAFC;
defparam \ramaddr~38 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y34_N10
cycloneive_lcell_comb \ramaddr~39 (
// Equation(s):
// \ramaddr~39_combout  = (\syif.tbCTRL~input_o  & (((\ramaddr~38_combout )))) # (!\syif.tbCTRL~input_o  & ((\ramaddr~38_combout  & (plif_exmemporto_l_21)) # (!\ramaddr~38_combout  & ((PCreg_21)))))

	.dataa(\syif.tbCTRL~input_o ),
	.datab(\CPU|DP|EXMEM|plif_exmem.porto_l [21]),
	.datac(\CPU|DP|PC|PCreg [21]),
	.datad(\ramaddr~38_combout ),
	.cin(gnd),
	.combout(\ramaddr~39_combout ),
	.cout());
// synopsys translate_off
defparam \ramaddr~39 .lut_mask = 16'hEE50;
defparam \ramaddr~39 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y34_N28
cycloneive_lcell_comb \ramaddr~40 (
// Equation(s):
// \ramaddr~40_combout  = (plif_exmemdmemWEN_l & (((plif_exmemporto_l_20)))) # (!plif_exmemdmemWEN_l & ((plif_exmemdmemREN_l & ((plif_exmemporto_l_20))) # (!plif_exmemdmemREN_l & (PCreg_20))))

	.dataa(\CPU|DP|PC|PCreg [20]),
	.datab(\CPU|DP|EXMEM|plif_exmem.dmemWEN_l~q ),
	.datac(\CPU|DP|EXMEM|plif_exmem.dmemREN_l~q ),
	.datad(\CPU|DP|EXMEM|plif_exmem.porto_l [20]),
	.cin(gnd),
	.combout(\ramaddr~40_combout ),
	.cout());
// synopsys translate_off
defparam \ramaddr~40 .lut_mask = 16'hFE02;
defparam \ramaddr~40 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y34_N0
cycloneive_lcell_comb \ramaddr~41 (
// Equation(s):
// \ramaddr~41_combout  = (\syif.tbCTRL~input_o  & (\syif.addr[20]~input_o )) # (!\syif.tbCTRL~input_o  & ((\ramaddr~40_combout )))

	.dataa(gnd),
	.datab(\syif.tbCTRL~input_o ),
	.datac(\syif.addr[20]~input_o ),
	.datad(\ramaddr~40_combout ),
	.cin(gnd),
	.combout(\ramaddr~41_combout ),
	.cout());
// synopsys translate_off
defparam \ramaddr~41 .lut_mask = 16'hF3C0;
defparam \ramaddr~41 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y34_N16
cycloneive_lcell_comb \ramaddr~42 (
// Equation(s):
// \ramaddr~42_combout  = (plif_exmemdmemWEN_l & (((plif_exmemporto_l_23)))) # (!plif_exmemdmemWEN_l & ((plif_exmemdmemREN_l & ((plif_exmemporto_l_23))) # (!plif_exmemdmemREN_l & (PCreg_23))))

	.dataa(\CPU|DP|PC|PCreg [23]),
	.datab(\CPU|DP|EXMEM|plif_exmem.dmemWEN_l~q ),
	.datac(\CPU|DP|EXMEM|plif_exmem.dmemREN_l~q ),
	.datad(\CPU|DP|EXMEM|plif_exmem.porto_l [23]),
	.cin(gnd),
	.combout(\ramaddr~42_combout ),
	.cout());
// synopsys translate_off
defparam \ramaddr~42 .lut_mask = 16'hFE02;
defparam \ramaddr~42 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y34_N18
cycloneive_lcell_comb \ramaddr~43 (
// Equation(s):
// \ramaddr~43_combout  = (\syif.tbCTRL~input_o  & (\syif.addr[23]~input_o )) # (!\syif.tbCTRL~input_o  & ((\ramaddr~42_combout )))

	.dataa(\syif.addr[23]~input_o ),
	.datab(gnd),
	.datac(\syif.tbCTRL~input_o ),
	.datad(\ramaddr~42_combout ),
	.cin(gnd),
	.combout(\ramaddr~43_combout ),
	.cout());
// synopsys translate_off
defparam \ramaddr~43 .lut_mask = 16'hAFA0;
defparam \ramaddr~43 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y34_N22
cycloneive_lcell_comb \ramaddr~44 (
// Equation(s):
// \ramaddr~44_combout  = (plif_exmemdmemWEN_l & (((plif_exmemporto_l_22)))) # (!plif_exmemdmemWEN_l & ((plif_exmemdmemREN_l & ((plif_exmemporto_l_22))) # (!plif_exmemdmemREN_l & (PCreg_22))))

	.dataa(\CPU|DP|PC|PCreg [22]),
	.datab(\CPU|DP|EXMEM|plif_exmem.dmemWEN_l~q ),
	.datac(\CPU|DP|EXMEM|plif_exmem.porto_l [22]),
	.datad(\CPU|DP|EXMEM|plif_exmem.dmemREN_l~q ),
	.cin(gnd),
	.combout(\ramaddr~44_combout ),
	.cout());
// synopsys translate_off
defparam \ramaddr~44 .lut_mask = 16'hF0E2;
defparam \ramaddr~44 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y34_N8
cycloneive_lcell_comb \ramaddr~45 (
// Equation(s):
// \ramaddr~45_combout  = (\syif.tbCTRL~input_o  & (\syif.addr[22]~input_o )) # (!\syif.tbCTRL~input_o  & ((\ramaddr~44_combout )))

	.dataa(\syif.tbCTRL~input_o ),
	.datab(\syif.addr[22]~input_o ),
	.datac(\ramaddr~44_combout ),
	.datad(gnd),
	.cin(gnd),
	.combout(\ramaddr~45_combout ),
	.cout());
// synopsys translate_off
defparam \ramaddr~45 .lut_mask = 16'hD8D8;
defparam \ramaddr~45 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y34_N14
cycloneive_lcell_comb \ramaddr~46 (
// Equation(s):
// \ramaddr~46_combout  = (\syif.tbCTRL~input_o  & (\syif.addr[25]~input_o )) # (!\syif.tbCTRL~input_o  & (((plif_exmemdmemREN_l) # (plif_exmemdmemWEN_l))))

	.dataa(\syif.tbCTRL~input_o ),
	.datab(\syif.addr[25]~input_o ),
	.datac(\CPU|DP|EXMEM|plif_exmem.dmemREN_l~q ),
	.datad(\CPU|DP|EXMEM|plif_exmem.dmemWEN_l~q ),
	.cin(gnd),
	.combout(\ramaddr~46_combout ),
	.cout());
// synopsys translate_off
defparam \ramaddr~46 .lut_mask = 16'hDDD8;
defparam \ramaddr~46 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y35_N4
cycloneive_lcell_comb \ramaddr~47 (
// Equation(s):
// \ramaddr~47_combout  = (\syif.tbCTRL~input_o  & (((\ramaddr~46_combout )))) # (!\syif.tbCTRL~input_o  & ((\ramaddr~46_combout  & ((plif_exmemporto_l_25))) # (!\ramaddr~46_combout  & (PCreg_25))))

	.dataa(\syif.tbCTRL~input_o ),
	.datab(\CPU|DP|PC|PCreg [25]),
	.datac(\ramaddr~46_combout ),
	.datad(\CPU|DP|EXMEM|plif_exmem.porto_l [25]),
	.cin(gnd),
	.combout(\ramaddr~47_combout ),
	.cout());
// synopsys translate_off
defparam \ramaddr~47 .lut_mask = 16'hF4A4;
defparam \ramaddr~47 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y35_N10
cycloneive_lcell_comb \ramaddr~48 (
// Equation(s):
// \ramaddr~48_combout  = (plif_exmemdmemWEN_l & (plif_exmemporto_l_24)) # (!plif_exmemdmemWEN_l & ((plif_exmemdmemREN_l & (plif_exmemporto_l_24)) # (!plif_exmemdmemREN_l & ((PCreg_24)))))

	.dataa(\CPU|DP|EXMEM|plif_exmem.porto_l [24]),
	.datab(\CPU|DP|PC|PCreg [24]),
	.datac(\CPU|DP|EXMEM|plif_exmem.dmemWEN_l~q ),
	.datad(\CPU|DP|EXMEM|plif_exmem.dmemREN_l~q ),
	.cin(gnd),
	.combout(\ramaddr~48_combout ),
	.cout());
// synopsys translate_off
defparam \ramaddr~48 .lut_mask = 16'hAAAC;
defparam \ramaddr~48 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y35_N8
cycloneive_lcell_comb \ramaddr~49 (
// Equation(s):
// \ramaddr~49_combout  = (\syif.tbCTRL~input_o  & (\syif.addr[24]~input_o )) # (!\syif.tbCTRL~input_o  & ((\ramaddr~48_combout )))

	.dataa(\syif.tbCTRL~input_o ),
	.datab(gnd),
	.datac(\syif.addr[24]~input_o ),
	.datad(\ramaddr~48_combout ),
	.cin(gnd),
	.combout(\ramaddr~49_combout ),
	.cout());
// synopsys translate_off
defparam \ramaddr~49 .lut_mask = 16'hF5A0;
defparam \ramaddr~49 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y33_N22
cycloneive_lcell_comb \ramaddr~50 (
// Equation(s):
// \ramaddr~50_combout  = (plif_exmemdmemREN_l & (plif_exmemporto_l_27)) # (!plif_exmemdmemREN_l & ((plif_exmemdmemWEN_l & (plif_exmemporto_l_27)) # (!plif_exmemdmemWEN_l & ((PCreg_27)))))

	.dataa(\CPU|DP|EXMEM|plif_exmem.porto_l [27]),
	.datab(\CPU|DP|PC|PCreg [27]),
	.datac(\CPU|DP|EXMEM|plif_exmem.dmemREN_l~q ),
	.datad(\CPU|DP|EXMEM|plif_exmem.dmemWEN_l~q ),
	.cin(gnd),
	.combout(\ramaddr~50_combout ),
	.cout());
// synopsys translate_off
defparam \ramaddr~50 .lut_mask = 16'hAAAC;
defparam \ramaddr~50 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y34_N6
cycloneive_lcell_comb \ramaddr~51 (
// Equation(s):
// \ramaddr~51_combout  = (\syif.tbCTRL~input_o  & (\syif.addr[27]~input_o )) # (!\syif.tbCTRL~input_o  & ((\ramaddr~50_combout )))

	.dataa(gnd),
	.datab(\syif.addr[27]~input_o ),
	.datac(\syif.tbCTRL~input_o ),
	.datad(\ramaddr~50_combout ),
	.cin(gnd),
	.combout(\ramaddr~51_combout ),
	.cout());
// synopsys translate_off
defparam \ramaddr~51 .lut_mask = 16'hCFC0;
defparam \ramaddr~51 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y36_N18
cycloneive_lcell_comb \ramaddr~52 (
// Equation(s):
// \ramaddr~52_combout  = (plif_exmemdmemWEN_l & (plif_exmemporto_l_26)) # (!plif_exmemdmemWEN_l & ((plif_exmemdmemREN_l & (plif_exmemporto_l_26)) # (!plif_exmemdmemREN_l & ((PCreg_26)))))

	.dataa(\CPU|DP|EXMEM|plif_exmem.dmemWEN_l~q ),
	.datab(\CPU|DP|EXMEM|plif_exmem.porto_l [26]),
	.datac(\CPU|DP|PC|PCreg [26]),
	.datad(\CPU|DP|EXMEM|plif_exmem.dmemREN_l~q ),
	.cin(gnd),
	.combout(\ramaddr~52_combout ),
	.cout());
// synopsys translate_off
defparam \ramaddr~52 .lut_mask = 16'hCCD8;
defparam \ramaddr~52 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y34_N16
cycloneive_lcell_comb \ramaddr~53 (
// Equation(s):
// \ramaddr~53_combout  = (\syif.tbCTRL~input_o  & (\syif.addr[26]~input_o )) # (!\syif.tbCTRL~input_o  & ((\ramaddr~52_combout )))

	.dataa(gnd),
	.datab(\syif.addr[26]~input_o ),
	.datac(\syif.tbCTRL~input_o ),
	.datad(\ramaddr~52_combout ),
	.cin(gnd),
	.combout(\ramaddr~53_combout ),
	.cout());
// synopsys translate_off
defparam \ramaddr~53 .lut_mask = 16'hCFC0;
defparam \ramaddr~53 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X50_Y34_N16
cycloneive_lcell_comb \ramaddr~54 (
// Equation(s):
// \ramaddr~54_combout  = (plif_exmemdmemREN_l & (((plif_exmemporto_l_29)))) # (!plif_exmemdmemREN_l & ((plif_exmemdmemWEN_l & ((plif_exmemporto_l_29))) # (!plif_exmemdmemWEN_l & (PCreg_29))))

	.dataa(\CPU|DP|PC|PCreg [29]),
	.datab(\CPU|DP|EXMEM|plif_exmem.dmemREN_l~q ),
	.datac(\CPU|DP|EXMEM|plif_exmem.dmemWEN_l~q ),
	.datad(\CPU|DP|EXMEM|plif_exmem.porto_l [29]),
	.cin(gnd),
	.combout(\ramaddr~54_combout ),
	.cout());
// synopsys translate_off
defparam \ramaddr~54 .lut_mask = 16'hFE02;
defparam \ramaddr~54 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X50_Y34_N12
cycloneive_lcell_comb \ramaddr~55 (
// Equation(s):
// \ramaddr~55_combout  = (\syif.tbCTRL~input_o  & (\syif.addr[29]~input_o )) # (!\syif.tbCTRL~input_o  & ((\ramaddr~54_combout )))

	.dataa(\syif.tbCTRL~input_o ),
	.datab(gnd),
	.datac(\syif.addr[29]~input_o ),
	.datad(\ramaddr~54_combout ),
	.cin(gnd),
	.combout(\ramaddr~55_combout ),
	.cout());
// synopsys translate_off
defparam \ramaddr~55 .lut_mask = 16'hF5A0;
defparam \ramaddr~55 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X50_Y34_N20
cycloneive_lcell_comb \ramaddr~56 (
// Equation(s):
// \ramaddr~56_combout  = (plif_exmemdmemREN_l & (((plif_exmemporto_l_28)))) # (!plif_exmemdmemREN_l & ((plif_exmemdmemWEN_l & ((plif_exmemporto_l_28))) # (!plif_exmemdmemWEN_l & (PCreg_28))))

	.dataa(\CPU|DP|EXMEM|plif_exmem.dmemREN_l~q ),
	.datab(\CPU|DP|PC|PCreg [28]),
	.datac(\CPU|DP|EXMEM|plif_exmem.dmemWEN_l~q ),
	.datad(\CPU|DP|EXMEM|plif_exmem.porto_l [28]),
	.cin(gnd),
	.combout(\ramaddr~56_combout ),
	.cout());
// synopsys translate_off
defparam \ramaddr~56 .lut_mask = 16'hFE04;
defparam \ramaddr~56 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X50_Y34_N26
cycloneive_lcell_comb \ramaddr~57 (
// Equation(s):
// \ramaddr~57_combout  = (\syif.tbCTRL~input_o  & (\syif.addr[28]~input_o )) # (!\syif.tbCTRL~input_o  & ((\ramaddr~56_combout )))

	.dataa(\syif.tbCTRL~input_o ),
	.datab(gnd),
	.datac(\syif.addr[28]~input_o ),
	.datad(\ramaddr~56_combout ),
	.cin(gnd),
	.combout(\ramaddr~57_combout ),
	.cout());
// synopsys translate_off
defparam \ramaddr~57 .lut_mask = 16'hF5A0;
defparam \ramaddr~57 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y34_N12
cycloneive_lcell_comb \ramaddr~58 (
// Equation(s):
// \ramaddr~58_combout  = (plif_exmemdmemREN_l & (((plif_exmemporto_l_31)))) # (!plif_exmemdmemREN_l & ((plif_exmemdmemWEN_l & (plif_exmemporto_l_31)) # (!plif_exmemdmemWEN_l & ((PCreg_31)))))

	.dataa(\CPU|DP|EXMEM|plif_exmem.dmemREN_l~q ),
	.datab(\CPU|DP|EXMEM|plif_exmem.dmemWEN_l~q ),
	.datac(\CPU|DP|EXMEM|plif_exmem.porto_l [31]),
	.datad(\CPU|DP|PC|PCreg [31]),
	.cin(gnd),
	.combout(\ramaddr~58_combout ),
	.cout());
// synopsys translate_off
defparam \ramaddr~58 .lut_mask = 16'hF1E0;
defparam \ramaddr~58 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y34_N2
cycloneive_lcell_comb \ramaddr~59 (
// Equation(s):
// \ramaddr~59_combout  = (\syif.tbCTRL~input_o  & (\syif.addr[31]~input_o )) # (!\syif.tbCTRL~input_o  & ((\ramaddr~58_combout )))

	.dataa(gnd),
	.datab(\syif.addr[31]~input_o ),
	.datac(\syif.tbCTRL~input_o ),
	.datad(\ramaddr~58_combout ),
	.cin(gnd),
	.combout(\ramaddr~59_combout ),
	.cout());
// synopsys translate_off
defparam \ramaddr~59 .lut_mask = 16'hCFC0;
defparam \ramaddr~59 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y34_N6
cycloneive_lcell_comb \ramaddr~60 (
// Equation(s):
// \ramaddr~60_combout  = (plif_exmemdmemWEN_l & (((plif_exmemporto_l_30)))) # (!plif_exmemdmemWEN_l & ((plif_exmemdmemREN_l & ((plif_exmemporto_l_30))) # (!plif_exmemdmemREN_l & (PCreg_30))))

	.dataa(\CPU|DP|PC|PCreg [30]),
	.datab(\CPU|DP|EXMEM|plif_exmem.dmemWEN_l~q ),
	.datac(\CPU|DP|EXMEM|plif_exmem.dmemREN_l~q ),
	.datad(\CPU|DP|EXMEM|plif_exmem.porto_l [30]),
	.cin(gnd),
	.combout(\ramaddr~60_combout ),
	.cout());
// synopsys translate_off
defparam \ramaddr~60 .lut_mask = 16'hFE02;
defparam \ramaddr~60 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y34_N24
cycloneive_lcell_comb \ramaddr~61 (
// Equation(s):
// \ramaddr~61_combout  = (\syif.tbCTRL~input_o  & (\syif.addr[30]~input_o )) # (!\syif.tbCTRL~input_o  & ((\ramaddr~60_combout )))

	.dataa(gnd),
	.datab(\syif.addr[30]~input_o ),
	.datac(\syif.tbCTRL~input_o ),
	.datad(\ramaddr~60_combout ),
	.cin(gnd),
	.combout(\ramaddr~61_combout ),
	.cout());
// synopsys translate_off
defparam \ramaddr~61 .lut_mask = 16'hCFC0;
defparam \ramaddr~61 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y34_N10
cycloneive_lcell_comb \ramWEN~0 (
// Equation(s):
// \ramWEN~0_combout  = (\syif.tbCTRL~input_o  & (!\syif.WEN~input_o )) # (!\syif.tbCTRL~input_o  & ((!plif_exmemdmemWEN_l)))

	.dataa(gnd),
	.datab(\syif.tbCTRL~input_o ),
	.datac(\syif.WEN~input_o ),
	.datad(\CPU|DP|EXMEM|plif_exmem.dmemWEN_l~q ),
	.cin(gnd),
	.combout(\ramWEN~0_combout ),
	.cout());
// synopsys translate_off
defparam \ramWEN~0 .lut_mask = 16'h0C3F;
defparam \ramWEN~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y33_N10
cycloneive_lcell_comb \ramREN~0 (
// Equation(s):
// \ramREN~0_combout  = (!\syif.tbCTRL~input_o  & ((plif_exmemdmemREN_l) # ((!dpifimemREN & !plif_exmemdmemWEN_l))))

	.dataa(\CPU|DP|EXMEM|plif_exmem.dmemREN_l~q ),
	.datab(\CPU|DP|dpif.imemREN~q ),
	.datac(\syif.tbCTRL~input_o ),
	.datad(\CPU|DP|EXMEM|plif_exmem.dmemWEN_l~q ),
	.cin(gnd),
	.combout(\ramREN~0_combout ),
	.cout());
// synopsys translate_off
defparam \ramREN~0 .lut_mask = 16'h0A0B;
defparam \ramREN~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y34_N28
cycloneive_lcell_comb \ramREN~1 (
// Equation(s):
// \ramREN~1_combout  = (!\ramREN~0_combout  & ((!\syif.tbCTRL~input_o ) # (!\syif.REN~input_o )))

	.dataa(\syif.REN~input_o ),
	.datab(gnd),
	.datac(\syif.tbCTRL~input_o ),
	.datad(\ramREN~0_combout ),
	.cin(gnd),
	.combout(\ramREN~1_combout ),
	.cout());
// synopsys translate_off
defparam \ramREN~1 .lut_mask = 16'h005F;
defparam \ramREN~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X59_Y1_N25
dffeas CPUCLK(
	.clk(\CLK~inputclkctrl_outclk ),
	.d(\CPUCLK~0_combout ),
	.asdata(vcc),
	.clrn(\nRST~inputclkctrl_outclk ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\CPUCLK~q ),
	.prn(vcc));
// synopsys translate_off
defparam CPUCLK.is_wysiwyg = "true";
defparam CPUCLK.power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X59_Y39_N18
cycloneive_lcell_comb \ramstore~0 (
// Equation(s):
// \ramstore~0_combout  = (\syif.tbCTRL~input_o  & (\syif.store[0]~input_o )) # (!\syif.tbCTRL~input_o  & ((plif_exmemrdat2_l_0)))

	.dataa(\syif.store[0]~input_o ),
	.datab(\syif.tbCTRL~input_o ),
	.datac(gnd),
	.datad(\CPU|DP|EXMEM|plif_exmem.rdat2_l [0]),
	.cin(gnd),
	.combout(\ramstore~0_combout ),
	.cout());
// synopsys translate_off
defparam \ramstore~0 .lut_mask = 16'hBB88;
defparam \ramstore~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X49_Y34_N2
cycloneive_lcell_comb \ramaddr~62 (
// Equation(s):
// \ramaddr~62_combout  = (\syif.tbCTRL~input_o  & (\syif.addr[1]~input_o )) # (!\syif.tbCTRL~input_o  & ((\ramaddr~0_combout )))

	.dataa(\syif.addr[1]~input_o ),
	.datab(\syif.tbCTRL~input_o ),
	.datac(gnd),
	.datad(\ramaddr~0_combout ),
	.cin(gnd),
	.combout(\ramaddr~62_combout ),
	.cout());
// synopsys translate_off
defparam \ramaddr~62 .lut_mask = 16'hBB88;
defparam \ramaddr~62 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X49_Y34_N14
cycloneive_lcell_comb \ramaddr~63 (
// Equation(s):
// \ramaddr~63_combout  = (\syif.tbCTRL~input_o  & (\syif.addr[0]~input_o )) # (!\syif.tbCTRL~input_o  & ((\ramaddr~1_combout )))

	.dataa(\syif.tbCTRL~input_o ),
	.datab(\syif.addr[0]~input_o ),
	.datac(\ramaddr~1_combout ),
	.datad(gnd),
	.cin(gnd),
	.combout(\ramaddr~63_combout ),
	.cout());
// synopsys translate_off
defparam \ramaddr~63 .lut_mask = 16'hD8D8;
defparam \ramaddr~63 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y25_N12
cycloneive_lcell_comb \ramstore~1 (
// Equation(s):
// \ramstore~1_combout  = (\syif.tbCTRL~input_o  & (\syif.store[1]~input_o )) # (!\syif.tbCTRL~input_o  & ((plif_exmemrdat2_l_1)))

	.dataa(\syif.tbCTRL~input_o ),
	.datab(gnd),
	.datac(\syif.store[1]~input_o ),
	.datad(\CPU|DP|EXMEM|plif_exmem.rdat2_l [1]),
	.cin(gnd),
	.combout(\ramstore~1_combout ),
	.cout());
// synopsys translate_off
defparam \ramstore~1 .lut_mask = 16'hF5A0;
defparam \ramstore~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y39_N4
cycloneive_lcell_comb \ramstore~2 (
// Equation(s):
// \ramstore~2_combout  = (\syif.tbCTRL~input_o  & ((\syif.store[2]~input_o ))) # (!\syif.tbCTRL~input_o  & (plif_exmemrdat2_l_2))

	.dataa(\CPU|DP|EXMEM|plif_exmem.rdat2_l [2]),
	.datab(\syif.store[2]~input_o ),
	.datac(gnd),
	.datad(\syif.tbCTRL~input_o ),
	.cin(gnd),
	.combout(\ramstore~2_combout ),
	.cout());
// synopsys translate_off
defparam \ramstore~2 .lut_mask = 16'hCCAA;
defparam \ramstore~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X52_Y34_N28
cycloneive_lcell_comb \ramstore~3 (
// Equation(s):
// \ramstore~3_combout  = (\syif.tbCTRL~input_o  & (\syif.store[3]~input_o )) # (!\syif.tbCTRL~input_o  & ((plif_exmemrdat2_l_3)))

	.dataa(\syif.store[3]~input_o ),
	.datab(\syif.tbCTRL~input_o ),
	.datac(gnd),
	.datad(\CPU|DP|EXMEM|plif_exmem.rdat2_l [3]),
	.cin(gnd),
	.combout(\ramstore~3_combout ),
	.cout());
// synopsys translate_off
defparam \ramstore~3 .lut_mask = 16'hBB88;
defparam \ramstore~3 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y34_N26
cycloneive_lcell_comb \ramstore~4 (
// Equation(s):
// \ramstore~4_combout  = (\syif.tbCTRL~input_o  & (\syif.store[4]~input_o )) # (!\syif.tbCTRL~input_o  & ((plif_exmemrdat2_l_4)))

	.dataa(\syif.tbCTRL~input_o ),
	.datab(gnd),
	.datac(\syif.store[4]~input_o ),
	.datad(\CPU|DP|EXMEM|plif_exmem.rdat2_l [4]),
	.cin(gnd),
	.combout(\ramstore~4_combout ),
	.cout());
// synopsys translate_off
defparam \ramstore~4 .lut_mask = 16'hF5A0;
defparam \ramstore~4 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y39_N8
cycloneive_lcell_comb \ramstore~5 (
// Equation(s):
// \ramstore~5_combout  = (\syif.tbCTRL~input_o  & (\syif.store[5]~input_o )) # (!\syif.tbCTRL~input_o  & ((plif_exmemrdat2_l_5)))

	.dataa(\syif.store[5]~input_o ),
	.datab(\syif.tbCTRL~input_o ),
	.datac(gnd),
	.datad(\CPU|DP|EXMEM|plif_exmem.rdat2_l [5]),
	.cin(gnd),
	.combout(\ramstore~5_combout ),
	.cout());
// synopsys translate_off
defparam \ramstore~5 .lut_mask = 16'hBB88;
defparam \ramstore~5 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y29_N26
cycloneive_lcell_comb \ramstore~6 (
// Equation(s):
// \ramstore~6_combout  = (\syif.tbCTRL~input_o  & (\syif.store[6]~input_o )) # (!\syif.tbCTRL~input_o  & ((plif_exmemrdat2_l_6)))

	.dataa(\syif.tbCTRL~input_o ),
	.datab(gnd),
	.datac(\syif.store[6]~input_o ),
	.datad(\CPU|DP|EXMEM|plif_exmem.rdat2_l [6]),
	.cin(gnd),
	.combout(\ramstore~6_combout ),
	.cout());
// synopsys translate_off
defparam \ramstore~6 .lut_mask = 16'hF5A0;
defparam \ramstore~6 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y34_N22
cycloneive_lcell_comb \ramstore~7 (
// Equation(s):
// \ramstore~7_combout  = (\syif.tbCTRL~input_o  & (\syif.store[7]~input_o )) # (!\syif.tbCTRL~input_o  & ((plif_exmemrdat2_l_7)))

	.dataa(\syif.store[7]~input_o ),
	.datab(gnd),
	.datac(\syif.tbCTRL~input_o ),
	.datad(\CPU|DP|EXMEM|plif_exmem.rdat2_l [7]),
	.cin(gnd),
	.combout(\ramstore~7_combout ),
	.cout());
// synopsys translate_off
defparam \ramstore~7 .lut_mask = 16'hAFA0;
defparam \ramstore~7 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X49_Y34_N26
cycloneive_lcell_comb \ramstore~8 (
// Equation(s):
// \ramstore~8_combout  = (\syif.tbCTRL~input_o  & (\syif.store[8]~input_o )) # (!\syif.tbCTRL~input_o  & ((plif_exmemrdat2_l_8)))

	.dataa(\syif.store[8]~input_o ),
	.datab(\syif.tbCTRL~input_o ),
	.datac(gnd),
	.datad(\CPU|DP|EXMEM|plif_exmem.rdat2_l [8]),
	.cin(gnd),
	.combout(\ramstore~8_combout ),
	.cout());
// synopsys translate_off
defparam \ramstore~8 .lut_mask = 16'hBB88;
defparam \ramstore~8 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y35_N30
cycloneive_lcell_comb \ramstore~9 (
// Equation(s):
// \ramstore~9_combout  = (\syif.tbCTRL~input_o  & (\syif.store[9]~input_o )) # (!\syif.tbCTRL~input_o  & ((plif_exmemrdat2_l_9)))

	.dataa(\syif.store[9]~input_o ),
	.datab(\syif.tbCTRL~input_o ),
	.datac(gnd),
	.datad(\CPU|DP|EXMEM|plif_exmem.rdat2_l [9]),
	.cin(gnd),
	.combout(\ramstore~9_combout ),
	.cout());
// synopsys translate_off
defparam \ramstore~9 .lut_mask = 16'hBB88;
defparam \ramstore~9 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X52_Y34_N8
cycloneive_lcell_comb \ramstore~10 (
// Equation(s):
// \ramstore~10_combout  = (\syif.tbCTRL~input_o  & (\syif.store[10]~input_o )) # (!\syif.tbCTRL~input_o  & ((plif_exmemrdat2_l_10)))

	.dataa(\syif.tbCTRL~input_o ),
	.datab(gnd),
	.datac(\syif.store[10]~input_o ),
	.datad(\CPU|DP|EXMEM|plif_exmem.rdat2_l [10]),
	.cin(gnd),
	.combout(\ramstore~10_combout ),
	.cout());
// synopsys translate_off
defparam \ramstore~10 .lut_mask = 16'hF5A0;
defparam \ramstore~10 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X63_Y27_N16
cycloneive_lcell_comb \ramstore~11 (
// Equation(s):
// \ramstore~11_combout  = (\syif.tbCTRL~input_o  & (\syif.store[11]~input_o )) # (!\syif.tbCTRL~input_o  & ((plif_exmemrdat2_l_11)))

	.dataa(gnd),
	.datab(\syif.store[11]~input_o ),
	.datac(\syif.tbCTRL~input_o ),
	.datad(\CPU|DP|EXMEM|plif_exmem.rdat2_l [11]),
	.cin(gnd),
	.combout(\ramstore~11_combout ),
	.cout());
// synopsys translate_off
defparam \ramstore~11 .lut_mask = 16'hCFC0;
defparam \ramstore~11 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y34_N8
cycloneive_lcell_comb \ramstore~12 (
// Equation(s):
// \ramstore~12_combout  = (\syif.tbCTRL~input_o  & (\syif.store[12]~input_o )) # (!\syif.tbCTRL~input_o  & ((plif_exmemrdat2_l_12)))

	.dataa(\syif.store[12]~input_o ),
	.datab(gnd),
	.datac(\syif.tbCTRL~input_o ),
	.datad(\CPU|DP|EXMEM|plif_exmem.rdat2_l [12]),
	.cin(gnd),
	.combout(\ramstore~12_combout ),
	.cout());
// synopsys translate_off
defparam \ramstore~12 .lut_mask = 16'hAFA0;
defparam \ramstore~12 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y39_N24
cycloneive_lcell_comb \ramstore~13 (
// Equation(s):
// \ramstore~13_combout  = (\syif.tbCTRL~input_o  & ((\syif.store[13]~input_o ))) # (!\syif.tbCTRL~input_o  & (plif_exmemrdat2_l_13))

	.dataa(\CPU|DP|EXMEM|plif_exmem.rdat2_l [13]),
	.datab(\syif.store[13]~input_o ),
	.datac(gnd),
	.datad(\syif.tbCTRL~input_o ),
	.cin(gnd),
	.combout(\ramstore~13_combout ),
	.cout());
// synopsys translate_off
defparam \ramstore~13 .lut_mask = 16'hCCAA;
defparam \ramstore~13 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y35_N12
cycloneive_lcell_comb \ramstore~14 (
// Equation(s):
// \ramstore~14_combout  = (\syif.tbCTRL~input_o  & ((\syif.store[14]~input_o ))) # (!\syif.tbCTRL~input_o  & (plif_exmemrdat2_l_14))

	.dataa(\syif.tbCTRL~input_o ),
	.datab(\CPU|DP|EXMEM|plif_exmem.rdat2_l [14]),
	.datac(gnd),
	.datad(\syif.store[14]~input_o ),
	.cin(gnd),
	.combout(\ramstore~14_combout ),
	.cout());
// synopsys translate_off
defparam \ramstore~14 .lut_mask = 16'hEE44;
defparam \ramstore~14 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X49_Y35_N28
cycloneive_lcell_comb \ramstore~15 (
// Equation(s):
// \ramstore~15_combout  = (\syif.tbCTRL~input_o  & ((\syif.store[15]~input_o ))) # (!\syif.tbCTRL~input_o  & (plif_exmemrdat2_l_15))

	.dataa(\CPU|DP|EXMEM|plif_exmem.rdat2_l [15]),
	.datab(\syif.store[15]~input_o ),
	.datac(gnd),
	.datad(\syif.tbCTRL~input_o ),
	.cin(gnd),
	.combout(\ramstore~15_combout ),
	.cout());
// synopsys translate_off
defparam \ramstore~15 .lut_mask = 16'hCCAA;
defparam \ramstore~15 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X49_Y30_N12
cycloneive_lcell_comb \ramstore~16 (
// Equation(s):
// \ramstore~16_combout  = (\syif.tbCTRL~input_o  & ((\syif.store[16]~input_o ))) # (!\syif.tbCTRL~input_o  & (plif_exmemrdat2_l_16))

	.dataa(\syif.tbCTRL~input_o ),
	.datab(gnd),
	.datac(\CPU|DP|EXMEM|plif_exmem.rdat2_l [16]),
	.datad(\syif.store[16]~input_o ),
	.cin(gnd),
	.combout(\ramstore~16_combout ),
	.cout());
// synopsys translate_off
defparam \ramstore~16 .lut_mask = 16'hFA50;
defparam \ramstore~16 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y39_N12
cycloneive_lcell_comb \ramstore~17 (
// Equation(s):
// \ramstore~17_combout  = (\syif.tbCTRL~input_o  & (\syif.store[17]~input_o )) # (!\syif.tbCTRL~input_o  & ((plif_exmemrdat2_l_17)))

	.dataa(gnd),
	.datab(\syif.store[17]~input_o ),
	.datac(\syif.tbCTRL~input_o ),
	.datad(\CPU|DP|EXMEM|plif_exmem.rdat2_l [17]),
	.cin(gnd),
	.combout(\ramstore~17_combout ),
	.cout());
// synopsys translate_off
defparam \ramstore~17 .lut_mask = 16'hCFC0;
defparam \ramstore~17 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y24_N12
cycloneive_lcell_comb \ramstore~18 (
// Equation(s):
// \ramstore~18_combout  = (\syif.tbCTRL~input_o  & (\syif.store[18]~input_o )) # (!\syif.tbCTRL~input_o  & ((plif_exmemrdat2_l_18)))

	.dataa(gnd),
	.datab(\syif.tbCTRL~input_o ),
	.datac(\syif.store[18]~input_o ),
	.datad(\CPU|DP|EXMEM|plif_exmem.rdat2_l [18]),
	.cin(gnd),
	.combout(\ramstore~18_combout ),
	.cout());
// synopsys translate_off
defparam \ramstore~18 .lut_mask = 16'hF3C0;
defparam \ramstore~18 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y34_N6
cycloneive_lcell_comb \ramstore~19 (
// Equation(s):
// \ramstore~19_combout  = (\syif.tbCTRL~input_o  & (\syif.store[19]~input_o )) # (!\syif.tbCTRL~input_o  & ((plif_exmemrdat2_l_19)))

	.dataa(gnd),
	.datab(\syif.store[19]~input_o ),
	.datac(\syif.tbCTRL~input_o ),
	.datad(\CPU|DP|EXMEM|plif_exmem.rdat2_l [19]),
	.cin(gnd),
	.combout(\ramstore~19_combout ),
	.cout());
// synopsys translate_off
defparam \ramstore~19 .lut_mask = 16'hCFC0;
defparam \ramstore~19 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y35_N20
cycloneive_lcell_comb \ramstore~20 (
// Equation(s):
// \ramstore~20_combout  = (\syif.tbCTRL~input_o  & (\syif.store[20]~input_o )) # (!\syif.tbCTRL~input_o  & ((plif_exmemrdat2_l_20)))

	.dataa(\syif.store[20]~input_o ),
	.datab(\syif.tbCTRL~input_o ),
	.datac(gnd),
	.datad(\CPU|DP|EXMEM|plif_exmem.rdat2_l [20]),
	.cin(gnd),
	.combout(\ramstore~20_combout ),
	.cout());
// synopsys translate_off
defparam \ramstore~20 .lut_mask = 16'hBB88;
defparam \ramstore~20 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y32_N26
cycloneive_lcell_comb \ramstore~21 (
// Equation(s):
// \ramstore~21_combout  = (\syif.tbCTRL~input_o  & (\syif.store[21]~input_o )) # (!\syif.tbCTRL~input_o  & ((plif_exmemrdat2_l_21)))

	.dataa(\syif.tbCTRL~input_o ),
	.datab(\syif.store[21]~input_o ),
	.datac(gnd),
	.datad(\CPU|DP|EXMEM|plif_exmem.rdat2_l [21]),
	.cin(gnd),
	.combout(\ramstore~21_combout ),
	.cout());
// synopsys translate_off
defparam \ramstore~21 .lut_mask = 16'hDD88;
defparam \ramstore~21 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y39_N30
cycloneive_lcell_comb \ramstore~22 (
// Equation(s):
// \ramstore~22_combout  = (\syif.tbCTRL~input_o  & (\syif.store[22]~input_o )) # (!\syif.tbCTRL~input_o  & ((plif_exmemrdat2_l_22)))

	.dataa(\syif.store[22]~input_o ),
	.datab(\syif.tbCTRL~input_o ),
	.datac(gnd),
	.datad(\CPU|DP|EXMEM|plif_exmem.rdat2_l [22]),
	.cin(gnd),
	.combout(\ramstore~22_combout ),
	.cout());
// synopsys translate_off
defparam \ramstore~22 .lut_mask = 16'hBB88;
defparam \ramstore~22 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X52_Y23_N0
cycloneive_lcell_comb \ramstore~23 (
// Equation(s):
// \ramstore~23_combout  = (\syif.tbCTRL~input_o  & (\syif.store[23]~input_o )) # (!\syif.tbCTRL~input_o  & ((plif_exmemrdat2_l_23)))

	.dataa(\syif.tbCTRL~input_o ),
	.datab(\syif.store[23]~input_o ),
	.datac(gnd),
	.datad(\CPU|DP|EXMEM|plif_exmem.rdat2_l [23]),
	.cin(gnd),
	.combout(\ramstore~23_combout ),
	.cout());
// synopsys translate_off
defparam \ramstore~23 .lut_mask = 16'hDD88;
defparam \ramstore~23 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y29_N8
cycloneive_lcell_comb \ramstore~24 (
// Equation(s):
// \ramstore~24_combout  = (\syif.tbCTRL~input_o  & (\syif.store[24]~input_o )) # (!\syif.tbCTRL~input_o  & ((plif_exmemrdat2_l_24)))

	.dataa(\syif.store[24]~input_o ),
	.datab(gnd),
	.datac(\syif.tbCTRL~input_o ),
	.datad(\CPU|DP|EXMEM|plif_exmem.rdat2_l [24]),
	.cin(gnd),
	.combout(\ramstore~24_combout ),
	.cout());
// synopsys translate_off
defparam \ramstore~24 .lut_mask = 16'hAFA0;
defparam \ramstore~24 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y32_N14
cycloneive_lcell_comb \ramstore~25 (
// Equation(s):
// \ramstore~25_combout  = (\syif.tbCTRL~input_o  & (\syif.store[25]~input_o )) # (!\syif.tbCTRL~input_o  & ((plif_exmemrdat2_l_25)))

	.dataa(\syif.tbCTRL~input_o ),
	.datab(gnd),
	.datac(\syif.store[25]~input_o ),
	.datad(\CPU|DP|EXMEM|plif_exmem.rdat2_l [25]),
	.cin(gnd),
	.combout(\ramstore~25_combout ),
	.cout());
// synopsys translate_off
defparam \ramstore~25 .lut_mask = 16'hF5A0;
defparam \ramstore~25 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y29_N2
cycloneive_lcell_comb \ramstore~26 (
// Equation(s):
// \ramstore~26_combout  = (\syif.tbCTRL~input_o  & (\syif.store[26]~input_o )) # (!\syif.tbCTRL~input_o  & ((plif_exmemrdat2_l_26)))

	.dataa(\syif.store[26]~input_o ),
	.datab(\CPU|DP|EXMEM|plif_exmem.rdat2_l [26]),
	.datac(\syif.tbCTRL~input_o ),
	.datad(gnd),
	.cin(gnd),
	.combout(\ramstore~26_combout ),
	.cout());
// synopsys translate_off
defparam \ramstore~26 .lut_mask = 16'hACAC;
defparam \ramstore~26 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X50_Y36_N4
cycloneive_lcell_comb \ramstore~27 (
// Equation(s):
// \ramstore~27_combout  = (\syif.tbCTRL~input_o  & (\syif.store[27]~input_o )) # (!\syif.tbCTRL~input_o  & ((plif_exmemrdat2_l_27)))

	.dataa(gnd),
	.datab(\syif.store[27]~input_o ),
	.datac(\syif.tbCTRL~input_o ),
	.datad(\CPU|DP|EXMEM|plif_exmem.rdat2_l [27]),
	.cin(gnd),
	.combout(\ramstore~27_combout ),
	.cout());
// synopsys translate_off
defparam \ramstore~27 .lut_mask = 16'hCFC0;
defparam \ramstore~27 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y35_N8
cycloneive_lcell_comb \ramstore~28 (
// Equation(s):
// \ramstore~28_combout  = (\syif.tbCTRL~input_o  & (\syif.store[28]~input_o )) # (!\syif.tbCTRL~input_o  & ((plif_exmemrdat2_l_28)))

	.dataa(\syif.store[28]~input_o ),
	.datab(\syif.tbCTRL~input_o ),
	.datac(gnd),
	.datad(\CPU|DP|EXMEM|plif_exmem.rdat2_l [28]),
	.cin(gnd),
	.combout(\ramstore~28_combout ),
	.cout());
// synopsys translate_off
defparam \ramstore~28 .lut_mask = 16'hBB88;
defparam \ramstore~28 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y34_N16
cycloneive_lcell_comb \ramstore~29 (
// Equation(s):
// \ramstore~29_combout  = (\syif.tbCTRL~input_o  & (\syif.store[29]~input_o )) # (!\syif.tbCTRL~input_o  & ((plif_exmemrdat2_l_29)))

	.dataa(\syif.tbCTRL~input_o ),
	.datab(\syif.store[29]~input_o ),
	.datac(gnd),
	.datad(\CPU|DP|EXMEM|plif_exmem.rdat2_l [29]),
	.cin(gnd),
	.combout(\ramstore~29_combout ),
	.cout());
// synopsys translate_off
defparam \ramstore~29 .lut_mask = 16'hDD88;
defparam \ramstore~29 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y32_N0
cycloneive_lcell_comb \ramstore~30 (
// Equation(s):
// \ramstore~30_combout  = (\syif.tbCTRL~input_o  & (\syif.store[30]~input_o )) # (!\syif.tbCTRL~input_o  & ((plif_exmemrdat2_l_30)))

	.dataa(\syif.tbCTRL~input_o ),
	.datab(gnd),
	.datac(\syif.store[30]~input_o ),
	.datad(\CPU|DP|EXMEM|plif_exmem.rdat2_l [30]),
	.cin(gnd),
	.combout(\ramstore~30_combout ),
	.cout());
// synopsys translate_off
defparam \ramstore~30 .lut_mask = 16'hF5A0;
defparam \ramstore~30 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y26_N20
cycloneive_lcell_comb \ramstore~31 (
// Equation(s):
// \ramstore~31_combout  = (\syif.tbCTRL~input_o  & (\syif.store[31]~input_o )) # (!\syif.tbCTRL~input_o  & ((plif_exmemrdat2_l_31)))

	.dataa(gnd),
	.datab(\syif.tbCTRL~input_o ),
	.datac(\syif.store[31]~input_o ),
	.datad(\CPU|DP|EXMEM|plif_exmem.rdat2_l [31]),
	.cin(gnd),
	.combout(\ramstore~31_combout ),
	.cout());
// synopsys translate_off
defparam \ramstore~31 .lut_mask = 16'hF3C0;
defparam \ramstore~31 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X59_Y1_N9
dffeas \count[3] (
	.clk(\CLK~inputclkctrl_outclk ),
	.d(\count[3]~0_combout ),
	.asdata(vcc),
	.clrn(\nRST~inputclkctrl_outclk ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(count[3]),
	.prn(vcc));
// synopsys translate_off
defparam \count[3] .is_wysiwyg = "true";
defparam \count[3] .power_up = "low";
// synopsys translate_on

// Location: FF_X59_Y1_N11
dffeas \count[2] (
	.clk(\CLK~inputclkctrl_outclk ),
	.d(\count[2]~1_combout ),
	.asdata(vcc),
	.clrn(\nRST~inputclkctrl_outclk ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(count[2]),
	.prn(vcc));
// synopsys translate_off
defparam \count[2] .is_wysiwyg = "true";
defparam \count[2] .power_up = "low";
// synopsys translate_on

// Location: FF_X59_Y1_N5
dffeas \count[1] (
	.clk(\CLK~inputclkctrl_outclk ),
	.d(\count[1]~2_combout ),
	.asdata(vcc),
	.clrn(\nRST~inputclkctrl_outclk ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(count[1]),
	.prn(vcc));
// synopsys translate_off
defparam \count[1] .is_wysiwyg = "true";
defparam \count[1] .power_up = "low";
// synopsys translate_on

// Location: FF_X59_Y1_N1
dffeas \count[0] (
	.clk(\CLK~inputclkctrl_outclk ),
	.d(\count~3_combout ),
	.asdata(vcc),
	.clrn(\nRST~inputclkctrl_outclk ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(count[0]),
	.prn(vcc));
// synopsys translate_off
defparam \count[0] .is_wysiwyg = "true";
defparam \count[0] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X59_Y1_N12
cycloneive_lcell_comb \Equal0~0 (
// Equation(s):
// \Equal0~0_combout  = (!count[2] & (!count[1] & (!count[3] & !count[0])))

	.dataa(count[2]),
	.datab(count[1]),
	.datac(count[3]),
	.datad(count[0]),
	.cin(gnd),
	.combout(\Equal0~0_combout ),
	.cout());
// synopsys translate_off
defparam \Equal0~0 .lut_mask = 16'h0001;
defparam \Equal0~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y1_N24
cycloneive_lcell_comb \CPUCLK~0 (
// Equation(s):
// \CPUCLK~0_combout  = \CPUCLK~q  $ (\Equal0~0_combout )

	.dataa(gnd),
	.datab(gnd),
	.datac(\CPUCLK~q ),
	.datad(\Equal0~0_combout ),
	.cin(gnd),
	.combout(\CPUCLK~0_combout ),
	.cout());
// synopsys translate_off
defparam \CPUCLK~0 .lut_mask = 16'h0FF0;
defparam \CPUCLK~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y1_N8
cycloneive_lcell_comb \count[3]~0 (
// Equation(s):
// \count[3]~0_combout  = count[3] $ (((count[2] & (count[1] & count[0]))))

	.dataa(count[2]),
	.datab(count[1]),
	.datac(count[3]),
	.datad(count[0]),
	.cin(gnd),
	.combout(\count[3]~0_combout ),
	.cout());
// synopsys translate_off
defparam \count[3]~0 .lut_mask = 16'h78F0;
defparam \count[3]~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y1_N10
cycloneive_lcell_comb \count[2]~1 (
// Equation(s):
// \count[2]~1_combout  = count[2] $ (((count[1] & count[0])))

	.dataa(gnd),
	.datab(count[1]),
	.datac(count[2]),
	.datad(count[0]),
	.cin(gnd),
	.combout(\count[2]~1_combout ),
	.cout());
// synopsys translate_off
defparam \count[2]~1 .lut_mask = 16'h3CF0;
defparam \count[2]~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y1_N4
cycloneive_lcell_comb \count[1]~2 (
// Equation(s):
// \count[1]~2_combout  = count[1] $ (count[0])

	.dataa(gnd),
	.datab(gnd),
	.datac(count[1]),
	.datad(count[0]),
	.cin(gnd),
	.combout(\count[1]~2_combout ),
	.cout());
// synopsys translate_off
defparam \count[1]~2 .lut_mask = 16'h0FF0;
defparam \count[1]~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y1_N0
cycloneive_lcell_comb \count~3 (
// Equation(s):
// \count~3_combout  = (!count[0] & ((count[2]) # ((count[1]) # (count[3]))))

	.dataa(count[2]),
	.datab(count[1]),
	.datac(count[0]),
	.datad(count[3]),
	.cin(gnd),
	.combout(\count~3_combout ),
	.cout());
// synopsys translate_off
defparam \count~3 .lut_mask = 16'h0F0E;
defparam \count~3 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y34_N20
cycloneive_lcell_comb \ramaddr~27_wirecell (
// Equation(s):
// \ramaddr~27_wirecell_combout  = !\ramaddr~27_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(\ramaddr~27_combout ),
	.datad(gnd),
	.cin(gnd),
	.combout(\ramaddr~27_wirecell_combout ),
	.cout());
// synopsys translate_off
defparam \ramaddr~27_wirecell .lut_mask = 16'h0F0F;
defparam \ramaddr~27_wirecell .sum_lutc_input = "datac";
// synopsys translate_on

// Location: JTAG_X1_Y37_N0
cycloneive_jtag altera_internal_jtag(
	.tms(\altera_reserved_tms~input_o ),
	.tck(\altera_reserved_tck~input_o ),
	.tdi(\altera_reserved_tdi~input_o ),
	.tdoutap(gnd),
	.tdouser(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|tdo~_wirecell_combout ),
	.tdo(\altera_internal_jtag~TDO ),
	.tmsutap(\altera_internal_jtag~TMSUTAP ),
	.tckutap(\altera_internal_jtag~TCKUTAP ),
	.tdiutap(\altera_internal_jtag~TDIUTAP ),
	.shiftuser(),
	.clkdruser(),
	.updateuser(),
	.runidleuser(),
	.usr1user());

// Location: FF_X42_Y33_N7
dffeas \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter[2] (
	.clk(\altera_internal_jtag~TCKUTAPclkctrl_outclk ),
	.d(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter[2]~15_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter[1]~22_combout ),
	.sload(gnd),
	.ena(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter[1]~23_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter [2]),
	.prn(vcc));
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter[2] .is_wysiwyg = "true";
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter[2] .power_up = "low";
// synopsys translate_on

// Location: FF_X42_Y33_N3
dffeas \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter[0] (
	.clk(\altera_internal_jtag~TCKUTAPclkctrl_outclk ),
	.d(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter[0]~11_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter[1]~22_combout ),
	.sload(gnd),
	.ena(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter[1]~23_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter [0]),
	.prn(vcc));
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter[0] .is_wysiwyg = "true";
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter[0] .power_up = "low";
// synopsys translate_on

// Location: FF_X42_Y33_N9
dffeas \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter[3] (
	.clk(\altera_internal_jtag~TCKUTAPclkctrl_outclk ),
	.d(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter[3]~18_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter[1]~22_combout ),
	.sload(gnd),
	.ena(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter[1]~23_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter [3]),
	.prn(vcc));
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter[3] .is_wysiwyg = "true";
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter[3] .power_up = "low";
// synopsys translate_on

// Location: FF_X42_Y33_N11
dffeas \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter[4] (
	.clk(\altera_internal_jtag~TCKUTAPclkctrl_outclk ),
	.d(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter[4]~20_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter[1]~22_combout ),
	.sload(gnd),
	.ena(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter[1]~23_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter [4]),
	.prn(vcc));
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter[4] .is_wysiwyg = "true";
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter[4] .power_up = "low";
// synopsys translate_on

// Location: FF_X42_Y33_N5
dffeas \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter[1] (
	.clk(\altera_internal_jtag~TCKUTAPclkctrl_outclk ),
	.d(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter[1]~13_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter[1]~22_combout ),
	.sload(gnd),
	.ena(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter[1]~23_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter [1]),
	.prn(vcc));
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter[1] .is_wysiwyg = "true";
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter[1] .power_up = "low";
// synopsys translate_on

// Location: FF_X45_Y33_N7
dffeas \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|tms_cnt[1] (
	.clk(\altera_internal_jtag~TCKUTAPclkctrl_outclk ),
	.d(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|tms_cnt~2_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!\altera_internal_jtag~TMSUTAP ),
	.sload(gnd),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|tms_cnt [1]),
	.prn(vcc));
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|tms_cnt[1] .is_wysiwyg = "true";
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|tms_cnt[1] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X42_Y33_N2
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter[0]~11 (
	.dataa(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter [0]),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(gnd),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter[0]~11_combout ),
	.cout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter[0]~12 ));
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter[0]~11 .lut_mask = 16'h55AA;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter[0]~11 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X42_Y33_N4
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter[1]~13 (
	.dataa(gnd),
	.datab(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter [1]),
	.datac(gnd),
	.datad(vcc),
	.cin(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter[0]~12 ),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter[1]~13_combout ),
	.cout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter[1]~14 ));
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter[1]~13 .lut_mask = 16'h3C3F;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter[1]~13 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X42_Y33_N6
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter[2]~15 (
	.dataa(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter [2]),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter[1]~14 ),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter[2]~15_combout ),
	.cout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter[2]~16 ));
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter[2]~15 .lut_mask = 16'hA50A;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter[2]~15 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X42_Y33_N8
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter[3]~18 (
	.dataa(gnd),
	.datab(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter [3]),
	.datac(gnd),
	.datad(vcc),
	.cin(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter[2]~16 ),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter[3]~18_combout ),
	.cout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter[3]~19 ));
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter[3]~18 .lut_mask = 16'h3C3F;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter[3]~18 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X42_Y33_N10
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter[4]~20 (
	.dataa(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter [4]),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.cin(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter[3]~19 ),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter[4]~20_combout ),
	.cout());
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter[4]~20 .lut_mask = 16'hA5A5;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter[4]~20 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: FF_X46_Y33_N13
dffeas \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irf_reg[1][0] (
	.clk(\altera_internal_jtag~TCKUTAPclkctrl_outclk ),
	.d(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irf_reg[1][0]~feeder_combout ),
	.asdata(vcc),
	.clrn(!\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|clr_reg~q ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irf_reg[1][0]~0_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irf_reg[1][0]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irf_reg[1][0] .is_wysiwyg = "true";
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irf_reg[1][0] .power_up = "low";
// synopsys translate_on

// Location: FF_X46_Y33_N11
dffeas \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irf_reg[1][1] (
	.clk(\altera_internal_jtag~TCKUTAPclkctrl_outclk ),
	.d(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irf_reg[1][1]~feeder_combout ),
	.asdata(vcc),
	.clrn(!\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|clr_reg~q ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irf_reg[1][0]~0_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irf_reg[1][1]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irf_reg[1][1] .is_wysiwyg = "true";
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irf_reg[1][1] .power_up = "low";
// synopsys translate_on

// Location: FF_X46_Y33_N1
dffeas \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irf_reg[1][2] (
	.clk(\altera_internal_jtag~TCKUTAPclkctrl_outclk ),
	.d(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irf_reg[1][2]~feeder_combout ),
	.asdata(vcc),
	.clrn(!\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|clr_reg~q ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irf_reg[1][0]~0_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irf_reg[1][2]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irf_reg[1][2] .is_wysiwyg = "true";
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irf_reg[1][2] .power_up = "low";
// synopsys translate_on

// Location: FF_X46_Y33_N23
dffeas \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irf_reg[1][3] (
	.clk(\altera_internal_jtag~TCKUTAPclkctrl_outclk ),
	.d(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irf_reg[1][3]~feeder_combout ),
	.asdata(vcc),
	.clrn(!\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|clr_reg~q ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irf_reg[1][0]~0_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irf_reg[1][3]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irf_reg[1][3] .is_wysiwyg = "true";
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irf_reg[1][3] .power_up = "low";
// synopsys translate_on

// Location: FF_X46_Y33_N29
dffeas \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irf_reg[1][4] (
	.clk(\altera_internal_jtag~TCKUTAPclkctrl_outclk ),
	.d(gnd),
	.asdata(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg [4]),
	.clrn(!\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|clr_reg~q ),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irf_reg[1][0]~0_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irf_reg[1][4]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irf_reg[1][4] .is_wysiwyg = "true";
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irf_reg[1][4] .power_up = "low";
// synopsys translate_on

// Location: FF_X45_Y33_N5
dffeas \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|node_ena[1]~reg0 (
	.clk(\altera_internal_jtag~TCKUTAPclkctrl_outclk ),
	.d(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|node_ena~3_combout ),
	.asdata(vcc),
	.clrn(!\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|clr_reg~q ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|node_ena[1]~reg0_q ),
	.prn(vcc));
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|node_ena[1]~reg0 .is_wysiwyg = "true";
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|node_ena[1]~reg0 .power_up = "low";
// synopsys translate_on

// Location: FF_X45_Y33_N17
dffeas \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_minor_ver_reg[0] (
	.clk(\altera_internal_jtag~TCKUTAPclkctrl_outclk ),
	.d(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_minor_ver_reg~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg_ena~0_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_minor_ver_reg [0]),
	.prn(vcc));
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_minor_ver_reg[0] .is_wysiwyg = "true";
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_minor_ver_reg[0] .power_up = "low";
// synopsys translate_on

// Location: FF_X42_Y33_N1
dffeas \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|WORD_SR[0] (
	.clk(\altera_internal_jtag~TCKUTAPclkctrl_outclk ),
	.d(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|WORD_SR~8_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|WORD_SR[1]~15_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|WORD_SR [0]),
	.prn(vcc));
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|WORD_SR[0] .is_wysiwyg = "true";
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|WORD_SR[0] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X46_Y33_N14
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|tdo~0 (
	.dataa(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_minor_ver_reg [0]),
	.datab(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg [0]),
	.datac(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|WORD_SR [0]),
	.datad(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg [2]),
	.cin(gnd),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|tdo~0_combout ),
	.cout());
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|tdo~0 .lut_mask = 16'hEE30;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|tdo~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X45_Y34_N12
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|reset_ena_reg_proc~0 (
	.dataa(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [7]),
	.datab(\altera_internal_jtag~TMSUTAP ),
	.datac(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [5]),
	.datad(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|virtual_ir_scan_reg~q ),
	.cin(gnd),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|reset_ena_reg_proc~0_combout ),
	.cout());
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|reset_ena_reg_proc~0 .lut_mask = 16'hC800;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|reset_ena_reg_proc~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X46_Y33_N18
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irf_reg[1][0]~0 (
	.dataa(gnd),
	.datab(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg [5]),
	.datac(gnd),
	.datad(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|reset_ena_reg_proc~0_combout ),
	.cin(gnd),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irf_reg[1][0]~0_combout ),
	.cout());
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irf_reg[1][0]~0 .lut_mask = 16'hCC00;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irf_reg[1][0]~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X43_Y33_N22
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|node_ena~0 (
	.dataa(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg [5]),
	.datab(\altera_internal_jtag~TDIUTAP ),
	.datac(\altera_internal_jtag~TMSUTAP ),
	.datad(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [4]),
	.cin(gnd),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|node_ena~0_combout ),
	.cout());
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|node_ena~0 .lut_mask = 16'hCAAA;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|node_ena~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X45_Y33_N26
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|node_ena~1 (
	.dataa(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|node_ena~0_combout ),
	.datab(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_mode_reg [1]),
	.datac(\altera_internal_jtag~TMSUTAP ),
	.datad(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [2]),
	.cin(gnd),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|node_ena~1_combout ),
	.cout());
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|node_ena~1 .lut_mask = 16'h0222;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|node_ena~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X43_Y33_N0
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|node_ena_proc~0 (
	.dataa(gnd),
	.datab(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [4]),
	.datac(\altera_internal_jtag~TMSUTAP ),
	.datad(gnd),
	.cin(gnd),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|node_ena_proc~0_combout ),
	.cout());
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|node_ena_proc~0 .lut_mask = 16'hC0C0;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|node_ena_proc~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X43_Y33_N26
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|node_ena~2 (
	.dataa(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [15]),
	.datab(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|node_ena_proc~0_combout ),
	.datac(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|virtual_ir_scan_reg~q ),
	.datad(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|virtual_dr_scan_reg~q ),
	.cin(gnd),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|node_ena~2_combout ),
	.cout());
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|node_ena~2 .lut_mask = 16'hE2E0;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|node_ena~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X45_Y33_N4
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|node_ena~3 (
	.dataa(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|node_ena~1_combout ),
	.datab(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|node_ena_proc~1_combout ),
	.datac(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|node_ena[1]~reg0_q ),
	.datad(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|node_ena~2_combout ),
	.cin(gnd),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|node_ena~3_combout ),
	.cout());
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|node_ena~3 .lut_mask = 16'hAA30;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|node_ena~3 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X43_Y34_N12
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|Equal0~0 (
	.dataa(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg [8]),
	.datab(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg [7]),
	.datac(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg [6]),
	.datad(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg [9]),
	.cin(gnd),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|Equal0~0_combout ),
	.cout());
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|Equal0~0 .lut_mask = 16'h0001;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|Equal0~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X40_Y33_N12
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg[3]~13 (
	.dataa(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg [2]),
	.datab(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg [0]),
	.datac(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg [3]),
	.datad(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg [1]),
	.cin(gnd),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg[3]~13_combout ),
	.cout());
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg[3]~13 .lut_mask = 16'h8000;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg[3]~13 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X45_Y32_N29
dffeas \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_mode_reg[0] (
	.clk(\altera_internal_jtag~TCKUTAPclkctrl_outclk ),
	.d(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_mode_reg[0]~4_combout ),
	.asdata(vcc),
	.clrn(!\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|clr_reg~q ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_mode_reg [0]),
	.prn(vcc));
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_mode_reg[0] .is_wysiwyg = "true";
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_mode_reg[0] .power_up = "low";
// synopsys translate_on

// Location: FF_X45_Y33_N15
dffeas \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_minor_ver_reg[1] (
	.clk(\altera_internal_jtag~TCKUTAPclkctrl_outclk ),
	.d(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_minor_ver_reg~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg_ena~0_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_minor_ver_reg [1]),
	.prn(vcc));
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_minor_ver_reg[1] .is_wysiwyg = "true";
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_minor_ver_reg[1] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X45_Y33_N16
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_minor_ver_reg~0 (
	.dataa(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [3]),
	.datab(gnd),
	.datac(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_minor_ver_reg [1]),
	.datad(gnd),
	.cin(gnd),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_minor_ver_reg~0_combout ),
	.cout());
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_minor_ver_reg~0 .lut_mask = 16'hFAFA;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_minor_ver_reg~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X42_Y33_N16
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|WORD_SR~6 (
	.dataa(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter [2]),
	.datab(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter [3]),
	.datac(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter [0]),
	.datad(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter [4]),
	.cin(gnd),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|WORD_SR~6_combout ),
	.cout());
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|WORD_SR~6 .lut_mask = 16'h8081;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|WORD_SR~6 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X42_Y33_N26
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|WORD_SR~7 (
	.dataa(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|clear_signal~combout ),
	.datab(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter [1]),
	.datac(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [4]),
	.datad(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|WORD_SR~6_combout ),
	.cin(gnd),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|WORD_SR~7_combout ),
	.cout());
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|WORD_SR~7 .lut_mask = 16'h0100;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|WORD_SR~7 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X42_Y33_N21
dffeas \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|WORD_SR[1] (
	.clk(\altera_internal_jtag~TCKUTAPclkctrl_outclk ),
	.d(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|WORD_SR~16_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|WORD_SR[1]~15_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|WORD_SR [1]),
	.prn(vcc));
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|WORD_SR[1] .is_wysiwyg = "true";
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|WORD_SR[1] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X42_Y33_N0
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|WORD_SR~8 (
	.dataa(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|clear_signal~combout ),
	.datab(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|WORD_SR [1]),
	.datac(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [4]),
	.datad(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|WORD_SR~7_combout ),
	.cin(gnd),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|WORD_SR~8_combout ),
	.cout());
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|WORD_SR~8 .lut_mask = 16'hFF40;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|WORD_SR~8 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X43_Y33_N10
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg~7 (
	.dataa(gnd),
	.datab(gnd),
	.datac(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_mode_reg [0]),
	.datad(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg [3]),
	.cin(gnd),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg~7_combout ),
	.cout());
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg~7 .lut_mask = 16'h0F00;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg~7 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X45_Y34_N13
dffeas \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|reset_ena_reg (
	.clk(\altera_internal_jtag~TCKUTAPclkctrl_outclk ),
	.d(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|reset_ena_reg_proc~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|reset_ena_reg~q ),
	.prn(vcc));
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|reset_ena_reg .is_wysiwyg = "true";
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|reset_ena_reg .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X40_Y33_N0
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg~15 (
	.dataa(gnd),
	.datab(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg [4]),
	.datac(gnd),
	.datad(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg [1]),
	.cin(gnd),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg~15_combout ),
	.cout());
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg~15 .lut_mask = 16'h0033;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg~15 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X48_Y33_N21
dffeas \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|identity_contrib_update_reg[1] (
	.clk(\altera_internal_jtag~TCKUTAPclkctrl_outclk ),
	.d(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|identity_contrib_update_reg[1]~feeder_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|identity_contrib_update_reg[0]~0_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|identity_contrib_update_reg [1]),
	.prn(vcc));
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|identity_contrib_update_reg[1] .is_wysiwyg = "true";
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|identity_contrib_update_reg[1] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X46_Y33_N30
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|Equal3~0 (
	.dataa(gnd),
	.datab(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg [0]),
	.datac(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg [2]),
	.datad(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg [1]),
	.cin(gnd),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|Equal3~0_combout ),
	.cout());
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|Equal3~0 .lut_mask = 16'h0C00;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|Equal3~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X45_Y32_N28
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_mode_reg[0]~4 (
	.dataa(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|Equal3~0_combout ),
	.datab(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg [5]),
	.datac(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_mode_reg [0]),
	.datad(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|reset_ena_reg_proc~0_combout ),
	.cin(gnd),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_mode_reg[0]~4_combout ),
	.cout());
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_mode_reg[0]~4 .lut_mask = 16'h22F0;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_mode_reg[0]~4 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X45_Y33_N19
dffeas \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_minor_ver_reg[2] (
	.clk(\altera_internal_jtag~TCKUTAPclkctrl_outclk ),
	.d(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_minor_ver_reg~2_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg_ena~0_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_minor_ver_reg [2]),
	.prn(vcc));
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_minor_ver_reg[2] .is_wysiwyg = "true";
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_minor_ver_reg[2] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X45_Y33_N14
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_minor_ver_reg~1 (
	.dataa(gnd),
	.datab(gnd),
	.datac(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [3]),
	.datad(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_minor_ver_reg [2]),
	.cin(gnd),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_minor_ver_reg~1_combout ),
	.cout());
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_minor_ver_reg~1 .lut_mask = 16'h0F00;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_minor_ver_reg~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X42_Y33_N14
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter[1]~17 (
	.dataa(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter [0]),
	.datab(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter [3]),
	.datac(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter [1]),
	.datad(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter [2]),
	.cin(gnd),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter[1]~17_combout ),
	.cout());
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter[1]~17 .lut_mask = 16'hFFFE;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter[1]~17 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X42_Y33_N25
dffeas \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|WORD_SR[2] (
	.clk(\altera_internal_jtag~TCKUTAPclkctrl_outclk ),
	.d(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|WORD_SR~12_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|WORD_SR[1]~15_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|WORD_SR [2]),
	.prn(vcc));
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|WORD_SR[2] .is_wysiwyg = "true";
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|WORD_SR[2] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X42_Y33_N22
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|WORD_SR~9 (
	.dataa(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter [2]),
	.datab(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter [1]),
	.datac(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [4]),
	.datad(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|WORD_SR [2]),
	.cin(gnd),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|WORD_SR~9_combout ),
	.cout());
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|WORD_SR~9 .lut_mask = 16'hF404;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|WORD_SR~9 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X45_Y33_N6
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|tms_cnt~2 (
	.dataa(gnd),
	.datab(gnd),
	.datac(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|tms_cnt [1]),
	.datad(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|tms_cnt [0]),
	.cin(gnd),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|tms_cnt~2_combout ),
	.cout());
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|tms_cnt~2 .lut_mask = 16'h0FF0;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|tms_cnt~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X41_Y33_N0
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg~16 (
	.dataa(gnd),
	.datab(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg [2]),
	.datac(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg [0]),
	.datad(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg [3]),
	.cin(gnd),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg~16_combout ),
	.cout());
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg~16 .lut_mask = 16'hFFCF;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg~16 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X40_Y33_N14
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg~17 (
	.dataa(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg [4]),
	.datab(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg [0]),
	.datac(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg [2]),
	.datad(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg [1]),
	.cin(gnd),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg~17_combout ),
	.cout());
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg~17 .lut_mask = 16'h4E08;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg~17 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X41_Y33_N2
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg~18 (
	.dataa(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg~17_combout ),
	.datab(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg [3]),
	.datac(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg~15_combout ),
	.datad(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg~16_combout ),
	.cin(gnd),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg~18_combout ),
	.cout());
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg~18 .lut_mask = 16'hF222;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg~18 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X45_Y33_N9
dffeas \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_minor_ver_reg[3] (
	.clk(\altera_internal_jtag~TCKUTAPclkctrl_outclk ),
	.d(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_minor_ver_reg~3_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg_ena~0_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_minor_ver_reg [3]),
	.prn(vcc));
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_minor_ver_reg[3] .is_wysiwyg = "true";
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_minor_ver_reg[3] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X45_Y33_N18
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_minor_ver_reg~2 (
	.dataa(gnd),
	.datab(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_minor_ver_reg [3]),
	.datac(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [3]),
	.datad(gnd),
	.cin(gnd),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_minor_ver_reg~2_combout ),
	.cout());
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_minor_ver_reg~2 .lut_mask = 16'hFCFC;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_minor_ver_reg~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X42_Y33_N28
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|WORD_SR~10 (
	.dataa(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter [0]),
	.datab(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter [3]),
	.datac(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter [1]),
	.datad(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter [4]),
	.cin(gnd),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|WORD_SR~10_combout ),
	.cout());
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|WORD_SR~10 .lut_mask = 16'hF0F1;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|WORD_SR~10 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X42_Y33_N18
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|WORD_SR~11 (
	.dataa(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|clear_signal~combout ),
	.datab(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|WORD_SR~10_combout ),
	.datac(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [4]),
	.datad(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter [2]),
	.cin(gnd),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|WORD_SR~11_combout ),
	.cout());
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|WORD_SR~11 .lut_mask = 16'h0004;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|WORD_SR~11 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X43_Y33_N7
dffeas \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|WORD_SR[3] (
	.clk(\altera_internal_jtag~TCKUTAPclkctrl_outclk ),
	.d(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|WORD_SR~14_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|WORD_SR[1]~15_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|WORD_SR [3]),
	.prn(vcc));
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|WORD_SR[3] .is_wysiwyg = "true";
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|WORD_SR[3] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X42_Y33_N24
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|WORD_SR~12 (
	.dataa(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|WORD_SR [3]),
	.datab(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [4]),
	.datac(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|clear_signal~combout ),
	.datad(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|WORD_SR~11_combout ),
	.cin(gnd),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|WORD_SR~12_combout ),
	.cout());
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|WORD_SR~12 .lut_mask = 16'hFF08;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|WORD_SR~12 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X45_Y33_N8
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_minor_ver_reg~3 (
	.dataa(gnd),
	.datab(\altera_internal_jtag~TDIUTAP ),
	.datac(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [3]),
	.datad(gnd),
	.cin(gnd),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_minor_ver_reg~3_combout ),
	.cout());
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_minor_ver_reg~3 .lut_mask = 16'h0C0C;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_minor_ver_reg~3 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X42_Y33_N12
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|WORD_SR~13 (
	.dataa(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter [0]),
	.datab(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter [1]),
	.datac(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [4]),
	.datad(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter [2]),
	.cin(gnd),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|WORD_SR~13_combout ),
	.cout());
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|WORD_SR~13 .lut_mask = 16'h0504;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|WORD_SR~13 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X43_Y33_N6
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|WORD_SR~14 (
	.dataa(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|WORD_SR~13_combout ),
	.datab(\altera_internal_jtag~TDIUTAP ),
	.datac(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [4]),
	.datad(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|clear_signal~combout ),
	.cin(gnd),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|WORD_SR~14_combout ),
	.cout());
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|WORD_SR~14 .lut_mask = 16'h00EA;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|WORD_SR~14 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X43_Y33_N8
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|WORD_SR[1]~15 (
	.dataa(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [3]),
	.datab(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|clear_signal~combout ),
	.datac(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [4]),
	.datad(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|virtual_dr_scan_reg~q ),
	.cin(gnd),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|WORD_SR[1]~15_combout ),
	.cout());
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|WORD_SR[1]~15 .lut_mask = 16'hFECC;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|WORD_SR[1]~15 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X42_Y33_N30
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter[1]~22 (
	.dataa(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter [4]),
	.datab(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|virtual_ir_scan_reg~q ),
	.datac(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter[1]~17_combout ),
	.datad(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [8]),
	.cin(gnd),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter[1]~22_combout ),
	.cout());
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter[1]~22 .lut_mask = 16'hCE0A;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter[1]~22 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X43_Y33_N2
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter[1]~23 (
	.dataa(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [3]),
	.datab(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|clear_signal~combout ),
	.datac(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [4]),
	.datad(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|virtual_dr_scan_reg~q ),
	.cin(gnd),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter[1]~23_combout ),
	.cout());
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter[1]~23 .lut_mask = 16'hCECC;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter[1]~23 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X42_Y33_N20
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|WORD_SR~16 (
	.dataa(gnd),
	.datab(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|virtual_ir_scan_reg~q ),
	.datac(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|WORD_SR~9_combout ),
	.datad(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [8]),
	.cin(gnd),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|WORD_SR~16_combout ),
	.cout());
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|WORD_SR~16 .lut_mask = 16'h30F0;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|WORD_SR~16 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X39_Y33_N10
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg~20 (
	.dataa(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg [3]),
	.datab(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg [4]),
	.datac(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg [2]),
	.datad(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg [0]),
	.cin(gnd),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg~20_combout ),
	.cout());
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg~20 .lut_mask = 16'h2106;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg~20 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X39_Y33_N20
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg~21 (
	.dataa(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg~20_combout ),
	.datab(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg [4]),
	.datac(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg [2]),
	.datad(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg [1]),
	.cin(gnd),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg~21_combout ),
	.cout());
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg~21 .lut_mask = 16'h2A2B;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg~21 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X39_Y33_N22
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg~22 (
	.dataa(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg [3]),
	.datab(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg [0]),
	.datac(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg [2]),
	.datad(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg [1]),
	.cin(gnd),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg~22_combout ),
	.cout());
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg~22 .lut_mask = 16'h5ED5;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg~22 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X39_Y33_N24
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg~23 (
	.dataa(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg~22_combout ),
	.datab(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg [4]),
	.datac(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg [2]),
	.datad(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg [1]),
	.cin(gnd),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg~23_combout ),
	.cout());
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg~23 .lut_mask = 16'h2628;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg~23 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: IOIBUF_X58_Y0_N8
cycloneive_io_ibuf \syif.tbCTRL~input (
	.i(\syif.tbCTRL ),
	.ibar(gnd),
	.o(\syif.tbCTRL~input_o ));
// synopsys translate_off
defparam \syif.tbCTRL~input .bus_hold = "false";
defparam \syif.tbCTRL~input .simulate_z_as = "z";
// synopsys translate_on

// Location: IOIBUF_X58_Y0_N1
cycloneive_io_ibuf \syif.addr[1]~input (
	.i(\syif.addr [1]),
	.ibar(gnd),
	.o(\syif.addr[1]~input_o ));
// synopsys translate_off
defparam \syif.addr[1]~input .bus_hold = "false";
defparam \syif.addr[1]~input .simulate_z_as = "z";
// synopsys translate_on

// Location: IOIBUF_X40_Y73_N1
cycloneive_io_ibuf \syif.addr[0]~input (
	.i(\syif.addr [0]),
	.ibar(gnd),
	.o(\syif.addr[0]~input_o ));
// synopsys translate_off
defparam \syif.addr[0]~input .bus_hold = "false";
defparam \syif.addr[0]~input .simulate_z_as = "z";
// synopsys translate_on

// Location: IOIBUF_X42_Y0_N15
cycloneive_io_ibuf \syif.addr[3]~input (
	.i(\syif.addr [3]),
	.ibar(gnd),
	.o(\syif.addr[3]~input_o ));
// synopsys translate_off
defparam \syif.addr[3]~input .bus_hold = "false";
defparam \syif.addr[3]~input .simulate_z_as = "z";
// synopsys translate_on

// Location: IOIBUF_X49_Y73_N15
cycloneive_io_ibuf \syif.addr[2]~input (
	.i(\syif.addr [2]),
	.ibar(gnd),
	.o(\syif.addr[2]~input_o ));
// synopsys translate_off
defparam \syif.addr[2]~input .bus_hold = "false";
defparam \syif.addr[2]~input .simulate_z_as = "z";
// synopsys translate_on

// Location: IOIBUF_X49_Y0_N8
cycloneive_io_ibuf \syif.addr[5]~input (
	.i(\syif.addr [5]),
	.ibar(gnd),
	.o(\syif.addr[5]~input_o ));
// synopsys translate_off
defparam \syif.addr[5]~input .bus_hold = "false";
defparam \syif.addr[5]~input .simulate_z_as = "z";
// synopsys translate_on

// Location: IOIBUF_X40_Y0_N22
cycloneive_io_ibuf \syif.addr[4]~input (
	.i(\syif.addr [4]),
	.ibar(gnd),
	.o(\syif.addr[4]~input_o ));
// synopsys translate_off
defparam \syif.addr[4]~input .bus_hold = "false";
defparam \syif.addr[4]~input .simulate_z_as = "z";
// synopsys translate_on

// Location: IOIBUF_X115_Y35_N15
cycloneive_io_ibuf \syif.addr[7]~input (
	.i(\syif.addr [7]),
	.ibar(gnd),
	.o(\syif.addr[7]~input_o ));
// synopsys translate_off
defparam \syif.addr[7]~input .bus_hold = "false";
defparam \syif.addr[7]~input .simulate_z_as = "z";
// synopsys translate_on

// Location: IOIBUF_X52_Y73_N22
cycloneive_io_ibuf \syif.addr[6]~input (
	.i(\syif.addr [6]),
	.ibar(gnd),
	.o(\syif.addr[6]~input_o ));
// synopsys translate_off
defparam \syif.addr[6]~input .bus_hold = "false";
defparam \syif.addr[6]~input .simulate_z_as = "z";
// synopsys translate_on

// Location: IOIBUF_X0_Y33_N22
cycloneive_io_ibuf \syif.addr[9]~input (
	.i(\syif.addr [9]),
	.ibar(gnd),
	.o(\syif.addr[9]~input_o ));
// synopsys translate_off
defparam \syif.addr[9]~input .bus_hold = "false";
defparam \syif.addr[9]~input .simulate_z_as = "z";
// synopsys translate_on

// Location: IOIBUF_X47_Y0_N1
cycloneive_io_ibuf \syif.addr[8]~input (
	.i(\syif.addr [8]),
	.ibar(gnd),
	.o(\syif.addr[8]~input_o ));
// synopsys translate_off
defparam \syif.addr[8]~input .bus_hold = "false";
defparam \syif.addr[8]~input .simulate_z_as = "z";
// synopsys translate_on

// Location: IOIBUF_X54_Y73_N1
cycloneive_io_ibuf \syif.addr[11]~input (
	.i(\syif.addr [11]),
	.ibar(gnd),
	.o(\syif.addr[11]~input_o ));
// synopsys translate_off
defparam \syif.addr[11]~input .bus_hold = "false";
defparam \syif.addr[11]~input .simulate_z_as = "z";
// synopsys translate_on

// Location: IOIBUF_X115_Y36_N1
cycloneive_io_ibuf \syif.addr[10]~input (
	.i(\syif.addr [10]),
	.ibar(gnd),
	.o(\syif.addr[10]~input_o ));
// synopsys translate_off
defparam \syif.addr[10]~input .bus_hold = "false";
defparam \syif.addr[10]~input .simulate_z_as = "z";
// synopsys translate_on

// Location: IOIBUF_X115_Y32_N1
cycloneive_io_ibuf \syif.addr[13]~input (
	.i(\syif.addr [13]),
	.ibar(gnd),
	.o(\syif.addr[13]~input_o ));
// synopsys translate_off
defparam \syif.addr[13]~input .bus_hold = "false";
defparam \syif.addr[13]~input .simulate_z_as = "z";
// synopsys translate_on

// Location: IOIBUF_X47_Y73_N15
cycloneive_io_ibuf \syif.addr[12]~input (
	.i(\syif.addr [12]),
	.ibar(gnd),
	.o(\syif.addr[12]~input_o ));
// synopsys translate_off
defparam \syif.addr[12]~input .bus_hold = "false";
defparam \syif.addr[12]~input .simulate_z_as = "z";
// synopsys translate_on

// Location: IOIBUF_X52_Y0_N15
cycloneive_io_ibuf \syif.addr[15]~input (
	.i(\syif.addr [15]),
	.ibar(gnd),
	.o(\syif.addr[15]~input_o ));
// synopsys translate_off
defparam \syif.addr[15]~input .bus_hold = "false";
defparam \syif.addr[15]~input .simulate_z_as = "z";
// synopsys translate_on

// Location: IOIBUF_X40_Y73_N8
cycloneive_io_ibuf \syif.addr[14]~input (
	.i(\syif.addr [14]),
	.ibar(gnd),
	.o(\syif.addr[14]~input_o ));
// synopsys translate_off
defparam \syif.addr[14]~input .bus_hold = "false";
defparam \syif.addr[14]~input .simulate_z_as = "z";
// synopsys translate_on

// Location: IOIBUF_X49_Y0_N22
cycloneive_io_ibuf \syif.addr[17]~input (
	.i(\syif.addr [17]),
	.ibar(gnd),
	.o(\syif.addr[17]~input_o ));
// synopsys translate_off
defparam \syif.addr[17]~input .bus_hold = "false";
defparam \syif.addr[17]~input .simulate_z_as = "z";
// synopsys translate_on

// Location: IOIBUF_X42_Y0_N22
cycloneive_io_ibuf \syif.addr[16]~input (
	.i(\syif.addr [16]),
	.ibar(gnd),
	.o(\syif.addr[16]~input_o ));
// synopsys translate_off
defparam \syif.addr[16]~input .bus_hold = "false";
defparam \syif.addr[16]~input .simulate_z_as = "z";
// synopsys translate_on

// Location: IOIBUF_X54_Y0_N8
cycloneive_io_ibuf \syif.addr[19]~input (
	.i(\syif.addr [19]),
	.ibar(gnd),
	.o(\syif.addr[19]~input_o ));
// synopsys translate_off
defparam \syif.addr[19]~input .bus_hold = "false";
defparam \syif.addr[19]~input .simulate_z_as = "z";
// synopsys translate_on

// Location: IOIBUF_X74_Y0_N8
cycloneive_io_ibuf \syif.addr[18]~input (
	.i(\syif.addr [18]),
	.ibar(gnd),
	.o(\syif.addr[18]~input_o ));
// synopsys translate_off
defparam \syif.addr[18]~input .bus_hold = "false";
defparam \syif.addr[18]~input .simulate_z_as = "z";
// synopsys translate_on

// Location: IOIBUF_X52_Y73_N15
cycloneive_io_ibuf \syif.addr[21]~input (
	.i(\syif.addr [21]),
	.ibar(gnd),
	.o(\syif.addr[21]~input_o ));
// synopsys translate_off
defparam \syif.addr[21]~input .bus_hold = "false";
defparam \syif.addr[21]~input .simulate_z_as = "z";
// synopsys translate_on

// Location: IOIBUF_X42_Y73_N8
cycloneive_io_ibuf \syif.addr[20]~input (
	.i(\syif.addr [20]),
	.ibar(gnd),
	.o(\syif.addr[20]~input_o ));
// synopsys translate_off
defparam \syif.addr[20]~input .bus_hold = "false";
defparam \syif.addr[20]~input .simulate_z_as = "z";
// synopsys translate_on

// Location: IOIBUF_X45_Y73_N8
cycloneive_io_ibuf \syif.addr[23]~input (
	.i(\syif.addr [23]),
	.ibar(gnd),
	.o(\syif.addr[23]~input_o ));
// synopsys translate_off
defparam \syif.addr[23]~input .bus_hold = "false";
defparam \syif.addr[23]~input .simulate_z_as = "z";
// synopsys translate_on

// Location: IOIBUF_X52_Y73_N1
cycloneive_io_ibuf \syif.addr[22]~input (
	.i(\syif.addr [22]),
	.ibar(gnd),
	.o(\syif.addr[22]~input_o ));
// synopsys translate_off
defparam \syif.addr[22]~input .bus_hold = "false";
defparam \syif.addr[22]~input .simulate_z_as = "z";
// synopsys translate_on

// Location: IOIBUF_X45_Y0_N15
cycloneive_io_ibuf \syif.addr[25]~input (
	.i(\syif.addr [25]),
	.ibar(gnd),
	.o(\syif.addr[25]~input_o ));
// synopsys translate_off
defparam \syif.addr[25]~input .bus_hold = "false";
defparam \syif.addr[25]~input .simulate_z_as = "z";
// synopsys translate_on

// Location: IOIBUF_X47_Y73_N1
cycloneive_io_ibuf \syif.addr[24]~input (
	.i(\syif.addr [24]),
	.ibar(gnd),
	.o(\syif.addr[24]~input_o ));
// synopsys translate_off
defparam \syif.addr[24]~input .bus_hold = "false";
defparam \syif.addr[24]~input .simulate_z_as = "z";
// synopsys translate_on

// Location: IOIBUF_X115_Y34_N15
cycloneive_io_ibuf \syif.addr[27]~input (
	.i(\syif.addr [27]),
	.ibar(gnd),
	.o(\syif.addr[27]~input_o ));
// synopsys translate_off
defparam \syif.addr[27]~input .bus_hold = "false";
defparam \syif.addr[27]~input .simulate_z_as = "z";
// synopsys translate_on

// Location: IOIBUF_X49_Y0_N15
cycloneive_io_ibuf \syif.addr[26]~input (
	.i(\syif.addr [26]),
	.ibar(gnd),
	.o(\syif.addr[26]~input_o ));
// synopsys translate_off
defparam \syif.addr[26]~input .bus_hold = "false";
defparam \syif.addr[26]~input .simulate_z_as = "z";
// synopsys translate_on

// Location: IOIBUF_X0_Y34_N15
cycloneive_io_ibuf \syif.addr[29]~input (
	.i(\syif.addr [29]),
	.ibar(gnd),
	.o(\syif.addr[29]~input_o ));
// synopsys translate_off
defparam \syif.addr[29]~input .bus_hold = "false";
defparam \syif.addr[29]~input .simulate_z_as = "z";
// synopsys translate_on

// Location: IOIBUF_X45_Y73_N1
cycloneive_io_ibuf \syif.addr[28]~input (
	.i(\syif.addr [28]),
	.ibar(gnd),
	.o(\syif.addr[28]~input_o ));
// synopsys translate_off
defparam \syif.addr[28]~input .bus_hold = "false";
defparam \syif.addr[28]~input .simulate_z_as = "z";
// synopsys translate_on

// Location: IOIBUF_X52_Y73_N8
cycloneive_io_ibuf \syif.addr[31]~input (
	.i(\syif.addr [31]),
	.ibar(gnd),
	.o(\syif.addr[31]~input_o ));
// synopsys translate_off
defparam \syif.addr[31]~input .bus_hold = "false";
defparam \syif.addr[31]~input .simulate_z_as = "z";
// synopsys translate_on

// Location: IOIBUF_X49_Y73_N22
cycloneive_io_ibuf \syif.addr[30]~input (
	.i(\syif.addr [30]),
	.ibar(gnd),
	.o(\syif.addr[30]~input_o ));
// synopsys translate_off
defparam \syif.addr[30]~input .bus_hold = "false";
defparam \syif.addr[30]~input .simulate_z_as = "z";
// synopsys translate_on

// Location: IOIBUF_X0_Y34_N22
cycloneive_io_ibuf \syif.WEN~input (
	.i(\syif.WEN ),
	.ibar(gnd),
	.o(\syif.WEN~input_o ));
// synopsys translate_off
defparam \syif.WEN~input .bus_hold = "false";
defparam \syif.WEN~input .simulate_z_as = "z";
// synopsys translate_on

// Location: IOIBUF_X115_Y34_N22
cycloneive_io_ibuf \syif.REN~input (
	.i(\syif.REN ),
	.ibar(gnd),
	.o(\syif.REN~input_o ));
// synopsys translate_off
defparam \syif.REN~input .bus_hold = "false";
defparam \syif.REN~input .simulate_z_as = "z";
// synopsys translate_on

// Location: IOIBUF_X0_Y36_N15
cycloneive_io_ibuf \nRST~input (
	.i(nRST),
	.ibar(gnd),
	.o(\nRST~input_o ));
// synopsys translate_off
defparam \nRST~input .bus_hold = "false";
defparam \nRST~input .simulate_z_as = "z";
// synopsys translate_on

// Location: IOIBUF_X0_Y36_N8
cycloneive_io_ibuf \CLK~input (
	.i(CLK),
	.ibar(gnd),
	.o(\CLK~input_o ));
// synopsys translate_off
defparam \CLK~input .bus_hold = "false";
defparam \CLK~input .simulate_z_as = "z";
// synopsys translate_on

// Location: IOIBUF_X67_Y73_N15
cycloneive_io_ibuf \syif.store[0]~input (
	.i(\syif.store [0]),
	.ibar(gnd),
	.o(\syif.store[0]~input_o ));
// synopsys translate_off
defparam \syif.store[0]~input .bus_hold = "false";
defparam \syif.store[0]~input .simulate_z_as = "z";
// synopsys translate_on

// Location: IOIBUF_X54_Y0_N22
cycloneive_io_ibuf \syif.store[1]~input (
	.i(\syif.store [1]),
	.ibar(gnd),
	.o(\syif.store[1]~input_o ));
// synopsys translate_off
defparam \syif.store[1]~input .bus_hold = "false";
defparam \syif.store[1]~input .simulate_z_as = "z";
// synopsys translate_on

// Location: IOIBUF_X60_Y73_N8
cycloneive_io_ibuf \syif.store[2]~input (
	.i(\syif.store [2]),
	.ibar(gnd),
	.o(\syif.store[2]~input_o ));
// synopsys translate_off
defparam \syif.store[2]~input .bus_hold = "false";
defparam \syif.store[2]~input .simulate_z_as = "z";
// synopsys translate_on

// Location: IOIBUF_X52_Y0_N1
cycloneive_io_ibuf \syif.store[3]~input (
	.i(\syif.store [3]),
	.ibar(gnd),
	.o(\syif.store[3]~input_o ));
// synopsys translate_off
defparam \syif.store[3]~input .bus_hold = "false";
defparam \syif.store[3]~input .simulate_z_as = "z";
// synopsys translate_on

// Location: IOIBUF_X0_Y34_N1
cycloneive_io_ibuf \syif.store[4]~input (
	.i(\syif.store [4]),
	.ibar(gnd),
	.o(\syif.store[4]~input_o ));
// synopsys translate_off
defparam \syif.store[4]~input .bus_hold = "false";
defparam \syif.store[4]~input .simulate_z_as = "z";
// synopsys translate_on

// Location: IOIBUF_X67_Y73_N1
cycloneive_io_ibuf \syif.store[5]~input (
	.i(\syif.store [5]),
	.ibar(gnd),
	.o(\syif.store[5]~input_o ));
// synopsys translate_off
defparam \syif.store[5]~input .bus_hold = "false";
defparam \syif.store[5]~input .simulate_z_as = "z";
// synopsys translate_on

// Location: IOIBUF_X54_Y0_N15
cycloneive_io_ibuf \syif.store[6]~input (
	.i(\syif.store [6]),
	.ibar(gnd),
	.o(\syif.store[6]~input_o ));
// synopsys translate_off
defparam \syif.store[6]~input .bus_hold = "false";
defparam \syif.store[6]~input .simulate_z_as = "z";
// synopsys translate_on

// Location: IOIBUF_X58_Y73_N22
cycloneive_io_ibuf \syif.store[7]~input (
	.i(\syif.store [7]),
	.ibar(gnd),
	.o(\syif.store[7]~input_o ));
// synopsys translate_off
defparam \syif.store[7]~input .bus_hold = "false";
defparam \syif.store[7]~input .simulate_z_as = "z";
// synopsys translate_on

// Location: IOIBUF_X0_Y34_N8
cycloneive_io_ibuf \syif.store[8]~input (
	.i(\syif.store [8]),
	.ibar(gnd),
	.o(\syif.store[8]~input_o ));
// synopsys translate_off
defparam \syif.store[8]~input .bus_hold = "false";
defparam \syif.store[8]~input .simulate_z_as = "z";
// synopsys translate_on

// Location: IOIBUF_X69_Y73_N22
cycloneive_io_ibuf \syif.store[9]~input (
	.i(\syif.store [9]),
	.ibar(gnd),
	.o(\syif.store[9]~input_o ));
// synopsys translate_off
defparam \syif.store[9]~input .bus_hold = "false";
defparam \syif.store[9]~input .simulate_z_as = "z";
// synopsys translate_on

// Location: IOIBUF_X52_Y0_N22
cycloneive_io_ibuf \syif.store[10]~input (
	.i(\syif.store [10]),
	.ibar(gnd),
	.o(\syif.store[10]~input_o ));
// synopsys translate_off
defparam \syif.store[10]~input .bus_hold = "false";
defparam \syif.store[10]~input .simulate_z_as = "z";
// synopsys translate_on

// Location: IOIBUF_X72_Y0_N8
cycloneive_io_ibuf \syif.store[11]~input (
	.i(\syif.store [11]),
	.ibar(gnd),
	.o(\syif.store[11]~input_o ));
// synopsys translate_off
defparam \syif.store[11]~input .bus_hold = "false";
defparam \syif.store[11]~input .simulate_z_as = "z";
// synopsys translate_on

// Location: IOIBUF_X58_Y73_N1
cycloneive_io_ibuf \syif.store[12]~input (
	.i(\syif.store [12]),
	.ibar(gnd),
	.o(\syif.store[12]~input_o ));
// synopsys translate_off
defparam \syif.store[12]~input .bus_hold = "false";
defparam \syif.store[12]~input .simulate_z_as = "z";
// synopsys translate_on

// Location: IOIBUF_X115_Y40_N8
cycloneive_io_ibuf \syif.store[13]~input (
	.i(\syif.store [13]),
	.ibar(gnd),
	.o(\syif.store[13]~input_o ));
// synopsys translate_off
defparam \syif.store[13]~input .bus_hold = "false";
defparam \syif.store[13]~input .simulate_z_as = "z";
// synopsys translate_on

// Location: IOIBUF_X54_Y73_N8
cycloneive_io_ibuf \syif.store[14]~input (
	.i(\syif.store [14]),
	.ibar(gnd),
	.o(\syif.store[14]~input_o ));
// synopsys translate_off
defparam \syif.store[14]~input .bus_hold = "false";
defparam \syif.store[14]~input .simulate_z_as = "z";
// synopsys translate_on

// Location: IOIBUF_X0_Y35_N15
cycloneive_io_ibuf \syif.store[15]~input (
	.i(\syif.store [15]),
	.ibar(gnd),
	.o(\syif.store[15]~input_o ));
// synopsys translate_off
defparam \syif.store[15]~input .bus_hold = "false";
defparam \syif.store[15]~input .simulate_z_as = "z";
// synopsys translate_on

// Location: IOIBUF_X0_Y30_N8
cycloneive_io_ibuf \syif.store[16]~input (
	.i(\syif.store [16]),
	.ibar(gnd),
	.o(\syif.store[16]~input_o ));
// synopsys translate_off
defparam \syif.store[16]~input .bus_hold = "false";
defparam \syif.store[16]~input .simulate_z_as = "z";
// synopsys translate_on

// Location: IOIBUF_X67_Y73_N8
cycloneive_io_ibuf \syif.store[17]~input (
	.i(\syif.store [17]),
	.ibar(gnd),
	.o(\syif.store[17]~input_o ));
// synopsys translate_off
defparam \syif.store[17]~input .bus_hold = "false";
defparam \syif.store[17]~input .simulate_z_as = "z";
// synopsys translate_on

// Location: IOIBUF_X56_Y0_N8
cycloneive_io_ibuf \syif.store[18]~input (
	.i(\syif.store [18]),
	.ibar(gnd),
	.o(\syif.store[18]~input_o ));
// synopsys translate_off
defparam \syif.store[18]~input .bus_hold = "false";
defparam \syif.store[18]~input .simulate_z_as = "z";
// synopsys translate_on

// Location: IOIBUF_X67_Y0_N8
cycloneive_io_ibuf \syif.store[19]~input (
	.i(\syif.store [19]),
	.ibar(gnd),
	.o(\syif.store[19]~input_o ));
// synopsys translate_off
defparam \syif.store[19]~input .bus_hold = "false";
defparam \syif.store[19]~input .simulate_z_as = "z";
// synopsys translate_on

// Location: IOIBUF_X38_Y73_N8
cycloneive_io_ibuf \syif.store[20]~input (
	.i(\syif.store [20]),
	.ibar(gnd),
	.o(\syif.store[20]~input_o ));
// synopsys translate_off
defparam \syif.store[20]~input .bus_hold = "false";
defparam \syif.store[20]~input .simulate_z_as = "z";
// synopsys translate_on

// Location: IOIBUF_X115_Y32_N8
cycloneive_io_ibuf \syif.store[21]~input (
	.i(\syif.store [21]),
	.ibar(gnd),
	.o(\syif.store[21]~input_o ));
// synopsys translate_off
defparam \syif.store[21]~input .bus_hold = "false";
defparam \syif.store[21]~input .simulate_z_as = "z";
// synopsys translate_on

// Location: IOIBUF_X60_Y73_N1
cycloneive_io_ibuf \syif.store[22]~input (
	.i(\syif.store [22]),
	.ibar(gnd),
	.o(\syif.store[22]~input_o ));
// synopsys translate_off
defparam \syif.store[22]~input .bus_hold = "false";
defparam \syif.store[22]~input .simulate_z_as = "z";
// synopsys translate_on

// Location: IOIBUF_X52_Y0_N8
cycloneive_io_ibuf \syif.store[23]~input (
	.i(\syif.store [23]),
	.ibar(gnd),
	.o(\syif.store[23]~input_o ));
// synopsys translate_off
defparam \syif.store[23]~input .bus_hold = "false";
defparam \syif.store[23]~input .simulate_z_as = "z";
// synopsys translate_on

// Location: IOIBUF_X0_Y29_N15
cycloneive_io_ibuf \syif.store[24]~input (
	.i(\syif.store [24]),
	.ibar(gnd),
	.o(\syif.store[24]~input_o ));
// synopsys translate_off
defparam \syif.store[24]~input .bus_hold = "false";
defparam \syif.store[24]~input .simulate_z_as = "z";
// synopsys translate_on

// Location: IOIBUF_X54_Y0_N1
cycloneive_io_ibuf \syif.store[25]~input (
	.i(\syif.store [25]),
	.ibar(gnd),
	.o(\syif.store[25]~input_o ));
// synopsys translate_off
defparam \syif.store[25]~input .bus_hold = "false";
defparam \syif.store[25]~input .simulate_z_as = "z";
// synopsys translate_on

// Location: IOIBUF_X45_Y0_N22
cycloneive_io_ibuf \syif.store[26]~input (
	.i(\syif.store [26]),
	.ibar(gnd),
	.o(\syif.store[26]~input_o ));
// synopsys translate_off
defparam \syif.store[26]~input .bus_hold = "false";
defparam \syif.store[26]~input .simulate_z_as = "z";
// synopsys translate_on

// Location: IOIBUF_X42_Y73_N1
cycloneive_io_ibuf \syif.store[27]~input (
	.i(\syif.store [27]),
	.ibar(gnd),
	.o(\syif.store[27]~input_o ));
// synopsys translate_off
defparam \syif.store[27]~input .bus_hold = "false";
defparam \syif.store[27]~input .simulate_z_as = "z";
// synopsys translate_on

// Location: IOIBUF_X65_Y73_N8
cycloneive_io_ibuf \syif.store[28]~input (
	.i(\syif.store [28]),
	.ibar(gnd),
	.o(\syif.store[28]~input_o ));
// synopsys translate_off
defparam \syif.store[28]~input .bus_hold = "false";
defparam \syif.store[28]~input .simulate_z_as = "z";
// synopsys translate_on

// Location: IOIBUF_X65_Y73_N15
cycloneive_io_ibuf \syif.store[29]~input (
	.i(\syif.store [29]),
	.ibar(gnd),
	.o(\syif.store[29]~input_o ));
// synopsys translate_off
defparam \syif.store[29]~input .bus_hold = "false";
defparam \syif.store[29]~input .simulate_z_as = "z";
// synopsys translate_on

// Location: IOIBUF_X69_Y0_N8
cycloneive_io_ibuf \syif.store[30]~input (
	.i(\syif.store [30]),
	.ibar(gnd),
	.o(\syif.store[30]~input_o ));
// synopsys translate_off
defparam \syif.store[30]~input .bus_hold = "false";
defparam \syif.store[30]~input .simulate_z_as = "z";
// synopsys translate_on

// Location: IOIBUF_X67_Y0_N1
cycloneive_io_ibuf \syif.store[31]~input (
	.i(\syif.store [31]),
	.ibar(gnd),
	.o(\syif.store[31]~input_o ));
// synopsys translate_off
defparam \syif.store[31]~input .bus_hold = "false";
defparam \syif.store[31]~input .simulate_z_as = "z";
// synopsys translate_on

// Location: CLKCTRL_G4
cycloneive_clkctrl \altera_internal_jtag~TCKUTAPclkctrl (
	.ena(vcc),
	.inclk({vcc,vcc,vcc,\altera_internal_jtag~TCKUTAP }),
	.clkselect(2'b00),
	.devclrn(devclrn),
	.devpor(devpor),
	.outclk(\altera_internal_jtag~TCKUTAPclkctrl_outclk ));
// synopsys translate_off
defparam \altera_internal_jtag~TCKUTAPclkctrl .clock_type = "global clock";
defparam \altera_internal_jtag~TCKUTAPclkctrl .ena_register_mode = "none";
// synopsys translate_on

// Location: CLKCTRL_G18
cycloneive_clkctrl \CPUCLK~clkctrl (
	.ena(vcc),
	.inclk({vcc,vcc,vcc,\CPUCLK~q }),
	.clkselect(2'b00),
	.devclrn(devclrn),
	.devpor(devpor),
	.outclk(\CPUCLK~clkctrl_outclk ));
// synopsys translate_off
defparam \CPUCLK~clkctrl .clock_type = "global clock";
defparam \CPUCLK~clkctrl .ena_register_mode = "none";
// synopsys translate_on

// Location: CLKCTRL_G1
cycloneive_clkctrl \nRST~inputclkctrl (
	.ena(vcc),
	.inclk({vcc,vcc,vcc,\nRST~input_o }),
	.clkselect(2'b00),
	.devclrn(devclrn),
	.devpor(devpor),
	.outclk(\nRST~inputclkctrl_outclk ));
// synopsys translate_off
defparam \nRST~inputclkctrl .clock_type = "global clock";
defparam \nRST~inputclkctrl .ena_register_mode = "none";
// synopsys translate_on

// Location: CLKCTRL_G2
cycloneive_clkctrl \CLK~inputclkctrl (
	.ena(vcc),
	.inclk({vcc,vcc,vcc,\CLK~input_o }),
	.clkselect(2'b00),
	.devclrn(devclrn),
	.devpor(devpor),
	.outclk(\CLK~inputclkctrl_outclk ));
// synopsys translate_off
defparam \CLK~inputclkctrl .clock_type = "global clock";
defparam \CLK~inputclkctrl .ena_register_mode = "none";
// synopsys translate_on

// Location: LCCOMB_X46_Y33_N22
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irf_reg[1][3]~feeder (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg [3]),
	.cin(gnd),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irf_reg[1][3]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irf_reg[1][3]~feeder .lut_mask = 16'hFF00;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irf_reg[1][3]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X46_Y33_N12
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irf_reg[1][0]~feeder (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg [0]),
	.cin(gnd),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irf_reg[1][0]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irf_reg[1][0]~feeder .lut_mask = 16'hFF00;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irf_reg[1][0]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X46_Y33_N0
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irf_reg[1][2]~feeder (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg [2]),
	.cin(gnd),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irf_reg[1][2]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irf_reg[1][2]~feeder .lut_mask = 16'hFF00;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irf_reg[1][2]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X46_Y33_N10
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irf_reg[1][1]~feeder (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg [1]),
	.cin(gnd),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irf_reg[1][1]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irf_reg[1][1]~feeder .lut_mask = 16'hFF00;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irf_reg[1][1]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X48_Y33_N20
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|identity_contrib_update_reg[1]~feeder (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|identity_contrib_shift_reg [1]),
	.cin(gnd),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|identity_contrib_update_reg[1]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|identity_contrib_update_reg[1]~feeder .lut_mask = 16'hFF00;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|identity_contrib_update_reg[1]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: IOOBUF_X49_Y0_N2
cycloneive_io_obuf \syif.halt~output (
	.i(\CPU|DP|EXMEM|plif_exmem.hlt_l~q ),
	.oe(vcc),
	.seriesterminationcontrol(16'b0000000000000000),
	.devoe(devoe),
	.o(\syif.halt ),
	.obar());
// synopsys translate_off
defparam \syif.halt~output .bus_hold = "false";
defparam \syif.halt~output .open_drain_output = "false";
// synopsys translate_on

// Location: IOOBUF_X0_Y32_N16
cycloneive_io_obuf \syif.load[0]~output (
	.i(\RAM|ramif.ramload[0]~0_combout ),
	.oe(vcc),
	.seriesterminationcontrol(16'b0000000000000000),
	.devoe(devoe),
	.o(\syif.load [0]),
	.obar());
// synopsys translate_off
defparam \syif.load[0]~output .bus_hold = "false";
defparam \syif.load[0]~output .open_drain_output = "false";
// synopsys translate_on

// Location: IOOBUF_X65_Y0_N9
cycloneive_io_obuf \syif.load[1]~output (
	.i(\RAM|ramif.ramload[1]~1_combout ),
	.oe(vcc),
	.seriesterminationcontrol(16'b0000000000000000),
	.devoe(devoe),
	.o(\syif.load [1]),
	.obar());
// synopsys translate_off
defparam \syif.load[1]~output .bus_hold = "false";
defparam \syif.load[1]~output .open_drain_output = "false";
// synopsys translate_on

// Location: IOOBUF_X60_Y0_N23
cycloneive_io_obuf \syif.load[2]~output (
	.i(\RAM|ramif.ramload[2]~2_combout ),
	.oe(vcc),
	.seriesterminationcontrol(16'b0000000000000000),
	.devoe(devoe),
	.o(\syif.load [2]),
	.obar());
// synopsys translate_off
defparam \syif.load[2]~output .bus_hold = "false";
defparam \syif.load[2]~output .open_drain_output = "false";
// synopsys translate_on

// Location: IOOBUF_X56_Y0_N16
cycloneive_io_obuf \syif.load[3]~output (
	.i(\RAM|ramif.ramload[3]~3_combout ),
	.oe(vcc),
	.seriesterminationcontrol(16'b0000000000000000),
	.devoe(devoe),
	.o(\syif.load [3]),
	.obar());
// synopsys translate_off
defparam \syif.load[3]~output .bus_hold = "false";
defparam \syif.load[3]~output .open_drain_output = "false";
// synopsys translate_on

// Location: IOOBUF_X67_Y0_N23
cycloneive_io_obuf \syif.load[4]~output (
	.i(\RAM|ramif.ramload[4]~4_combout ),
	.oe(vcc),
	.seriesterminationcontrol(16'b0000000000000000),
	.devoe(devoe),
	.o(\syif.load [4]),
	.obar());
// synopsys translate_off
defparam \syif.load[4]~output .bus_hold = "false";
defparam \syif.load[4]~output .open_drain_output = "false";
// synopsys translate_on

// Location: IOOBUF_X60_Y0_N2
cycloneive_io_obuf \syif.load[5]~output (
	.i(\RAM|ramif.ramload[5]~5_combout ),
	.oe(vcc),
	.seriesterminationcontrol(16'b0000000000000000),
	.devoe(devoe),
	.o(\syif.load [5]),
	.obar());
// synopsys translate_off
defparam \syif.load[5]~output .bus_hold = "false";
defparam \syif.load[5]~output .open_drain_output = "false";
// synopsys translate_on

// Location: IOOBUF_X56_Y0_N23
cycloneive_io_obuf \syif.load[6]~output (
	.i(\RAM|ramif.ramload[6]~6_combout ),
	.oe(vcc),
	.seriesterminationcontrol(16'b0000000000000000),
	.devoe(devoe),
	.o(\syif.load [6]),
	.obar());
// synopsys translate_off
defparam \syif.load[6]~output .bus_hold = "false";
defparam \syif.load[6]~output .open_drain_output = "false";
// synopsys translate_on

// Location: IOOBUF_X0_Y30_N2
cycloneive_io_obuf \syif.load[7]~output (
	.i(\RAM|ramif.ramload[7]~7_combout ),
	.oe(vcc),
	.seriesterminationcontrol(16'b0000000000000000),
	.devoe(devoe),
	.o(\syif.load [7]),
	.obar());
// synopsys translate_off
defparam \syif.load[7]~output .bus_hold = "false";
defparam \syif.load[7]~output .open_drain_output = "false";
// synopsys translate_on

// Location: IOOBUF_X0_Y32_N23
cycloneive_io_obuf \syif.load[8]~output (
	.i(\RAM|ramif.ramload[8]~8_combout ),
	.oe(vcc),
	.seriesterminationcontrol(16'b0000000000000000),
	.devoe(devoe),
	.o(\syif.load [8]),
	.obar());
// synopsys translate_off
defparam \syif.load[8]~output .bus_hold = "false";
defparam \syif.load[8]~output .open_drain_output = "false";
// synopsys translate_on

// Location: IOOBUF_X65_Y0_N2
cycloneive_io_obuf \syif.load[9]~output (
	.i(\RAM|ramif.ramload[9]~9_combout ),
	.oe(vcc),
	.seriesterminationcontrol(16'b0000000000000000),
	.devoe(devoe),
	.o(\syif.load [9]),
	.obar());
// synopsys translate_off
defparam \syif.load[9]~output .bus_hold = "false";
defparam \syif.load[9]~output .open_drain_output = "false";
// synopsys translate_on

// Location: IOOBUF_X60_Y73_N16
cycloneive_io_obuf \syif.load[10]~output (
	.i(\RAM|ramif.ramload[10]~10_combout ),
	.oe(vcc),
	.seriesterminationcontrol(16'b0000000000000000),
	.devoe(devoe),
	.o(\syif.load [10]),
	.obar());
// synopsys translate_off
defparam \syif.load[10]~output .bus_hold = "false";
defparam \syif.load[10]~output .open_drain_output = "false";
// synopsys translate_on

// Location: IOOBUF_X60_Y0_N16
cycloneive_io_obuf \syif.load[11]~output (
	.i(\RAM|ramif.ramload[11]~11_combout ),
	.oe(vcc),
	.seriesterminationcontrol(16'b0000000000000000),
	.devoe(devoe),
	.o(\syif.load [11]),
	.obar());
// synopsys translate_off
defparam \syif.load[11]~output .bus_hold = "false";
defparam \syif.load[11]~output .open_drain_output = "false";
// synopsys translate_on

// Location: IOOBUF_X56_Y0_N2
cycloneive_io_obuf \syif.load[12]~output (
	.i(\RAM|ramif.ramload[12]~12_combout ),
	.oe(vcc),
	.seriesterminationcontrol(16'b0000000000000000),
	.devoe(devoe),
	.o(\syif.load [12]),
	.obar());
// synopsys translate_off
defparam \syif.load[12]~output .bus_hold = "false";
defparam \syif.load[12]~output .open_drain_output = "false";
// synopsys translate_on

// Location: IOOBUF_X47_Y0_N9
cycloneive_io_obuf \syif.load[13]~output (
	.i(\RAM|ramif.ramload[13]~13_combout ),
	.oe(vcc),
	.seriesterminationcontrol(16'b0000000000000000),
	.devoe(devoe),
	.o(\syif.load [13]),
	.obar());
// synopsys translate_off
defparam \syif.load[13]~output .bus_hold = "false";
defparam \syif.load[13]~output .open_drain_output = "false";
// synopsys translate_on

// Location: IOOBUF_X62_Y0_N16
cycloneive_io_obuf \syif.load[14]~output (
	.i(\RAM|ramif.ramload[14]~14_combout ),
	.oe(vcc),
	.seriesterminationcontrol(16'b0000000000000000),
	.devoe(devoe),
	.o(\syif.load [14]),
	.obar());
// synopsys translate_off
defparam \syif.load[14]~output .bus_hold = "false";
defparam \syif.load[14]~output .open_drain_output = "false";
// synopsys translate_on

// Location: IOOBUF_X62_Y73_N23
cycloneive_io_obuf \syif.load[15]~output (
	.i(\RAM|ramif.ramload[15]~15_combout ),
	.oe(vcc),
	.seriesterminationcontrol(16'b0000000000000000),
	.devoe(devoe),
	.o(\syif.load [15]),
	.obar());
// synopsys translate_off
defparam \syif.load[15]~output .bus_hold = "false";
defparam \syif.load[15]~output .open_drain_output = "false";
// synopsys translate_on

// Location: IOOBUF_X0_Y35_N9
cycloneive_io_obuf \syif.load[16]~output (
	.i(\RAM|ramif.ramload[16]~16_combout ),
	.oe(vcc),
	.seriesterminationcontrol(16'b0000000000000000),
	.devoe(devoe),
	.o(\syif.load [16]),
	.obar());
// synopsys translate_off
defparam \syif.load[16]~output .bus_hold = "false";
defparam \syif.load[16]~output .open_drain_output = "false";
// synopsys translate_on

// Location: IOOBUF_X69_Y0_N2
cycloneive_io_obuf \syif.load[17]~output (
	.i(\RAM|ramif.ramload[17]~17_combout ),
	.oe(vcc),
	.seriesterminationcontrol(16'b0000000000000000),
	.devoe(devoe),
	.o(\syif.load [17]),
	.obar());
// synopsys translate_off
defparam \syif.load[17]~output .bus_hold = "false";
defparam \syif.load[17]~output .open_drain_output = "false";
// synopsys translate_on

// Location: IOOBUF_X62_Y73_N16
cycloneive_io_obuf \syif.load[18]~output (
	.i(\RAM|ramif.ramload[18]~18_combout ),
	.oe(vcc),
	.seriesterminationcontrol(16'b0000000000000000),
	.devoe(devoe),
	.o(\syif.load [18]),
	.obar());
// synopsys translate_off
defparam \syif.load[18]~output .bus_hold = "false";
defparam \syif.load[18]~output .open_drain_output = "false";
// synopsys translate_on

// Location: IOOBUF_X65_Y73_N23
cycloneive_io_obuf \syif.load[19]~output (
	.i(\RAM|ramif.ramload[19]~19_combout ),
	.oe(vcc),
	.seriesterminationcontrol(16'b0000000000000000),
	.devoe(devoe),
	.o(\syif.load [19]),
	.obar());
// synopsys translate_off
defparam \syif.load[19]~output .bus_hold = "false";
defparam \syif.load[19]~output .open_drain_output = "false";
// synopsys translate_on

// Location: IOOBUF_X65_Y0_N23
cycloneive_io_obuf \syif.load[20]~output (
	.i(\RAM|ramif.ramload[20]~20_combout ),
	.oe(vcc),
	.seriesterminationcontrol(16'b0000000000000000),
	.devoe(devoe),
	.o(\syif.load [20]),
	.obar());
// synopsys translate_off
defparam \syif.load[20]~output .bus_hold = "false";
defparam \syif.load[20]~output .open_drain_output = "false";
// synopsys translate_on

// Location: IOOBUF_X58_Y73_N9
cycloneive_io_obuf \syif.load[21]~output (
	.i(\RAM|ramif.ramload[21]~21_combout ),
	.oe(vcc),
	.seriesterminationcontrol(16'b0000000000000000),
	.devoe(devoe),
	.o(\syif.load [21]),
	.obar());
// synopsys translate_off
defparam \syif.load[21]~output .bus_hold = "false";
defparam \syif.load[21]~output .open_drain_output = "false";
// synopsys translate_on

// Location: IOOBUF_X72_Y0_N2
cycloneive_io_obuf \syif.load[22]~output (
	.i(\RAM|ramif.ramload[22]~22_combout ),
	.oe(vcc),
	.seriesterminationcontrol(16'b0000000000000000),
	.devoe(devoe),
	.o(\syif.load [22]),
	.obar());
// synopsys translate_off
defparam \syif.load[22]~output .bus_hold = "false";
defparam \syif.load[22]~output .open_drain_output = "false";
// synopsys translate_on

// Location: IOOBUF_X67_Y0_N16
cycloneive_io_obuf \syif.load[23]~output (
	.i(\RAM|ramif.ramload[23]~23_combout ),
	.oe(vcc),
	.seriesterminationcontrol(16'b0000000000000000),
	.devoe(devoe),
	.o(\syif.load [23]),
	.obar());
// synopsys translate_off
defparam \syif.load[23]~output .bus_hold = "false";
defparam \syif.load[23]~output .open_drain_output = "false";
// synopsys translate_on

// Location: IOOBUF_X60_Y73_N23
cycloneive_io_obuf \syif.load[24]~output (
	.i(\RAM|ramif.ramload[24]~24_combout ),
	.oe(vcc),
	.seriesterminationcontrol(16'b0000000000000000),
	.devoe(devoe),
	.o(\syif.load [24]),
	.obar());
// synopsys translate_off
defparam \syif.load[24]~output .bus_hold = "false";
defparam \syif.load[24]~output .open_drain_output = "false";
// synopsys translate_on

// Location: IOOBUF_X115_Y35_N23
cycloneive_io_obuf \syif.load[25]~output (
	.i(\RAM|ramif.ramload[25]~25_combout ),
	.oe(vcc),
	.seriesterminationcontrol(16'b0000000000000000),
	.devoe(devoe),
	.o(\syif.load [25]),
	.obar());
// synopsys translate_off
defparam \syif.load[25]~output .bus_hold = "false";
defparam \syif.load[25]~output .open_drain_output = "false";
// synopsys translate_on

// Location: IOOBUF_X58_Y73_N16
cycloneive_io_obuf \syif.load[26]~output (
	.i(\RAM|ramif.ramload[26]~26_combout ),
	.oe(vcc),
	.seriesterminationcontrol(16'b0000000000000000),
	.devoe(devoe),
	.o(\syif.load [26]),
	.obar());
// synopsys translate_off
defparam \syif.load[26]~output .bus_hold = "false";
defparam \syif.load[26]~output .open_drain_output = "false";
// synopsys translate_on

// Location: IOOBUF_X74_Y0_N23
cycloneive_io_obuf \syif.load[27]~output (
	.i(\RAM|ramif.ramload[27]~27_combout ),
	.oe(vcc),
	.seriesterminationcontrol(16'b0000000000000000),
	.devoe(devoe),
	.o(\syif.load [27]),
	.obar());
// synopsys translate_off
defparam \syif.load[27]~output .bus_hold = "false";
defparam \syif.load[27]~output .open_drain_output = "false";
// synopsys translate_on

// Location: IOOBUF_X65_Y0_N16
cycloneive_io_obuf \syif.load[28]~output (
	.i(\RAM|ramif.ramload[28]~28_combout ),
	.oe(vcc),
	.seriesterminationcontrol(16'b0000000000000000),
	.devoe(devoe),
	.o(\syif.load [28]),
	.obar());
// synopsys translate_off
defparam \syif.load[28]~output .bus_hold = "false";
defparam \syif.load[28]~output .open_drain_output = "false";
// synopsys translate_on

// Location: IOOBUF_X60_Y0_N9
cycloneive_io_obuf \syif.load[29]~output (
	.i(\RAM|ramif.ramload[29]~29_combout ),
	.oe(vcc),
	.seriesterminationcontrol(16'b0000000000000000),
	.devoe(devoe),
	.o(\syif.load [29]),
	.obar());
// synopsys translate_off
defparam \syif.load[29]~output .bus_hold = "false";
defparam \syif.load[29]~output .open_drain_output = "false";
// synopsys translate_on

// Location: IOOBUF_X62_Y0_N23
cycloneive_io_obuf \syif.load[30]~output (
	.i(\RAM|ramif.ramload[30]~30_combout ),
	.oe(vcc),
	.seriesterminationcontrol(16'b0000000000000000),
	.devoe(devoe),
	.o(\syif.load [30]),
	.obar());
// synopsys translate_off
defparam \syif.load[30]~output .bus_hold = "false";
defparam \syif.load[30]~output .open_drain_output = "false";
// synopsys translate_on

// Location: IOOBUF_X0_Y31_N16
cycloneive_io_obuf \syif.load[31]~output (
	.i(\RAM|ramif.ramload[31]~31_combout ),
	.oe(vcc),
	.seriesterminationcontrol(16'b0000000000000000),
	.devoe(devoe),
	.o(\syif.load [31]),
	.obar());
// synopsys translate_off
defparam \syif.load[31]~output .bus_hold = "false";
defparam \syif.load[31]~output .open_drain_output = "false";
// synopsys translate_on

// Location: IOOBUF_X0_Y37_N1
cycloneive_io_obuf \altera_reserved_tdo~output (
	.i(\altera_internal_jtag~TDO ),
	.oe(vcc),
	.seriesterminationcontrol(16'b0000000000000000),
	.devoe(devoe),
	.o(altera_reserved_tdo),
	.obar());
// synopsys translate_off
defparam \altera_reserved_tdo~output .bus_hold = "false";
defparam \altera_reserved_tdo~output .open_drain_output = "false";
// synopsys translate_on

// Location: IOIBUF_X0_Y38_N1
cycloneive_io_ibuf \altera_reserved_tms~input (
	.i(altera_reserved_tms),
	.ibar(gnd),
	.o(\altera_reserved_tms~input_o ));
// synopsys translate_off
defparam \altera_reserved_tms~input .bus_hold = "false";
defparam \altera_reserved_tms~input .simulate_z_as = "z";
// synopsys translate_on

// Location: IOIBUF_X0_Y39_N1
cycloneive_io_ibuf \altera_reserved_tck~input (
	.i(altera_reserved_tck),
	.ibar(gnd),
	.o(\altera_reserved_tck~input_o ));
// synopsys translate_off
defparam \altera_reserved_tck~input .bus_hold = "false";
defparam \altera_reserved_tck~input .simulate_z_as = "z";
// synopsys translate_on

// Location: IOIBUF_X0_Y40_N1
cycloneive_io_ibuf \altera_reserved_tdi~input (
	.i(altera_reserved_tdi),
	.ibar(gnd),
	.o(\altera_reserved_tdi~input_o ));
// synopsys translate_off
defparam \altera_reserved_tdi~input .bus_hold = "false";
defparam \altera_reserved_tdi~input .simulate_z_as = "z";
// synopsys translate_on

// Location: LCCOMB_X45_Y32_N0
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg[5]~0 (
	.dataa(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [4]),
	.datab(gnd),
	.datac(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg [5]),
	.datad(\altera_internal_jtag~TDIUTAP ),
	.cin(gnd),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg[5]~0_combout ),
	.cout());
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg[5]~0 .lut_mask = 16'hFA50;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg[5]~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X45_Y32_N22
cycloneive_lcell_comb \~QIC_CREATED_GND~I (
// Equation(s):
// \~QIC_CREATED_GND~I_combout  = GND

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\~QIC_CREATED_GND~I_combout ),
	.cout());
// synopsys translate_off
defparam \~QIC_CREATED_GND~I .lut_mask = 16'h0000;
defparam \~QIC_CREATED_GND~I .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X45_Y34_N8
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state~6 (
	.dataa(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [5]),
	.datab(gnd),
	.datac(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [6]),
	.datad(gnd),
	.cin(gnd),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state~6_combout ),
	.cout());
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state~6 .lut_mask = 16'hFAFA;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state~6 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X45_Y34_N9
dffeas \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state[6] (
	.clk(\altera_internal_jtag~TCKUTAPclkctrl_outclk ),
	.d(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state~6_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\altera_internal_jtag~TMSUTAP ),
	.sload(gnd),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [6]),
	.prn(vcc));
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state[6] .is_wysiwyg = "true";
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state[6] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X45_Y34_N10
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state~7 (
	.dataa(gnd),
	.datab(\altera_internal_jtag~TMSUTAP ),
	.datac(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [6]),
	.datad(gnd),
	.cin(gnd),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state~7_combout ),
	.cout());
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state~7 .lut_mask = 16'hC0C0;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state~7 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X45_Y34_N11
dffeas \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state[7] (
	.clk(\altera_internal_jtag~TCKUTAPclkctrl_outclk ),
	.d(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state~7_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [7]),
	.prn(vcc));
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state[7] .is_wysiwyg = "true";
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state[7] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X45_Y34_N22
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state~4 (
	.dataa(gnd),
	.datab(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [3]),
	.datac(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [4]),
	.datad(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [7]),
	.cin(gnd),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state~4_combout ),
	.cout());
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state~4 .lut_mask = 16'hFFFC;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state~4 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X45_Y34_N23
dffeas \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state[4] (
	.clk(\altera_internal_jtag~TCKUTAPclkctrl_outclk ),
	.d(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state~4_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\altera_internal_jtag~TMSUTAP ),
	.sload(gnd),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [4]),
	.prn(vcc));
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state[4] .is_wysiwyg = "true";
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state[4] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X45_Y34_N20
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state~5 (
	.dataa(gnd),
	.datab(\altera_internal_jtag~TMSUTAP ),
	.datac(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [4]),
	.datad(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [3]),
	.cin(gnd),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state~5_combout ),
	.cout());
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state~5 .lut_mask = 16'hCCC0;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state~5 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X45_Y34_N21
dffeas \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state[5] (
	.clk(\altera_internal_jtag~TCKUTAPclkctrl_outclk ),
	.d(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state~5_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [5]),
	.prn(vcc));
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state[5] .is_wysiwyg = "true";
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state[5] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X45_Y34_N24
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irf_proc~0 (
	.dataa(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [7]),
	.datab(\altera_internal_jtag~TMSUTAP ),
	.datac(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [5]),
	.datad(gnd),
	.cin(gnd),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irf_proc~0_combout ),
	.cout());
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irf_proc~0 .lut_mask = 16'hC8C8;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irf_proc~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X45_Y34_N25
dffeas \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state[8] (
	.clk(\altera_internal_jtag~TCKUTAPclkctrl_outclk ),
	.d(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irf_proc~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [8]),
	.prn(vcc));
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state[8] .is_wysiwyg = "true";
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state[8] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X45_Y33_N28
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|tms_cnt~1 (
	.dataa(gnd),
	.datab(\altera_internal_jtag~TMSUTAP ),
	.datac(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|tms_cnt [0]),
	.datad(gnd),
	.cin(gnd),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|tms_cnt~1_combout ),
	.cout());
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|tms_cnt~1 .lut_mask = 16'h0C0C;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|tms_cnt~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X45_Y33_N29
dffeas \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|tms_cnt[0] (
	.clk(\altera_internal_jtag~TCKUTAPclkctrl_outclk ),
	.d(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|tms_cnt~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|tms_cnt [0]),
	.prn(vcc));
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|tms_cnt[0] .is_wysiwyg = "true";
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|tms_cnt[0] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X45_Y33_N0
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|tms_cnt~0 (
	.dataa(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|tms_cnt [1]),
	.datab(gnd),
	.datac(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|tms_cnt [2]),
	.datad(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|tms_cnt [0]),
	.cin(gnd),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|tms_cnt~0_combout ),
	.cout());
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|tms_cnt~0 .lut_mask = 16'h5AF0;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|tms_cnt~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X45_Y33_N1
dffeas \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|tms_cnt[2] (
	.clk(\altera_internal_jtag~TCKUTAPclkctrl_outclk ),
	.d(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|tms_cnt~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!\altera_internal_jtag~TMSUTAP ),
	.sload(gnd),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|tms_cnt [2]),
	.prn(vcc));
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|tms_cnt[2] .is_wysiwyg = "true";
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|tms_cnt[2] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X45_Y33_N22
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state~0 (
	.dataa(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [9]),
	.datab(\altera_internal_jtag~TMSUTAP ),
	.datac(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [0]),
	.datad(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|tms_cnt [2]),
	.cin(gnd),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state~0_combout ),
	.cout());
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state~0 .lut_mask = 16'h3373;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X45_Y33_N23
dffeas \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state[0] (
	.clk(\altera_internal_jtag~TCKUTAPclkctrl_outclk ),
	.d(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [0]),
	.prn(vcc));
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state[0] .is_wysiwyg = "true";
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state[0] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X45_Y34_N4
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state~1 (
	.dataa(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [15]),
	.datab(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [8]),
	.datac(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [1]),
	.datad(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [0]),
	.cin(gnd),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state~1_combout ),
	.cout());
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state~1 .lut_mask = 16'hFEFF;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X45_Y34_N5
dffeas \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state[1] (
	.clk(\altera_internal_jtag~TCKUTAPclkctrl_outclk ),
	.d(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\altera_internal_jtag~TMSUTAP ),
	.sload(gnd),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [1]),
	.prn(vcc));
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state[1] .is_wysiwyg = "true";
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state[1] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X45_Y33_N20
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|node_ena_proc~1 (
	.dataa(gnd),
	.datab(gnd),
	.datac(\altera_internal_jtag~TMSUTAP ),
	.datad(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [2]),
	.cin(gnd),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|node_ena_proc~1_combout ),
	.cout());
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|node_ena_proc~1 .lut_mask = 16'hF000;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|node_ena_proc~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X45_Y33_N12
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state[9]~feeder (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|node_ena_proc~1_combout ),
	.cin(gnd),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state[9]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state[9]~feeder .lut_mask = 16'hFF00;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state[9]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X45_Y33_N13
dffeas \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state[9] (
	.clk(\altera_internal_jtag~TCKUTAPclkctrl_outclk ),
	.d(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state[9]~feeder_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [9]),
	.prn(vcc));
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state[9] .is_wysiwyg = "true";
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state[9] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X45_Y33_N10
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state~8 (
	.dataa(gnd),
	.datab(gnd),
	.datac(\altera_internal_jtag~TMSUTAP ),
	.datad(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [9]),
	.cin(gnd),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state~8_combout ),
	.cout());
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state~8 .lut_mask = 16'h0F00;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state~8 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X45_Y33_N11
dffeas \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state[10] (
	.clk(\altera_internal_jtag~TCKUTAPclkctrl_outclk ),
	.d(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state~8_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [10]),
	.prn(vcc));
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state[10] .is_wysiwyg = "true";
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state[10] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X45_Y34_N0
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state~11 (
	.dataa(gnd),
	.datab(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [12]),
	.datac(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [13]),
	.datad(gnd),
	.cin(gnd),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state~11_combout ),
	.cout());
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state~11 .lut_mask = 16'hFCFC;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state~11 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X45_Y34_N1
dffeas \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state[13] (
	.clk(\altera_internal_jtag~TCKUTAPclkctrl_outclk ),
	.d(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state~11_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\altera_internal_jtag~TMSUTAP ),
	.sload(gnd),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [13]),
	.prn(vcc));
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state[13] .is_wysiwyg = "true";
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state[13] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X45_Y34_N28
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state~12 (
	.dataa(gnd),
	.datab(\altera_internal_jtag~TMSUTAP ),
	.datac(gnd),
	.datad(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [13]),
	.cin(gnd),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state~12_combout ),
	.cout());
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state~12 .lut_mask = 16'hCC00;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state~12 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X45_Y34_N29
dffeas \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state[14] (
	.clk(\altera_internal_jtag~TCKUTAPclkctrl_outclk ),
	.d(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state~12_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [14]),
	.prn(vcc));
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state[14] .is_wysiwyg = "true";
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state[14] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X45_Y34_N2
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state~9 (
	.dataa(gnd),
	.datab(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [10]),
	.datac(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [11]),
	.datad(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [14]),
	.cin(gnd),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state~9_combout ),
	.cout());
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state~9 .lut_mask = 16'hFFFC;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state~9 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X45_Y34_N3
dffeas \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state[11] (
	.clk(\altera_internal_jtag~TCKUTAPclkctrl_outclk ),
	.d(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state~9_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\altera_internal_jtag~TMSUTAP ),
	.sload(gnd),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [11]),
	.prn(vcc));
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state[11] .is_wysiwyg = "true";
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state[11] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X45_Y34_N14
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state~10 (
	.dataa(gnd),
	.datab(\altera_internal_jtag~TMSUTAP ),
	.datac(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [10]),
	.datad(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [11]),
	.cin(gnd),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state~10_combout ),
	.cout());
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state~10 .lut_mask = 16'hCCC0;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state~10 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X45_Y34_N15
dffeas \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state[12] (
	.clk(\altera_internal_jtag~TCKUTAPclkctrl_outclk ),
	.d(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state~10_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [12]),
	.prn(vcc));
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state[12] .is_wysiwyg = "true";
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state[12] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X45_Y34_N30
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|virtual_ir_dr_scan_proc~0 (
	.dataa(gnd),
	.datab(\altera_internal_jtag~TMSUTAP ),
	.datac(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [12]),
	.datad(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [14]),
	.cin(gnd),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|virtual_ir_dr_scan_proc~0_combout ),
	.cout());
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|virtual_ir_dr_scan_proc~0 .lut_mask = 16'hCCC0;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|virtual_ir_dr_scan_proc~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X45_Y34_N31
dffeas \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state[15] (
	.clk(\altera_internal_jtag~TCKUTAPclkctrl_outclk ),
	.d(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|virtual_ir_dr_scan_proc~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [15]),
	.prn(vcc));
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state[15] .is_wysiwyg = "true";
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state[15] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X45_Y34_N16
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state~2 (
	.dataa(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [8]),
	.datab(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [1]),
	.datac(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [15]),
	.datad(\altera_internal_jtag~TMSUTAP ),
	.cin(gnd),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state~2_combout ),
	.cout());
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state~2 .lut_mask = 16'hFE00;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X45_Y34_N17
dffeas \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state[2] (
	.clk(\altera_internal_jtag~TCKUTAPclkctrl_outclk ),
	.d(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state~2_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [2]),
	.prn(vcc));
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state[2] .is_wysiwyg = "true";
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state[2] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X45_Y34_N26
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state~3 (
	.dataa(gnd),
	.datab(\altera_internal_jtag~TMSUTAP ),
	.datac(gnd),
	.datad(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [2]),
	.cin(gnd),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state~3_combout ),
	.cout());
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state~3 .lut_mask = 16'h3300;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state~3 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X45_Y34_N27
dffeas \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state[3] (
	.clk(\altera_internal_jtag~TCKUTAPclkctrl_outclk ),
	.d(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state~3_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [3]),
	.prn(vcc));
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state[3] .is_wysiwyg = "true";
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state[3] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X46_Y33_N24
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg~5 (
	.dataa(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg [3]),
	.datab(gnd),
	.datac(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [3]),
	.datad(\RAM|altsyncram_component|auto_generated|mgl_prim2|ir_loaded_address_reg [1]),
	.cin(gnd),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg~5_combout ),
	.cout());
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg~5 .lut_mask = 16'hFA0A;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg~5 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X43_Y34_N0
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg[9]~feeder (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(\altera_internal_jtag~TDIUTAP ),
	.cin(gnd),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg[9]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg[9]~feeder .lut_mask = 16'hFF00;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg[9]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X43_Y34_N1
dffeas \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg[9] (
	.clk(\altera_internal_jtag~TCKUTAPclkctrl_outclk ),
	.d(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg[9]~feeder_combout ),
	.asdata(vcc),
	.clrn(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [0]),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [11]),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg [9]),
	.prn(vcc));
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg[9] .is_wysiwyg = "true";
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg[9] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X43_Y34_N10
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg[8]~feeder (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg [9]),
	.cin(gnd),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg[8]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg[8]~feeder .lut_mask = 16'hFF00;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg[8]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X43_Y34_N11
dffeas \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg[8] (
	.clk(\altera_internal_jtag~TCKUTAPclkctrl_outclk ),
	.d(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg[8]~feeder_combout ),
	.asdata(vcc),
	.clrn(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [0]),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [11]),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg [8]),
	.prn(vcc));
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg[8] .is_wysiwyg = "true";
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg[8] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X43_Y34_N20
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg[7]~feeder (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg [8]),
	.cin(gnd),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg[7]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg[7]~feeder .lut_mask = 16'hFF00;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg[7]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X43_Y34_N21
dffeas \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg[7] (
	.clk(\altera_internal_jtag~TCKUTAPclkctrl_outclk ),
	.d(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg[7]~feeder_combout ),
	.asdata(vcc),
	.clrn(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [0]),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [11]),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg [7]),
	.prn(vcc));
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg[7] .is_wysiwyg = "true";
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg[7] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X43_Y34_N22
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg[6]~feeder (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg [7]),
	.cin(gnd),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg[6]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg[6]~feeder .lut_mask = 16'hFF00;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg[6]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X43_Y34_N23
dffeas \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg[6] (
	.clk(\altera_internal_jtag~TCKUTAPclkctrl_outclk ),
	.d(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg[6]~feeder_combout ),
	.asdata(vcc),
	.clrn(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [0]),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [11]),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg [6]),
	.prn(vcc));
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg[6] .is_wysiwyg = "true";
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg[6] .power_up = "low";
// synopsys translate_on

// Location: FF_X43_Y34_N29
dffeas \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg[5] (
	.clk(\altera_internal_jtag~TCKUTAPclkctrl_outclk ),
	.d(gnd),
	.asdata(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg [6]),
	.clrn(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [0]),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [11]),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg [5]),
	.prn(vcc));
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg[5] .is_wysiwyg = "true";
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg[5] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X43_Y34_N2
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg[4]~feeder (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg [5]),
	.cin(gnd),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg[4]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg[4]~feeder .lut_mask = 16'hFF00;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg[4]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X43_Y34_N3
dffeas \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg[4] (
	.clk(\altera_internal_jtag~TCKUTAPclkctrl_outclk ),
	.d(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg[4]~feeder_combout ),
	.asdata(vcc),
	.clrn(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [0]),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [11]),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg [4]),
	.prn(vcc));
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg[4] .is_wysiwyg = "true";
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg[4] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X43_Y34_N18
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg[3]~feeder (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg [4]),
	.cin(gnd),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg[3]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg[3]~feeder .lut_mask = 16'hFF00;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg[3]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X43_Y34_N19
dffeas \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg[3] (
	.clk(\altera_internal_jtag~TCKUTAPclkctrl_outclk ),
	.d(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg[3]~feeder_combout ),
	.asdata(vcc),
	.clrn(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [0]),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [11]),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg [3]),
	.prn(vcc));
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg[3] .is_wysiwyg = "true";
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg[3] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X43_Y34_N24
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg[2]~0 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg [3]),
	.cin(gnd),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg[2]~0_combout ),
	.cout());
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg[2]~0 .lut_mask = 16'h00FF;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg[2]~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X43_Y34_N25
dffeas \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg[2] (
	.clk(\altera_internal_jtag~TCKUTAPclkctrl_outclk ),
	.d(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg[2]~0_combout ),
	.asdata(vcc),
	.clrn(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [0]),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [11]),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg [2]),
	.prn(vcc));
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg[2] .is_wysiwyg = "true";
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg[2] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X43_Y34_N4
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg[1]~feeder (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg [2]),
	.cin(gnd),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg[1]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg[1]~feeder .lut_mask = 16'hFF00;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg[1]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X43_Y34_N5
dffeas \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg[1] (
	.clk(\altera_internal_jtag~TCKUTAPclkctrl_outclk ),
	.d(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg[1]~feeder_combout ),
	.asdata(vcc),
	.clrn(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [0]),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [11]),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg [1]),
	.prn(vcc));
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg[1] .is_wysiwyg = "true";
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg[1] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X43_Y34_N14
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg[0]~1 (
	.dataa(gnd),
	.datab(gnd),
	.datac(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg [1]),
	.datad(gnd),
	.cin(gnd),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg[0]~1_combout ),
	.cout());
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg[0]~1 .lut_mask = 16'h0F0F;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg[0]~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X43_Y34_N15
dffeas \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg[0] (
	.clk(\altera_internal_jtag~TCKUTAPclkctrl_outclk ),
	.d(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg[0]~1_combout ),
	.asdata(vcc),
	.clrn(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [0]),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [11]),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg [0]),
	.prn(vcc));
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg[0] .is_wysiwyg = "true";
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg[0] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X43_Y34_N6
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|Equal0~1 (
	.dataa(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg [5]),
	.datab(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg [2]),
	.datac(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg [3]),
	.datad(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg [4]),
	.cin(gnd),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|Equal0~1_combout ),
	.cout());
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|Equal0~1 .lut_mask = 16'h0010;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|Equal0~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X43_Y34_N16
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|Equal1~0 (
	.dataa(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|Equal0~0_combout ),
	.datab(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg [1]),
	.datac(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg [0]),
	.datad(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|Equal0~1_combout ),
	.cin(gnd),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|Equal1~0_combout ),
	.cout());
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|Equal1~0 .lut_mask = 16'h0200;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|Equal1~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X43_Y34_N17
dffeas \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|virtual_ir_scan_reg (
	.clk(\altera_internal_jtag~TCKUTAPclkctrl_outclk ),
	.d(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|Equal1~0_combout ),
	.asdata(vcc),
	.clrn(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [0]),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|virtual_ir_dr_scan_proc~0_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|virtual_ir_scan_reg~q ),
	.prn(vcc));
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|virtual_ir_scan_reg .is_wysiwyg = "true";
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|virtual_ir_scan_reg .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X43_Y33_N12
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg[3]~1 (
	.dataa(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg~7_combout ),
	.datab(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg[2]~3_combout ),
	.datac(gnd),
	.datad(\RAM|altsyncram_component|auto_generated|mgl_prim2|ir_loaded_address_reg [2]),
	.cin(gnd),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg[3]~1_combout ),
	.cout());
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg[3]~1 .lut_mask = 16'hEE22;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg[3]~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X46_Y33_N8
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg~9 (
	.dataa(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [3]),
	.datab(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg [5]),
	.datac(gnd),
	.datad(\RAM|altsyncram_component|auto_generated|mgl_prim2|ir_loaded_address_reg [3]),
	.cin(gnd),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg~9_combout ),
	.cout());
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg~9 .lut_mask = 16'hEE44;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg~9 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X46_Y33_N9
dffeas \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg[4] (
	.clk(\altera_internal_jtag~TCKUTAPclkctrl_outclk ),
	.d(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg~9_combout ),
	.asdata(vcc),
	.clrn(!\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|clr_reg~q ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg[0]~4_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg [4]),
	.prn(vcc));
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg[4] .is_wysiwyg = "true";
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg[4] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X43_Y33_N4
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg~8 (
	.dataa(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg [3]),
	.datab(gnd),
	.datac(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [4]),
	.datad(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg [4]),
	.cin(gnd),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg~8_combout ),
	.cout());
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg~8 .lut_mask = 16'hFA0A;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg~8 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X43_Y33_N13
dffeas \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg[3] (
	.clk(\altera_internal_jtag~TCKUTAPclkctrl_outclk ),
	.d(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg[3]~1_combout ),
	.asdata(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg~8_combout ),
	.clrn(!\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|clr_reg~q ),
	.aload(gnd),
	.sclr(gnd),
	.sload(!\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [3]),
	.ena(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|virtual_ir_scan_reg~q ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg [3]),
	.prn(vcc));
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg[3] .is_wysiwyg = "true";
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg[3] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X43_Y33_N20
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg[2]~3 (
	.dataa(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_mode_reg [0]),
	.datab(gnd),
	.datac(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg [5]),
	.datad(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg [3]),
	.cin(gnd),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg[2]~3_combout ),
	.cout());
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg[2]~3 .lut_mask = 16'hFA50;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg[2]~3 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X43_Y33_N18
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg[0]~4 (
	.dataa(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [3]),
	.datab(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [4]),
	.datac(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|virtual_ir_scan_reg~q ),
	.datad(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg[2]~3_combout ),
	.cin(gnd),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg[0]~4_combout ),
	.cout());
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg[0]~4 .lut_mask = 16'hE040;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg[0]~4 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X46_Y33_N25
dffeas \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg[2] (
	.clk(\altera_internal_jtag~TCKUTAPclkctrl_outclk ),
	.d(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg~5_combout ),
	.asdata(vcc),
	.clrn(!\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|clr_reg~q ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg[0]~4_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg [2]),
	.prn(vcc));
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg[2] .is_wysiwyg = "true";
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg[2] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X46_Y33_N20
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg~6 (
	.dataa(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [3]),
	.datab(gnd),
	.datac(\RAM|altsyncram_component|auto_generated|mgl_prim2|ir_loaded_address_reg [0]),
	.datad(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg [2]),
	.cin(gnd),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg~6_combout ),
	.cout());
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg~6 .lut_mask = 16'hF5A0;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg~6 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X46_Y33_N21
dffeas \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg[1] (
	.clk(\altera_internal_jtag~TCKUTAPclkctrl_outclk ),
	.d(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg~6_combout ),
	.asdata(vcc),
	.clrn(!\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|clr_reg~q ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg[0]~4_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg [1]),
	.prn(vcc));
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg[1] .is_wysiwyg = "true";
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg[1] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X46_Y33_N2
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg~2 (
	.dataa(gnd),
	.datab(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg [1]),
	.datac(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [3]),
	.datad(\RAM|altsyncram_component|auto_generated|mgl_prim2|is_in_use_reg~q ),
	.cin(gnd),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg~2_combout ),
	.cout());
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg~2 .lut_mask = 16'hFC0C;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X46_Y33_N3
dffeas \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg[0] (
	.clk(\altera_internal_jtag~TCKUTAPclkctrl_outclk ),
	.d(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg~2_combout ),
	.asdata(vcc),
	.clrn(!\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|clr_reg~q ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg[0]~4_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg [0]),
	.prn(vcc));
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg[0] .is_wysiwyg = "true";
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg[0] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X46_Y33_N6
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_mode_reg[1]~0 (
	.dataa(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg [2]),
	.datab(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg [1]),
	.datac(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_mode_reg [1]),
	.datad(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg [0]),
	.cin(gnd),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_mode_reg[1]~0_combout ),
	.cout());
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_mode_reg[1]~0 .lut_mask = 16'h21E0;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_mode_reg[1]~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X45_Y33_N24
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_mode_reg[1]~1 (
	.dataa(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|reset_ena_reg_proc~0_combout ),
	.datab(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg [5]),
	.datac(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_mode_reg [1]),
	.datad(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_mode_reg[1]~0_combout ),
	.cin(gnd),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_mode_reg[1]~1_combout ),
	.cout());
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_mode_reg[1]~1 .lut_mask = 16'hD2F0;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_mode_reg[1]~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X45_Y33_N25
dffeas \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_mode_reg[1] (
	.clk(\altera_internal_jtag~TCKUTAPclkctrl_outclk ),
	.d(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_mode_reg[1]~1_combout ),
	.asdata(vcc),
	.clrn(!\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|clr_reg~q ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_mode_reg [1]),
	.prn(vcc));
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_mode_reg[1] .is_wysiwyg = "true";
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_mode_reg[1] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X46_Y33_N4
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_mode_reg[2]~2 (
	.dataa(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg [2]),
	.datab(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg [1]),
	.datac(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_mode_reg [1]),
	.datad(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg [0]),
	.cin(gnd),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_mode_reg[2]~2_combout ),
	.cout());
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_mode_reg[2]~2 .lut_mask = 16'h0800;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_mode_reg[2]~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X45_Y34_N18
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_mode_reg[2]~3 (
	.dataa(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|reset_ena_reg~q ),
	.datab(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg [5]),
	.datac(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_mode_reg [2]),
	.datad(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_mode_reg[2]~2_combout ),
	.cin(gnd),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_mode_reg[2]~3_combout ),
	.cout());
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_mode_reg[2]~3 .lut_mask = 16'h7250;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_mode_reg[2]~3 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X45_Y34_N19
dffeas \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_mode_reg[2] (
	.clk(\altera_internal_jtag~TCKUTAPclkctrl_outclk ),
	.d(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_mode_reg[2]~3_combout ),
	.asdata(vcc),
	.clrn(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|virtual_ir_scan_reg~q ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_mode_reg [2]),
	.prn(vcc));
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_mode_reg[2] .is_wysiwyg = "true";
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_mode_reg[2] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X45_Y34_N6
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|clr_reg_proc~0 (
	.dataa(gnd),
	.datab(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_mode_reg [2]),
	.datac(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [1]),
	.datad(gnd),
	.cin(gnd),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|clr_reg_proc~0_combout ),
	.cout());
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|clr_reg_proc~0 .lut_mask = 16'hC0C0;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|clr_reg_proc~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X45_Y34_N7
dffeas \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|clr_reg (
	.clk(\altera_internal_jtag~TCKUTAPclkctrl_outclk ),
	.d(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|clr_reg_proc~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|clr_reg~q ),
	.prn(vcc));
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|clr_reg .is_wysiwyg = "true";
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|clr_reg .power_up = "low";
// synopsys translate_on

// Location: FF_X45_Y32_N1
dffeas \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg[5] (
	.clk(\altera_internal_jtag~TCKUTAPclkctrl_outclk ),
	.d(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg[5]~0_combout ),
	.asdata(\~QIC_CREATED_GND~I_combout ),
	.clrn(!\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|clr_reg~q ),
	.aload(gnd),
	.sclr(gnd),
	.sload(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [3]),
	.ena(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|virtual_ir_scan_reg~q ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg [5]),
	.prn(vcc));
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg[5] .is_wysiwyg = "true";
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg[5] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X45_Y32_N6
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|tdo_bypass_reg~0 (
	.dataa(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [4]),
	.datab(gnd),
	.datac(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|tdo_bypass_reg~q ),
	.datad(\altera_internal_jtag~TDIUTAP ),
	.cin(gnd),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|tdo_bypass_reg~0_combout ),
	.cout());
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|tdo_bypass_reg~0 .lut_mask = 16'hFA50;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|tdo_bypass_reg~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X45_Y32_N7
dffeas \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|tdo_bypass_reg (
	.clk(\altera_internal_jtag~TCKUTAPclkctrl_outclk ),
	.d(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|tdo_bypass_reg~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|tdo_bypass_reg~q ),
	.prn(vcc));
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|tdo_bypass_reg .is_wysiwyg = "true";
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|tdo_bypass_reg .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X47_Y33_N10
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|tdo~1 (
	.dataa(gnd),
	.datab(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg [1]),
	.datac(\RAM|altsyncram_component|auto_generated|mgl_prim2|tdo~1_combout ),
	.datad(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg [5]),
	.cin(gnd),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|tdo~1_combout ),
	.cout());
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|tdo~1 .lut_mask = 16'hF0CC;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|tdo~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X47_Y33_N28
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|tdo~2 (
	.dataa(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|tdo~0_combout ),
	.datab(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg [5]),
	.datac(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|tdo_bypass_reg~q ),
	.datad(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|tdo~1_combout ),
	.cin(gnd),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|tdo~2_combout ),
	.cout());
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|tdo~2 .lut_mask = 16'hFC22;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|tdo~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X40_Y33_N16
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg[0]~5 (
	.dataa(gnd),
	.datab(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg [0]),
	.datac(gnd),
	.datad(vcc),
	.cin(gnd),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg[0]~5_combout ),
	.cout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg[0]~6 ));
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg[0]~5 .lut_mask = 16'h33CC;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg[0]~5 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X43_Y33_N28
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|clear_signal (
	.dataa(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [8]),
	.datab(gnd),
	.datac(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|virtual_ir_scan_reg~q ),
	.datad(gnd),
	.cin(gnd),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|clear_signal~combout ),
	.cout());
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|clear_signal .lut_mask = 16'hA0A0;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|clear_signal .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X40_Y33_N20
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg[2]~9 (
	.dataa(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg [2]),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg[1]~8 ),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg[2]~9_combout ),
	.cout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg[2]~10 ));
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg[2]~9 .lut_mask = 16'h5AAF;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg[2]~9 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X43_Y34_N30
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|Equal0~2 (
	.dataa(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|Equal0~0_combout ),
	.datab(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg [1]),
	.datac(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg [0]),
	.datad(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|Equal0~1_combout ),
	.cin(gnd),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|Equal0~2_combout ),
	.cout());
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|Equal0~2 .lut_mask = 16'h0800;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|Equal0~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X43_Y34_N31
dffeas \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|virtual_dr_scan_reg (
	.clk(\altera_internal_jtag~TCKUTAPclkctrl_outclk ),
	.d(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|Equal0~2_combout ),
	.asdata(vcc),
	.clrn(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [0]),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|virtual_ir_dr_scan_proc~0_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|virtual_dr_scan_reg~q ),
	.prn(vcc));
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|virtual_dr_scan_reg .is_wysiwyg = "true";
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|virtual_dr_scan_reg .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X47_Y33_N4
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg[4]~12 (
	.dataa(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [8]),
	.datab(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|virtual_ir_scan_reg~q ),
	.datac(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [3]),
	.datad(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|virtual_dr_scan_reg~q ),
	.cin(gnd),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg[4]~12_combout ),
	.cout());
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg[4]~12 .lut_mask = 16'hF888;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg[4]~12 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X40_Y33_N21
dffeas \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg[2] (
	.clk(\altera_internal_jtag~TCKUTAPclkctrl_outclk ),
	.d(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg[2]~9_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg[4]~11_combout ),
	.ena(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg[4]~12_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg [2]),
	.prn(vcc));
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg[2] .is_wysiwyg = "true";
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg[2] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X40_Y33_N22
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg[3]~13 (
	.dataa(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg [3]),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg[2]~10 ),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg[3]~13_combout ),
	.cout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg[3]~14 ));
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg[3]~13 .lut_mask = 16'hA505;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg[3]~13 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: FF_X40_Y33_N23
dffeas \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg[3] (
	.clk(\altera_internal_jtag~TCKUTAPclkctrl_outclk ),
	.d(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg[3]~13_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg[4]~11_combout ),
	.ena(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg[4]~12_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg [3]),
	.prn(vcc));
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg[3] .is_wysiwyg = "true";
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg[3] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X41_Y33_N12
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg~12 (
	.dataa(gnd),
	.datab(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg [2]),
	.datac(gnd),
	.datad(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg [3]),
	.cin(gnd),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg~12_combout ),
	.cout());
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg~12 .lut_mask = 16'h0033;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg~12 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X41_Y33_N18
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg[4]~11 (
	.dataa(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg~15_combout ),
	.datab(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|clear_signal~combout ),
	.datac(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg [0]),
	.datad(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg~12_combout ),
	.cin(gnd),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg[4]~11_combout ),
	.cout());
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg[4]~11 .lut_mask = 16'hCECC;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg[4]~11 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X40_Y33_N17
dffeas \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg[0] (
	.clk(\altera_internal_jtag~TCKUTAPclkctrl_outclk ),
	.d(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg[0]~5_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg[4]~11_combout ),
	.ena(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg[4]~12_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg [0]),
	.prn(vcc));
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg[0] .is_wysiwyg = "true";
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg[0] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X40_Y33_N18
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg[1]~7 (
	.dataa(gnd),
	.datab(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg [1]),
	.datac(gnd),
	.datad(vcc),
	.cin(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg[0]~6 ),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg[1]~7_combout ),
	.cout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg[1]~8 ));
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg[1]~7 .lut_mask = 16'hC303;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg[1]~7 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: FF_X40_Y33_N19
dffeas \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg[1] (
	.clk(\altera_internal_jtag~TCKUTAPclkctrl_outclk ),
	.d(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg[1]~7_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg[4]~11_combout ),
	.ena(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg[4]~12_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg [1]),
	.prn(vcc));
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg[1] .is_wysiwyg = "true";
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg[1] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X40_Y33_N24
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg[4]~15 (
	.dataa(gnd),
	.datab(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg [4]),
	.datac(gnd),
	.datad(gnd),
	.cin(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg[3]~14 ),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg[4]~15_combout ),
	.cout());
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg[4]~15 .lut_mask = 16'h3C3C;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg[4]~15 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: FF_X40_Y33_N25
dffeas \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg[4] (
	.clk(\altera_internal_jtag~TCKUTAPclkctrl_outclk ),
	.d(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg[4]~15_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg[4]~11_combout ),
	.ena(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg[4]~12_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg [4]),
	.prn(vcc));
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg[4] .is_wysiwyg = "true";
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg[4] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X40_Y33_N6
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg[3]~14 (
	.dataa(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg[3]~13_combout ),
	.datab(gnd),
	.datac(gnd),
	.datad(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg [4]),
	.cin(gnd),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg[3]~14_combout ),
	.cout());
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg[3]~14 .lut_mask = 16'hAA00;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg[3]~14 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X48_Y33_N22
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|identity_contrib_shift_reg[3]~feeder (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(\altera_internal_jtag~TDIUTAP ),
	.cin(gnd),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|identity_contrib_shift_reg[3]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|identity_contrib_shift_reg[3]~feeder .lut_mask = 16'hFF00;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|identity_contrib_shift_reg[3]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X47_Y33_N20
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|identity_contrib_shift_reg[0]~0 (
	.dataa(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg [0]),
	.datab(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg [2]),
	.datac(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|virtual_dr_scan_reg~q ),
	.datad(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg [1]),
	.cin(gnd),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|identity_contrib_shift_reg[0]~0_combout ),
	.cout());
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|identity_contrib_shift_reg[0]~0 .lut_mask = 16'h4000;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|identity_contrib_shift_reg[0]~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X47_Y33_N0
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|identity_contrib_shift_reg[0]~1 (
	.dataa(gnd),
	.datab(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg [5]),
	.datac(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [4]),
	.datad(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|identity_contrib_shift_reg[0]~0_combout ),
	.cin(gnd),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|identity_contrib_shift_reg[0]~1_combout ),
	.cout());
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|identity_contrib_shift_reg[0]~1 .lut_mask = 16'h3000;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|identity_contrib_shift_reg[0]~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X48_Y33_N23
dffeas \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|identity_contrib_shift_reg[3] (
	.clk(\altera_internal_jtag~TCKUTAPclkctrl_outclk ),
	.d(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|identity_contrib_shift_reg[3]~feeder_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|identity_contrib_shift_reg[0]~1_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|identity_contrib_shift_reg [3]),
	.prn(vcc));
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|identity_contrib_shift_reg[3] .is_wysiwyg = "true";
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|identity_contrib_shift_reg[3] .power_up = "low";
// synopsys translate_on

// Location: FF_X48_Y33_N11
dffeas \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|identity_contrib_shift_reg[2] (
	.clk(\altera_internal_jtag~TCKUTAPclkctrl_outclk ),
	.d(gnd),
	.asdata(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|identity_contrib_shift_reg [3]),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|identity_contrib_shift_reg[0]~1_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|identity_contrib_shift_reg [2]),
	.prn(vcc));
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|identity_contrib_shift_reg[2] .is_wysiwyg = "true";
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|identity_contrib_shift_reg[2] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X48_Y33_N18
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|identity_contrib_shift_reg[1]~feeder (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|identity_contrib_shift_reg [2]),
	.cin(gnd),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|identity_contrib_shift_reg[1]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|identity_contrib_shift_reg[1]~feeder .lut_mask = 16'hFF00;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|identity_contrib_shift_reg[1]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X48_Y33_N19
dffeas \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|identity_contrib_shift_reg[1] (
	.clk(\altera_internal_jtag~TCKUTAPclkctrl_outclk ),
	.d(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|identity_contrib_shift_reg[1]~feeder_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|identity_contrib_shift_reg[0]~1_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|identity_contrib_shift_reg [1]),
	.prn(vcc));
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|identity_contrib_shift_reg[1] .is_wysiwyg = "true";
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|identity_contrib_shift_reg[1] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X48_Y33_N2
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|identity_contrib_shift_reg[0]~feeder (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|identity_contrib_shift_reg [1]),
	.cin(gnd),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|identity_contrib_shift_reg[0]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|identity_contrib_shift_reg[0]~feeder .lut_mask = 16'hFF00;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|identity_contrib_shift_reg[0]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X48_Y33_N3
dffeas \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|identity_contrib_shift_reg[0] (
	.clk(\altera_internal_jtag~TCKUTAPclkctrl_outclk ),
	.d(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|identity_contrib_shift_reg[0]~feeder_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|identity_contrib_shift_reg[0]~1_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|identity_contrib_shift_reg [0]),
	.prn(vcc));
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|identity_contrib_shift_reg[0] .is_wysiwyg = "true";
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|identity_contrib_shift_reg[0] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X48_Y33_N24
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|identity_contrib_update_reg[0]~feeder (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|identity_contrib_shift_reg [0]),
	.cin(gnd),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|identity_contrib_update_reg[0]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|identity_contrib_update_reg[0]~feeder .lut_mask = 16'hFF00;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|identity_contrib_update_reg[0]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X47_Y33_N6
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|identity_contrib_update_reg[0]~0 (
	.dataa(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [8]),
	.datab(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg [5]),
	.datac(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [4]),
	.datad(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|identity_contrib_shift_reg[0]~0_combout ),
	.cin(gnd),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|identity_contrib_update_reg[0]~0_combout ),
	.cout());
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|identity_contrib_update_reg[0]~0 .lut_mask = 16'h0200;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|identity_contrib_update_reg[0]~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X48_Y33_N25
dffeas \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|identity_contrib_update_reg[0] (
	.clk(\altera_internal_jtag~TCKUTAPclkctrl_outclk ),
	.d(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|identity_contrib_update_reg[0]~feeder_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|identity_contrib_update_reg[0]~0_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|identity_contrib_update_reg [0]),
	.prn(vcc));
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|identity_contrib_update_reg[0] .is_wysiwyg = "true";
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|identity_contrib_update_reg[0] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X47_Y33_N26
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg[0]~0 (
	.dataa(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg~23_combout ),
	.datab(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg[3]~14_combout ),
	.datac(gnd),
	.datad(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|identity_contrib_update_reg [0]),
	.cin(gnd),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg[0]~0_combout ),
	.cout());
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg[0]~0 .lut_mask = 16'hEE22;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg[0]~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X39_Y33_N2
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg~11 (
	.dataa(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg [3]),
	.datab(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg [4]),
	.datac(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg [2]),
	.datad(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg [0]),
	.cin(gnd),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg~11_combout ),
	.cout());
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg~11 .lut_mask = 16'h1024;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg~11 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X39_Y33_N4
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg~10 (
	.dataa(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg [3]),
	.datab(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg [4]),
	.datac(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg [2]),
	.datad(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg [0]),
	.cin(gnd),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg~10_combout ),
	.cout());
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg~10 .lut_mask = 16'h3714;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg~10 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X39_Y33_N12
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg~19 (
	.dataa(gnd),
	.datab(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg~11_combout ),
	.datac(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg~10_combout ),
	.datad(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg [1]),
	.cin(gnd),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg~19_combout ),
	.cout());
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg~19 .lut_mask = 16'hCCF0;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg~19 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X47_Y33_N30
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg[1]~1 (
	.dataa(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|identity_contrib_update_reg [1]),
	.datab(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg[3]~14_combout ),
	.datac(gnd),
	.datad(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg~19_combout ),
	.cin(gnd),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg[1]~1_combout ),
	.cout());
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg[1]~1 .lut_mask = 16'hBB88;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg[1]~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X48_Y33_N4
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|identity_contrib_update_reg[2]~feeder (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|identity_contrib_shift_reg [2]),
	.cin(gnd),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|identity_contrib_update_reg[2]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|identity_contrib_update_reg[2]~feeder .lut_mask = 16'hFF00;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|identity_contrib_update_reg[2]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X48_Y33_N5
dffeas \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|identity_contrib_update_reg[2] (
	.clk(\altera_internal_jtag~TCKUTAPclkctrl_outclk ),
	.d(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|identity_contrib_update_reg[2]~feeder_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|identity_contrib_update_reg[0]~0_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|identity_contrib_update_reg [2]),
	.prn(vcc));
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|identity_contrib_update_reg[2] .is_wysiwyg = "true";
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|identity_contrib_update_reg[2] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X47_Y33_N14
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg[2]~2 (
	.dataa(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg~18_combout ),
	.datab(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg[3]~14_combout ),
	.datac(gnd),
	.datad(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|identity_contrib_update_reg [2]),
	.cin(gnd),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg[2]~2_combout ),
	.cout());
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg[2]~2 .lut_mask = 16'hEE22;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg[2]~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X48_Y33_N17
dffeas \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|identity_contrib_update_reg[3] (
	.clk(\altera_internal_jtag~TCKUTAPclkctrl_outclk ),
	.d(gnd),
	.asdata(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|identity_contrib_shift_reg [3]),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|identity_contrib_update_reg[0]~0_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|identity_contrib_update_reg [3]),
	.prn(vcc));
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|identity_contrib_update_reg[3] .is_wysiwyg = "true";
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|identity_contrib_update_reg[3] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X47_Y33_N8
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg[3]~3 (
	.dataa(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg~21_combout ),
	.datab(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg[3]~14_combout ),
	.datac(gnd),
	.datad(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|identity_contrib_update_reg [3]),
	.cin(gnd),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg[3]~3_combout ),
	.cout());
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg[3]~3 .lut_mask = 16'hEE22;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg[3]~3 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X47_Y33_N16
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_proc~0 (
	.dataa(gnd),
	.datab(gnd),
	.datac(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [3]),
	.datad(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|virtual_dr_scan_reg~q ),
	.cin(gnd),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_proc~0_combout ),
	.cout());
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_proc~0 .lut_mask = 16'h0FFF;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_proc~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X47_Y33_N24
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg_ena (
	.dataa(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [4]),
	.datab(gnd),
	.datac(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [3]),
	.datad(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|virtual_dr_scan_reg~q ),
	.cin(gnd),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg_ena~combout ),
	.cout());
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg_ena .lut_mask = 16'hFA00;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg_ena .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X47_Y33_N9
dffeas \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg[3] (
	.clk(\altera_internal_jtag~TCKUTAPclkctrl_outclk ),
	.d(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg[3]~3_combout ),
	.asdata(\altera_internal_jtag~TDIUTAP ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_proc~0_combout ),
	.ena(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg_ena~combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg [3]),
	.prn(vcc));
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg[3] .is_wysiwyg = "true";
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg[3] .power_up = "low";
// synopsys translate_on

// Location: FF_X47_Y33_N15
dffeas \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg[2] (
	.clk(\altera_internal_jtag~TCKUTAPclkctrl_outclk ),
	.d(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg[2]~2_combout ),
	.asdata(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg [3]),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_proc~0_combout ),
	.ena(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg_ena~combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg [2]),
	.prn(vcc));
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg[2] .is_wysiwyg = "true";
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg[2] .power_up = "low";
// synopsys translate_on

// Location: FF_X47_Y33_N31
dffeas \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg[1] (
	.clk(\altera_internal_jtag~TCKUTAPclkctrl_outclk ),
	.d(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg[1]~1_combout ),
	.asdata(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg [2]),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_proc~0_combout ),
	.ena(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg_ena~combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg [1]),
	.prn(vcc));
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg[1] .is_wysiwyg = "true";
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg[1] .power_up = "low";
// synopsys translate_on

// Location: FF_X47_Y33_N27
dffeas \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg[0] (
	.clk(\altera_internal_jtag~TCKUTAPclkctrl_outclk ),
	.d(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg[0]~0_combout ),
	.asdata(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg [1]),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_proc~0_combout ),
	.ena(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg_ena~combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg [0]),
	.prn(vcc));
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg[0] .is_wysiwyg = "true";
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg[0] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X47_Y33_N12
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|tdo~3 (
	.dataa(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|tdo~0_combout ),
	.datab(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg [5]),
	.datac(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|tdo_bypass_reg~q ),
	.datad(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|tdo~1_combout ),
	.cin(gnd),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|tdo~3_combout ),
	.cout());
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|tdo~3 .lut_mask = 16'hFC10;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|tdo~3 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X47_Y33_N18
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|tdo~4 (
	.dataa(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg [0]),
	.datab(gnd),
	.datac(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|virtual_ir_scan_reg~q ),
	.datad(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|tdo~3_combout ),
	.cin(gnd),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|tdo~4_combout ),
	.cout());
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|tdo~4 .lut_mask = 16'hFAF0;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|tdo~4 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X47_Y33_N22
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|tdo~5 (
	.dataa(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg [0]),
	.datab(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|tdo~2_combout ),
	.datac(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg [0]),
	.datad(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|tdo~4_combout ),
	.cin(gnd),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|tdo~5_combout ),
	.cout());
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|tdo~5 .lut_mask = 16'h553B;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|tdo~5 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X45_Y33_N30
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg_ena~0 (
	.dataa(gnd),
	.datab(gnd),
	.datac(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [3]),
	.datad(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [4]),
	.cin(gnd),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg_ena~0_combout ),
	.cout());
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg_ena~0 .lut_mask = 16'hFFF0;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg_ena~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X47_Y33_N23
dffeas \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|tdo (
	.clk(!\altera_internal_jtag~TCKUTAPclkctrl_outclk ),
	.d(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|tdo~5_combout ),
	.asdata(vcc),
	.clrn(!\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [8]),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg_ena~0_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|tdo~q ),
	.prn(vcc));
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|tdo .is_wysiwyg = "true";
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|tdo .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X16_Y37_N0
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|tdo~_wirecell (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|tdo~q ),
	.cin(gnd),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|tdo~_wirecell_combout ),
	.cout());
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|tdo~_wirecell .lut_mask = 16'h00FF;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|tdo~_wirecell .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X81_Y16_N0
cycloneive_lcell_comb \auto_hub|~GND (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\auto_hub|~GND~combout ),
	.cout());
// synopsys translate_off
defparam \auto_hub|~GND .lut_mask = 16'h0000;
defparam \auto_hub|~GND .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X46_Y33_N16
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|clr_reg~_wirecell (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|clr_reg~q ),
	.cin(gnd),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|clr_reg~_wirecell_combout ),
	.cout());
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|clr_reg~_wirecell .lut_mask = 16'h00FF;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|clr_reg~_wirecell .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X45_Y33_N2
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state[0]~_wirecell (
	.dataa(gnd),
	.datab(gnd),
	.datac(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [0]),
	.datad(gnd),
	.cin(gnd),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state[0]~_wirecell_combout ),
	.cout());
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state[0]~_wirecell .lut_mask = 16'h0F0F;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state[0]~_wirecell .sum_lutc_input = "datac";
// synopsys translate_on

endmodule

module pipeline (
	PCreg_1,
	PCreg_0,
	plif_exmemhlt_l,
	plif_exmemporto_l_1,
	plif_exmemdmemWEN_l,
	plif_exmemdmemREN_l,
	plif_exmemporto_l_0,
	plif_exmemporto_l_3,
	PCreg_3,
	plif_exmemporto_l_2,
	PCreg_2,
	plif_exmemporto_l_5,
	PCreg_5,
	plif_exmemporto_l_4,
	PCreg_4,
	plif_exmemporto_l_7,
	PCreg_7,
	plif_exmemporto_l_6,
	PCreg_6,
	plif_exmemporto_l_9,
	PCreg_9,
	plif_exmemporto_l_8,
	PCreg_8,
	plif_exmemporto_l_11,
	PCreg_11,
	plif_exmemporto_l_10,
	PCreg_10,
	plif_exmemporto_l_13,
	PCreg_13,
	plif_exmemporto_l_12,
	PCreg_12,
	plif_exmemporto_l_15,
	PCreg_15,
	plif_exmemporto_l_14,
	PCreg_14,
	plif_exmemporto_l_17,
	PCreg_17,
	plif_exmemporto_l_16,
	PCreg_16,
	plif_exmemporto_l_19,
	PCreg_19,
	plif_exmemporto_l_18,
	PCreg_18,
	plif_exmemporto_l_21,
	PCreg_21,
	plif_exmemporto_l_20,
	PCreg_20,
	plif_exmemporto_l_23,
	PCreg_23,
	plif_exmemporto_l_22,
	PCreg_22,
	plif_exmemporto_l_25,
	PCreg_25,
	plif_exmemporto_l_24,
	PCreg_24,
	plif_exmemporto_l_27,
	PCreg_27,
	plif_exmemporto_l_26,
	PCreg_26,
	plif_exmemporto_l_29,
	PCreg_29,
	plif_exmemporto_l_28,
	PCreg_28,
	plif_exmemporto_l_31,
	PCreg_31,
	plif_exmemporto_l_30,
	PCreg_30,
	dpifimemREN,
	always1,
	ramiframload_0,
	ramiframload_1,
	ramiframload_2,
	ramiframload_3,
	ramiframload_4,
	ramiframload_5,
	ramiframload_6,
	ramiframload_7,
	ramiframload_8,
	ramiframload_9,
	ramiframload_10,
	ramiframload_11,
	ramiframload_12,
	ramiframload_13,
	ramiframload_14,
	ramiframload_15,
	ramiframload_16,
	ramiframload_17,
	ramiframload_18,
	ramiframload_19,
	ramiframload_20,
	ramiframload_21,
	ramiframload_22,
	ramiframload_23,
	ramiframload_24,
	ramiframload_25,
	ramiframload_26,
	ramiframload_27,
	ramiframload_28,
	ramiframload_29,
	ramiframload_30,
	ramiframload_31,
	plif_exmemrdat2_l_0,
	plif_exmemrdat2_l_1,
	plif_exmemrdat2_l_2,
	plif_exmemrdat2_l_3,
	plif_exmemrdat2_l_4,
	plif_exmemrdat2_l_5,
	plif_exmemrdat2_l_6,
	plif_exmemrdat2_l_7,
	plif_exmemrdat2_l_8,
	plif_exmemrdat2_l_9,
	plif_exmemrdat2_l_10,
	plif_exmemrdat2_l_11,
	plif_exmemrdat2_l_12,
	plif_exmemrdat2_l_13,
	plif_exmemrdat2_l_14,
	plif_exmemrdat2_l_15,
	plif_exmemrdat2_l_16,
	plif_exmemrdat2_l_17,
	plif_exmemrdat2_l_18,
	plif_exmemrdat2_l_19,
	plif_exmemrdat2_l_20,
	plif_exmemrdat2_l_21,
	plif_exmemrdat2_l_22,
	plif_exmemrdat2_l_23,
	plif_exmemrdat2_l_24,
	plif_exmemrdat2_l_25,
	plif_exmemrdat2_l_26,
	plif_exmemrdat2_l_27,
	plif_exmemrdat2_l_28,
	plif_exmemrdat2_l_29,
	plif_exmemrdat2_l_30,
	plif_exmemrdat2_l_31,
	nRST,
	CLK,
	nRST1,
	devpor,
	devclrn,
	devoe);
output 	PCreg_1;
output 	PCreg_0;
output 	plif_exmemhlt_l;
output 	plif_exmemporto_l_1;
output 	plif_exmemdmemWEN_l;
output 	plif_exmemdmemREN_l;
output 	plif_exmemporto_l_0;
output 	plif_exmemporto_l_3;
output 	PCreg_3;
output 	plif_exmemporto_l_2;
output 	PCreg_2;
output 	plif_exmemporto_l_5;
output 	PCreg_5;
output 	plif_exmemporto_l_4;
output 	PCreg_4;
output 	plif_exmemporto_l_7;
output 	PCreg_7;
output 	plif_exmemporto_l_6;
output 	PCreg_6;
output 	plif_exmemporto_l_9;
output 	PCreg_9;
output 	plif_exmemporto_l_8;
output 	PCreg_8;
output 	plif_exmemporto_l_11;
output 	PCreg_11;
output 	plif_exmemporto_l_10;
output 	PCreg_10;
output 	plif_exmemporto_l_13;
output 	PCreg_13;
output 	plif_exmemporto_l_12;
output 	PCreg_12;
output 	plif_exmemporto_l_15;
output 	PCreg_15;
output 	plif_exmemporto_l_14;
output 	PCreg_14;
output 	plif_exmemporto_l_17;
output 	PCreg_17;
output 	plif_exmemporto_l_16;
output 	PCreg_16;
output 	plif_exmemporto_l_19;
output 	PCreg_19;
output 	plif_exmemporto_l_18;
output 	PCreg_18;
output 	plif_exmemporto_l_21;
output 	PCreg_21;
output 	plif_exmemporto_l_20;
output 	PCreg_20;
output 	plif_exmemporto_l_23;
output 	PCreg_23;
output 	plif_exmemporto_l_22;
output 	PCreg_22;
output 	plif_exmemporto_l_25;
output 	PCreg_25;
output 	plif_exmemporto_l_24;
output 	PCreg_24;
output 	plif_exmemporto_l_27;
output 	PCreg_27;
output 	plif_exmemporto_l_26;
output 	PCreg_26;
output 	plif_exmemporto_l_29;
output 	PCreg_29;
output 	plif_exmemporto_l_28;
output 	PCreg_28;
output 	plif_exmemporto_l_31;
output 	PCreg_31;
output 	plif_exmemporto_l_30;
output 	PCreg_30;
output 	dpifimemREN;
input 	always1;
input 	ramiframload_0;
input 	ramiframload_1;
input 	ramiframload_2;
input 	ramiframload_3;
input 	ramiframload_4;
input 	ramiframload_5;
input 	ramiframload_6;
input 	ramiframload_7;
input 	ramiframload_8;
input 	ramiframload_9;
input 	ramiframload_10;
input 	ramiframload_11;
input 	ramiframload_12;
input 	ramiframload_13;
input 	ramiframload_14;
input 	ramiframload_15;
input 	ramiframload_16;
input 	ramiframload_17;
input 	ramiframload_18;
input 	ramiframload_19;
input 	ramiframload_20;
input 	ramiframload_21;
input 	ramiframload_22;
input 	ramiframload_23;
input 	ramiframload_24;
input 	ramiframload_25;
input 	ramiframload_26;
input 	ramiframload_27;
input 	ramiframload_28;
input 	ramiframload_29;
input 	ramiframload_30;
input 	ramiframload_31;
output 	plif_exmemrdat2_l_0;
output 	plif_exmemrdat2_l_1;
output 	plif_exmemrdat2_l_2;
output 	plif_exmemrdat2_l_3;
output 	plif_exmemrdat2_l_4;
output 	plif_exmemrdat2_l_5;
output 	plif_exmemrdat2_l_6;
output 	plif_exmemrdat2_l_7;
output 	plif_exmemrdat2_l_8;
output 	plif_exmemrdat2_l_9;
output 	plif_exmemrdat2_l_10;
output 	plif_exmemrdat2_l_11;
output 	plif_exmemrdat2_l_12;
output 	plif_exmemrdat2_l_13;
output 	plif_exmemrdat2_l_14;
output 	plif_exmemrdat2_l_15;
output 	plif_exmemrdat2_l_16;
output 	plif_exmemrdat2_l_17;
output 	plif_exmemrdat2_l_18;
output 	plif_exmemrdat2_l_19;
output 	plif_exmemrdat2_l_20;
output 	plif_exmemrdat2_l_21;
output 	plif_exmemrdat2_l_22;
output 	plif_exmemrdat2_l_23;
output 	plif_exmemrdat2_l_24;
output 	plif_exmemrdat2_l_25;
output 	plif_exmemrdat2_l_26;
output 	plif_exmemrdat2_l_27;
output 	plif_exmemrdat2_l_28;
output 	plif_exmemrdat2_l_29;
output 	plif_exmemrdat2_l_30;
output 	plif_exmemrdat2_l_31;
input 	nRST;
input 	CLK;
input 	nRST1;

// Design Ports Information

input 	devpor;
input 	devclrn;
input 	devoe;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
assign unknown = 1'bx;

wire \CC|always0~0_combout ;
wire \CC|ccif.iwait[0]~2_combout ;
wire [31:0] \CM|instr ;


memory_control CC(
	.plif_exmemdmemWEN_l(plif_exmemdmemWEN_l),
	.plif_exmemdmemREN_l(plif_exmemdmemREN_l),
	.dpifimemREN(dpifimemREN),
	.always1(always1),
	.always0(\CC|always0~0_combout ),
	.ccifiwait_0(\CC|ccif.iwait[0]~2_combout ),
	.devpor(devpor),
	.devclrn(devclrn),
	.devoe(devoe));

caches CM(
	.ramiframload_0(ramiframload_0),
	.ramiframload_1(ramiframload_1),
	.ramiframload_2(ramiframload_2),
	.ramiframload_3(ramiframload_3),
	.ramiframload_4(ramiframload_4),
	.ramiframload_5(ramiframload_5),
	.ramiframload_6(ramiframload_6),
	.ramiframload_7(ramiframload_7),
	.ramiframload_8(ramiframload_8),
	.ramiframload_9(ramiframload_9),
	.ramiframload_10(ramiframload_10),
	.ramiframload_11(ramiframload_11),
	.ramiframload_12(ramiframload_12),
	.ramiframload_13(ramiframload_13),
	.ramiframload_14(ramiframload_14),
	.ramiframload_15(ramiframload_15),
	.ramiframload_16(ramiframload_16),
	.ramiframload_17(ramiframload_17),
	.ramiframload_18(ramiframload_18),
	.ramiframload_19(ramiframload_19),
	.ramiframload_20(ramiframload_20),
	.ramiframload_21(ramiframload_21),
	.ramiframload_22(ramiframload_22),
	.ramiframload_23(ramiframload_23),
	.ramiframload_24(ramiframload_24),
	.ramiframload_25(ramiframload_25),
	.ramiframload_26(ramiframload_26),
	.ramiframload_27(ramiframload_27),
	.ramiframload_28(ramiframload_28),
	.ramiframload_29(ramiframload_29),
	.ramiframload_30(ramiframload_30),
	.ramiframload_31(ramiframload_31),
	.instr_31(\CM|instr [31]),
	.instr_29(\CM|instr [29]),
	.instr_27(\CM|instr [27]),
	.instr_26(\CM|instr [26]),
	.instr_28(\CM|instr [28]),
	.instr_30(\CM|instr [30]),
	.instr_5(\CM|instr [5]),
	.instr_1(\CM|instr [1]),
	.instr_0(\CM|instr [0]),
	.instr_2(\CM|instr [2]),
	.instr_3(\CM|instr [3]),
	.instr_4(\CM|instr [4]),
	.instr_22(\CM|instr [22]),
	.instr_21(\CM|instr [21]),
	.instr_24(\CM|instr [24]),
	.instr_23(\CM|instr [23]),
	.instr_25(\CM|instr [25]),
	.instr_17(\CM|instr [17]),
	.instr_16(\CM|instr [16]),
	.instr_19(\CM|instr [19]),
	.instr_18(\CM|instr [18]),
	.instr_20(\CM|instr [20]),
	.instr_15(\CM|instr [15]),
	.instr_14(\CM|instr [14]),
	.instr_13(\CM|instr [13]),
	.instr_12(\CM|instr [12]),
	.instr_11(\CM|instr [11]),
	.instr_10(\CM|instr [10]),
	.instr_9(\CM|instr [9]),
	.instr_8(\CM|instr [8]),
	.instr_7(\CM|instr [7]),
	.instr_6(\CM|instr [6]),
	.ccifiwait_0(\CC|ccif.iwait[0]~2_combout ),
	.nRST(nRST),
	.CLK(CLK),
	.devpor(devpor),
	.devclrn(devclrn),
	.devoe(devoe));

datapath DP(
	.PCreg_1(PCreg_1),
	.PCreg_0(PCreg_0),
	.plif_exmemhlt_l(plif_exmemhlt_l),
	.plif_exmemporto_l_1(plif_exmemporto_l_1),
	.plif_exmemdmemWEN_l(plif_exmemdmemWEN_l),
	.plif_exmemdmemREN_l(plif_exmemdmemREN_l),
	.plif_exmemporto_l_0(plif_exmemporto_l_0),
	.plif_exmemporto_l_3(plif_exmemporto_l_3),
	.PCreg_3(PCreg_3),
	.plif_exmemporto_l_2(plif_exmemporto_l_2),
	.PCreg_2(PCreg_2),
	.plif_exmemporto_l_5(plif_exmemporto_l_5),
	.PCreg_5(PCreg_5),
	.plif_exmemporto_l_4(plif_exmemporto_l_4),
	.PCreg_4(PCreg_4),
	.plif_exmemporto_l_7(plif_exmemporto_l_7),
	.PCreg_7(PCreg_7),
	.plif_exmemporto_l_6(plif_exmemporto_l_6),
	.PCreg_6(PCreg_6),
	.plif_exmemporto_l_9(plif_exmemporto_l_9),
	.PCreg_9(PCreg_9),
	.plif_exmemporto_l_8(plif_exmemporto_l_8),
	.PCreg_8(PCreg_8),
	.plif_exmemporto_l_11(plif_exmemporto_l_11),
	.PCreg_11(PCreg_11),
	.plif_exmemporto_l_10(plif_exmemporto_l_10),
	.PCreg_10(PCreg_10),
	.plif_exmemporto_l_13(plif_exmemporto_l_13),
	.PCreg_13(PCreg_13),
	.plif_exmemporto_l_12(plif_exmemporto_l_12),
	.PCreg_12(PCreg_12),
	.plif_exmemporto_l_15(plif_exmemporto_l_15),
	.PCreg_15(PCreg_15),
	.plif_exmemporto_l_14(plif_exmemporto_l_14),
	.PCreg_14(PCreg_14),
	.plif_exmemporto_l_17(plif_exmemporto_l_17),
	.PCreg_17(PCreg_17),
	.plif_exmemporto_l_16(plif_exmemporto_l_16),
	.PCreg_16(PCreg_16),
	.plif_exmemporto_l_19(plif_exmemporto_l_19),
	.PCreg_19(PCreg_19),
	.plif_exmemporto_l_18(plif_exmemporto_l_18),
	.PCreg_18(PCreg_18),
	.plif_exmemporto_l_21(plif_exmemporto_l_21),
	.PCreg_21(PCreg_21),
	.plif_exmemporto_l_20(plif_exmemporto_l_20),
	.PCreg_20(PCreg_20),
	.plif_exmemporto_l_23(plif_exmemporto_l_23),
	.PCreg_23(PCreg_23),
	.plif_exmemporto_l_22(plif_exmemporto_l_22),
	.PCreg_22(PCreg_22),
	.plif_exmemporto_l_25(plif_exmemporto_l_25),
	.PCreg_25(PCreg_25),
	.plif_exmemporto_l_24(plif_exmemporto_l_24),
	.PCreg_24(PCreg_24),
	.plif_exmemporto_l_27(plif_exmemporto_l_27),
	.PCreg_27(PCreg_27),
	.plif_exmemporto_l_26(plif_exmemporto_l_26),
	.PCreg_26(PCreg_26),
	.plif_exmemporto_l_29(plif_exmemporto_l_29),
	.PCreg_29(PCreg_29),
	.plif_exmemporto_l_28(plif_exmemporto_l_28),
	.PCreg_28(PCreg_28),
	.plif_exmemporto_l_31(plif_exmemporto_l_31),
	.PCreg_31(PCreg_31),
	.plif_exmemporto_l_30(plif_exmemporto_l_30),
	.PCreg_30(PCreg_30),
	.dpifimemREN(dpifimemREN),
	.always1(always1),
	.ramiframload_0(ramiframload_0),
	.ramiframload_1(ramiframload_1),
	.ramiframload_2(ramiframload_2),
	.ramiframload_3(ramiframload_3),
	.ramiframload_4(ramiframload_4),
	.ramiframload_5(ramiframload_5),
	.ramiframload_6(ramiframload_6),
	.ramiframload_7(ramiframload_7),
	.ramiframload_8(ramiframload_8),
	.ramiframload_9(ramiframload_9),
	.ramiframload_10(ramiframload_10),
	.ramiframload_11(ramiframload_11),
	.ramiframload_12(ramiframload_12),
	.ramiframload_13(ramiframload_13),
	.ramiframload_14(ramiframload_14),
	.ramiframload_15(ramiframload_15),
	.ramiframload_16(ramiframload_16),
	.ramiframload_17(ramiframload_17),
	.ramiframload_18(ramiframload_18),
	.ramiframload_19(ramiframload_19),
	.ramiframload_20(ramiframload_20),
	.ramiframload_21(ramiframload_21),
	.ramiframload_22(ramiframload_22),
	.ramiframload_23(ramiframload_23),
	.ramiframload_24(ramiframload_24),
	.ramiframload_25(ramiframload_25),
	.ramiframload_26(ramiframload_26),
	.ramiframload_27(ramiframload_27),
	.ramiframload_28(ramiframload_28),
	.ramiframload_29(ramiframload_29),
	.ramiframload_30(ramiframload_30),
	.ramiframload_31(ramiframload_31),
	.always0(\CC|always0~0_combout ),
	.plif_exmemrdat2_l_0(plif_exmemrdat2_l_0),
	.plif_exmemrdat2_l_1(plif_exmemrdat2_l_1),
	.plif_exmemrdat2_l_2(plif_exmemrdat2_l_2),
	.plif_exmemrdat2_l_3(plif_exmemrdat2_l_3),
	.plif_exmemrdat2_l_4(plif_exmemrdat2_l_4),
	.plif_exmemrdat2_l_5(plif_exmemrdat2_l_5),
	.plif_exmemrdat2_l_6(plif_exmemrdat2_l_6),
	.plif_exmemrdat2_l_7(plif_exmemrdat2_l_7),
	.plif_exmemrdat2_l_8(plif_exmemrdat2_l_8),
	.plif_exmemrdat2_l_9(plif_exmemrdat2_l_9),
	.plif_exmemrdat2_l_10(plif_exmemrdat2_l_10),
	.plif_exmemrdat2_l_11(plif_exmemrdat2_l_11),
	.plif_exmemrdat2_l_12(plif_exmemrdat2_l_12),
	.plif_exmemrdat2_l_13(plif_exmemrdat2_l_13),
	.plif_exmemrdat2_l_14(plif_exmemrdat2_l_14),
	.plif_exmemrdat2_l_15(plif_exmemrdat2_l_15),
	.plif_exmemrdat2_l_16(plif_exmemrdat2_l_16),
	.plif_exmemrdat2_l_17(plif_exmemrdat2_l_17),
	.plif_exmemrdat2_l_18(plif_exmemrdat2_l_18),
	.plif_exmemrdat2_l_19(plif_exmemrdat2_l_19),
	.plif_exmemrdat2_l_20(plif_exmemrdat2_l_20),
	.plif_exmemrdat2_l_21(plif_exmemrdat2_l_21),
	.plif_exmemrdat2_l_22(plif_exmemrdat2_l_22),
	.plif_exmemrdat2_l_23(plif_exmemrdat2_l_23),
	.plif_exmemrdat2_l_24(plif_exmemrdat2_l_24),
	.plif_exmemrdat2_l_25(plif_exmemrdat2_l_25),
	.plif_exmemrdat2_l_26(plif_exmemrdat2_l_26),
	.plif_exmemrdat2_l_27(plif_exmemrdat2_l_27),
	.plif_exmemrdat2_l_28(plif_exmemrdat2_l_28),
	.plif_exmemrdat2_l_29(plif_exmemrdat2_l_29),
	.plif_exmemrdat2_l_30(plif_exmemrdat2_l_30),
	.plif_exmemrdat2_l_31(plif_exmemrdat2_l_31),
	.instr_31(\CM|instr [31]),
	.instr_29(\CM|instr [29]),
	.instr_27(\CM|instr [27]),
	.instr_26(\CM|instr [26]),
	.instr_28(\CM|instr [28]),
	.instr_30(\CM|instr [30]),
	.instr_5(\CM|instr [5]),
	.instr_1(\CM|instr [1]),
	.instr_0(\CM|instr [0]),
	.instr_2(\CM|instr [2]),
	.instr_3(\CM|instr [3]),
	.instr_4(\CM|instr [4]),
	.instr_22(\CM|instr [22]),
	.instr_21(\CM|instr [21]),
	.instr_24(\CM|instr [24]),
	.instr_23(\CM|instr [23]),
	.instr_25(\CM|instr [25]),
	.instr_17(\CM|instr [17]),
	.instr_16(\CM|instr [16]),
	.instr_19(\CM|instr [19]),
	.instr_18(\CM|instr [18]),
	.instr_20(\CM|instr [20]),
	.instr_15(\CM|instr [15]),
	.instr_14(\CM|instr [14]),
	.instr_13(\CM|instr [13]),
	.instr_12(\CM|instr [12]),
	.instr_11(\CM|instr [11]),
	.instr_10(\CM|instr [10]),
	.instr_9(\CM|instr [9]),
	.instr_8(\CM|instr [8]),
	.instr_7(\CM|instr [7]),
	.instr_6(\CM|instr [6]),
	.ccifiwait_0(\CC|ccif.iwait[0]~2_combout ),
	.CLK(CLK),
	.nRST(nRST1),
	.devpor(devpor),
	.devclrn(devclrn),
	.devoe(devoe));

endmodule

module caches (
	ramiframload_0,
	ramiframload_1,
	ramiframload_2,
	ramiframload_3,
	ramiframload_4,
	ramiframload_5,
	ramiframload_6,
	ramiframload_7,
	ramiframload_8,
	ramiframload_9,
	ramiframload_10,
	ramiframload_11,
	ramiframload_12,
	ramiframload_13,
	ramiframload_14,
	ramiframload_15,
	ramiframload_16,
	ramiframload_17,
	ramiframload_18,
	ramiframload_19,
	ramiframload_20,
	ramiframload_21,
	ramiframload_22,
	ramiframload_23,
	ramiframload_24,
	ramiframload_25,
	ramiframload_26,
	ramiframload_27,
	ramiframload_28,
	ramiframload_29,
	ramiframload_30,
	ramiframload_31,
	instr_31,
	instr_29,
	instr_27,
	instr_26,
	instr_28,
	instr_30,
	instr_5,
	instr_1,
	instr_0,
	instr_2,
	instr_3,
	instr_4,
	instr_22,
	instr_21,
	instr_24,
	instr_23,
	instr_25,
	instr_17,
	instr_16,
	instr_19,
	instr_18,
	instr_20,
	instr_15,
	instr_14,
	instr_13,
	instr_12,
	instr_11,
	instr_10,
	instr_9,
	instr_8,
	instr_7,
	instr_6,
	ccifiwait_0,
	nRST,
	CLK,
	devpor,
	devclrn,
	devoe);
input 	ramiframload_0;
input 	ramiframload_1;
input 	ramiframload_2;
input 	ramiframload_3;
input 	ramiframload_4;
input 	ramiframload_5;
input 	ramiframload_6;
input 	ramiframload_7;
input 	ramiframload_8;
input 	ramiframload_9;
input 	ramiframload_10;
input 	ramiframload_11;
input 	ramiframload_12;
input 	ramiframload_13;
input 	ramiframload_14;
input 	ramiframload_15;
input 	ramiframload_16;
input 	ramiframload_17;
input 	ramiframload_18;
input 	ramiframload_19;
input 	ramiframload_20;
input 	ramiframload_21;
input 	ramiframload_22;
input 	ramiframload_23;
input 	ramiframload_24;
input 	ramiframload_25;
input 	ramiframload_26;
input 	ramiframload_27;
input 	ramiframload_28;
input 	ramiframload_29;
input 	ramiframload_30;
input 	ramiframload_31;
output 	instr_31;
output 	instr_29;
output 	instr_27;
output 	instr_26;
output 	instr_28;
output 	instr_30;
output 	instr_5;
output 	instr_1;
output 	instr_0;
output 	instr_2;
output 	instr_3;
output 	instr_4;
output 	instr_22;
output 	instr_21;
output 	instr_24;
output 	instr_23;
output 	instr_25;
output 	instr_17;
output 	instr_16;
output 	instr_19;
output 	instr_18;
output 	instr_20;
output 	instr_15;
output 	instr_14;
output 	instr_13;
output 	instr_12;
output 	instr_11;
output 	instr_10;
output 	instr_9;
output 	instr_8;
output 	instr_7;
output 	instr_6;
input 	ccifiwait_0;
input 	nRST;
input 	CLK;

// Design Ports Information

input 	devpor;
input 	devclrn;
input 	devoe;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
assign unknown = 1'bx;

wire \instr~0_combout ;
wire \instr~1_combout ;
wire \instr[29]~feeder_combout ;
wire \instr~2_combout ;
wire \instr[27]~feeder_combout ;
wire \instr~3_combout ;
wire \instr[26]~feeder_combout ;
wire \instr~4_combout ;
wire \instr~5_combout ;
wire \instr[30]~feeder_combout ;
wire \instr~6_combout ;
wire \instr[5]~feeder_combout ;
wire \instr~7_combout ;
wire \instr[1]~feeder_combout ;
wire \instr~8_combout ;
wire \instr~9_combout ;
wire \instr[2]~feeder_combout ;
wire \instr~10_combout ;
wire \instr[3]~feeder_combout ;
wire \instr~11_combout ;
wire \instr~12_combout ;
wire \instr~13_combout ;
wire \instr[21]~feeder_combout ;
wire \instr~14_combout ;
wire \instr~15_combout ;
wire \instr[23]~feeder_combout ;
wire \instr~16_combout ;
wire \instr[25]~feeder_combout ;
wire \instr~17_combout ;
wire \instr[17]~feeder_combout ;
wire \instr~18_combout ;
wire \instr[16]~feeder_combout ;
wire \instr~19_combout ;
wire \instr[19]~feeder_combout ;
wire \instr~20_combout ;
wire \instr~21_combout ;
wire \instr[20]~feeder_combout ;
wire \instr~22_combout ;
wire \instr[15]~feeder_combout ;
wire \instr~23_combout ;
wire \instr[14]~feeder_combout ;
wire \instr~24_combout ;
wire \instr~25_combout ;
wire \instr[12]~feeder_combout ;
wire \instr~26_combout ;
wire \instr[11]~feeder_combout ;
wire \instr~27_combout ;
wire \instr~28_combout ;
wire \instr[9]~feeder_combout ;
wire \instr~29_combout ;
wire \instr[8]~feeder_combout ;
wire \instr~30_combout ;
wire \instr[7]~feeder_combout ;
wire \instr~31_combout ;
wire \instr[6]~feeder_combout ;


// Location: FF_X54_Y30_N17
dffeas \instr[31] (
	.clk(CLK),
	.d(gnd),
	.asdata(\instr~0_combout ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(instr_31),
	.prn(vcc));
// synopsys translate_off
defparam \instr[31] .is_wysiwyg = "true";
defparam \instr[31] .power_up = "low";
// synopsys translate_on

// Location: FF_X54_Y30_N7
dffeas \instr[29] (
	.clk(CLK),
	.d(\instr[29]~feeder_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(instr_29),
	.prn(vcc));
// synopsys translate_off
defparam \instr[29] .is_wysiwyg = "true";
defparam \instr[29] .power_up = "low";
// synopsys translate_on

// Location: FF_X54_Y30_N21
dffeas \instr[27] (
	.clk(CLK),
	.d(\instr[27]~feeder_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(instr_27),
	.prn(vcc));
// synopsys translate_off
defparam \instr[27] .is_wysiwyg = "true";
defparam \instr[27] .power_up = "low";
// synopsys translate_on

// Location: FF_X58_Y30_N5
dffeas \instr[26] (
	.clk(CLK),
	.d(\instr[26]~feeder_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(instr_26),
	.prn(vcc));
// synopsys translate_off
defparam \instr[26] .is_wysiwyg = "true";
defparam \instr[26] .power_up = "low";
// synopsys translate_on

// Location: FF_X58_Y30_N15
dffeas \instr[28] (
	.clk(CLK),
	.d(gnd),
	.asdata(\instr~4_combout ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(instr_28),
	.prn(vcc));
// synopsys translate_off
defparam \instr[28] .is_wysiwyg = "true";
defparam \instr[28] .power_up = "low";
// synopsys translate_on

// Location: FF_X54_Y30_N15
dffeas \instr[30] (
	.clk(CLK),
	.d(\instr[30]~feeder_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(instr_30),
	.prn(vcc));
// synopsys translate_off
defparam \instr[30] .is_wysiwyg = "true";
defparam \instr[30] .power_up = "low";
// synopsys translate_on

// Location: FF_X58_Y30_N9
dffeas \instr[5] (
	.clk(CLK),
	.d(\instr[5]~feeder_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(instr_5),
	.prn(vcc));
// synopsys translate_off
defparam \instr[5] .is_wysiwyg = "true";
defparam \instr[5] .power_up = "low";
// synopsys translate_on

// Location: FF_X55_Y30_N9
dffeas \instr[1] (
	.clk(CLK),
	.d(\instr[1]~feeder_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(instr_1),
	.prn(vcc));
// synopsys translate_off
defparam \instr[1] .is_wysiwyg = "true";
defparam \instr[1] .power_up = "low";
// synopsys translate_on

// Location: FF_X56_Y33_N23
dffeas \instr[0] (
	.clk(CLK),
	.d(gnd),
	.asdata(\instr~8_combout ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(instr_0),
	.prn(vcc));
// synopsys translate_off
defparam \instr[0] .is_wysiwyg = "true";
defparam \instr[0] .power_up = "low";
// synopsys translate_on

// Location: FF_X56_Y29_N5
dffeas \instr[2] (
	.clk(CLK),
	.d(\instr[2]~feeder_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(instr_2),
	.prn(vcc));
// synopsys translate_off
defparam \instr[2] .is_wysiwyg = "true";
defparam \instr[2] .power_up = "low";
// synopsys translate_on

// Location: FF_X55_Y30_N31
dffeas \instr[3] (
	.clk(CLK),
	.d(\instr[3]~feeder_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(instr_3),
	.prn(vcc));
// synopsys translate_off
defparam \instr[3] .is_wysiwyg = "true";
defparam \instr[3] .power_up = "low";
// synopsys translate_on

// Location: FF_X56_Y33_N11
dffeas \instr[4] (
	.clk(CLK),
	.d(gnd),
	.asdata(\instr~11_combout ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(instr_4),
	.prn(vcc));
// synopsys translate_off
defparam \instr[4] .is_wysiwyg = "true";
defparam \instr[4] .power_up = "low";
// synopsys translate_on

// Location: FF_X59_Y32_N27
dffeas \instr[22] (
	.clk(CLK),
	.d(gnd),
	.asdata(\instr~12_combout ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(instr_22),
	.prn(vcc));
// synopsys translate_off
defparam \instr[22] .is_wysiwyg = "true";
defparam \instr[22] .power_up = "low";
// synopsys translate_on

// Location: FF_X59_Y32_N9
dffeas \instr[21] (
	.clk(CLK),
	.d(\instr[21]~feeder_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(instr_21),
	.prn(vcc));
// synopsys translate_off
defparam \instr[21] .is_wysiwyg = "true";
defparam \instr[21] .power_up = "low";
// synopsys translate_on

// Location: FF_X59_Y32_N29
dffeas \instr[24] (
	.clk(CLK),
	.d(gnd),
	.asdata(\instr~14_combout ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(instr_24),
	.prn(vcc));
// synopsys translate_off
defparam \instr[24] .is_wysiwyg = "true";
defparam \instr[24] .power_up = "low";
// synopsys translate_on

// Location: FF_X59_Y32_N31
dffeas \instr[23] (
	.clk(CLK),
	.d(\instr[23]~feeder_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(instr_23),
	.prn(vcc));
// synopsys translate_off
defparam \instr[23] .is_wysiwyg = "true";
defparam \instr[23] .power_up = "low";
// synopsys translate_on

// Location: FF_X59_Y33_N5
dffeas \instr[25] (
	.clk(CLK),
	.d(\instr[25]~feeder_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(instr_25),
	.prn(vcc));
// synopsys translate_off
defparam \instr[25] .is_wysiwyg = "true";
defparam \instr[25] .power_up = "low";
// synopsys translate_on

// Location: FF_X59_Y31_N5
dffeas \instr[17] (
	.clk(CLK),
	.d(\instr[17]~feeder_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(instr_17),
	.prn(vcc));
// synopsys translate_off
defparam \instr[17] .is_wysiwyg = "true";
defparam \instr[17] .power_up = "low";
// synopsys translate_on

// Location: FF_X59_Y31_N27
dffeas \instr[16] (
	.clk(CLK),
	.d(\instr[16]~feeder_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(instr_16),
	.prn(vcc));
// synopsys translate_off
defparam \instr[16] .is_wysiwyg = "true";
defparam \instr[16] .power_up = "low";
// synopsys translate_on

// Location: FF_X59_Y33_N27
dffeas \instr[19] (
	.clk(CLK),
	.d(\instr[19]~feeder_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(instr_19),
	.prn(vcc));
// synopsys translate_off
defparam \instr[19] .is_wysiwyg = "true";
defparam \instr[19] .power_up = "low";
// synopsys translate_on

// Location: FF_X59_Y31_N9
dffeas \instr[18] (
	.clk(CLK),
	.d(gnd),
	.asdata(\instr~20_combout ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(instr_18),
	.prn(vcc));
// synopsys translate_off
defparam \instr[18] .is_wysiwyg = "true";
defparam \instr[18] .power_up = "low";
// synopsys translate_on

// Location: FF_X59_Y33_N9
dffeas \instr[20] (
	.clk(CLK),
	.d(\instr[20]~feeder_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(instr_20),
	.prn(vcc));
// synopsys translate_off
defparam \instr[20] .is_wysiwyg = "true";
defparam \instr[20] .power_up = "low";
// synopsys translate_on

// Location: FF_X59_Y33_N23
dffeas \instr[15] (
	.clk(CLK),
	.d(\instr[15]~feeder_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(instr_15),
	.prn(vcc));
// synopsys translate_off
defparam \instr[15] .is_wysiwyg = "true";
defparam \instr[15] .power_up = "low";
// synopsys translate_on

// Location: FF_X57_Y31_N15
dffeas \instr[14] (
	.clk(CLK),
	.d(\instr[14]~feeder_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(instr_14),
	.prn(vcc));
// synopsys translate_off
defparam \instr[14] .is_wysiwyg = "true";
defparam \instr[14] .power_up = "low";
// synopsys translate_on

// Location: FF_X56_Y33_N5
dffeas \instr[13] (
	.clk(CLK),
	.d(gnd),
	.asdata(\instr~24_combout ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(instr_13),
	.prn(vcc));
// synopsys translate_off
defparam \instr[13] .is_wysiwyg = "true";
defparam \instr[13] .power_up = "low";
// synopsys translate_on

// Location: FF_X57_Y31_N9
dffeas \instr[12] (
	.clk(CLK),
	.d(\instr[12]~feeder_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(instr_12),
	.prn(vcc));
// synopsys translate_off
defparam \instr[12] .is_wysiwyg = "true";
defparam \instr[12] .power_up = "low";
// synopsys translate_on

// Location: FF_X56_Y29_N7
dffeas \instr[11] (
	.clk(CLK),
	.d(\instr[11]~feeder_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(instr_11),
	.prn(vcc));
// synopsys translate_off
defparam \instr[11] .is_wysiwyg = "true";
defparam \instr[11] .power_up = "low";
// synopsys translate_on

// Location: FF_X58_Y30_N27
dffeas \instr[10] (
	.clk(CLK),
	.d(gnd),
	.asdata(\instr~27_combout ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(instr_10),
	.prn(vcc));
// synopsys translate_off
defparam \instr[10] .is_wysiwyg = "true";
defparam \instr[10] .power_up = "low";
// synopsys translate_on

// Location: FF_X57_Y31_N31
dffeas \instr[9] (
	.clk(CLK),
	.d(\instr[9]~feeder_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(instr_9),
	.prn(vcc));
// synopsys translate_off
defparam \instr[9] .is_wysiwyg = "true";
defparam \instr[9] .power_up = "low";
// synopsys translate_on

// Location: FF_X56_Y29_N17
dffeas \instr[8] (
	.clk(CLK),
	.d(\instr[8]~feeder_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(instr_8),
	.prn(vcc));
// synopsys translate_off
defparam \instr[8] .is_wysiwyg = "true";
defparam \instr[8] .power_up = "low";
// synopsys translate_on

// Location: FF_X55_Y30_N5
dffeas \instr[7] (
	.clk(CLK),
	.d(\instr[7]~feeder_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(instr_7),
	.prn(vcc));
// synopsys translate_off
defparam \instr[7] .is_wysiwyg = "true";
defparam \instr[7] .power_up = "low";
// synopsys translate_on

// Location: FF_X55_Y30_N23
dffeas \instr[6] (
	.clk(CLK),
	.d(\instr[6]~feeder_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(instr_6),
	.prn(vcc));
// synopsys translate_off
defparam \instr[6] .is_wysiwyg = "true";
defparam \instr[6] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X54_Y30_N28
cycloneive_lcell_comb \instr~0 (
// Equation(s):
// \instr~0_combout  = (\nRST~input_o  & ((ccifiwait_0 & ((instr_31))) # (!ccifiwait_0 & (ramiframload_31))))

	.dataa(ramiframload_31),
	.datab(instr_31),
	.datac(ccifiwait_0),
	.datad(nRST),
	.cin(gnd),
	.combout(\instr~0_combout ),
	.cout());
// synopsys translate_off
defparam \instr~0 .lut_mask = 16'hCA00;
defparam \instr~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y30_N18
cycloneive_lcell_comb \instr~1 (
// Equation(s):
// \instr~1_combout  = (\nRST~input_o  & ((ccifiwait_0 & (instr_29)) # (!ccifiwait_0 & ((ramiframload_29)))))

	.dataa(instr_29),
	.datab(nRST),
	.datac(ccifiwait_0),
	.datad(ramiframload_29),
	.cin(gnd),
	.combout(\instr~1_combout ),
	.cout());
// synopsys translate_off
defparam \instr~1 .lut_mask = 16'h8C80;
defparam \instr~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y30_N6
cycloneive_lcell_comb \instr[29]~feeder (
// Equation(s):
// \instr[29]~feeder_combout  = \instr~1_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(\instr~1_combout ),
	.cin(gnd),
	.combout(\instr[29]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \instr[29]~feeder .lut_mask = 16'hFF00;
defparam \instr[29]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y30_N0
cycloneive_lcell_comb \instr~2 (
// Equation(s):
// \instr~2_combout  = (\nRST~input_o  & ((ccifiwait_0 & ((instr_27))) # (!ccifiwait_0 & (ramiframload_27))))

	.dataa(ramiframload_27),
	.datab(instr_27),
	.datac(ccifiwait_0),
	.datad(nRST),
	.cin(gnd),
	.combout(\instr~2_combout ),
	.cout());
// synopsys translate_off
defparam \instr~2 .lut_mask = 16'hCA00;
defparam \instr~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y30_N20
cycloneive_lcell_comb \instr[27]~feeder (
// Equation(s):
// \instr[27]~feeder_combout  = \instr~2_combout 

	.dataa(gnd),
	.datab(\instr~2_combout ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\instr[27]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \instr[27]~feeder .lut_mask = 16'hCCCC;
defparam \instr[27]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y30_N0
cycloneive_lcell_comb \instr~3 (
// Equation(s):
// \instr~3_combout  = (\nRST~input_o  & ((ccifiwait_0 & ((instr_26))) # (!ccifiwait_0 & (ramiframload_26))))

	.dataa(nRST),
	.datab(ramiframload_26),
	.datac(ccifiwait_0),
	.datad(instr_26),
	.cin(gnd),
	.combout(\instr~3_combout ),
	.cout());
// synopsys translate_off
defparam \instr~3 .lut_mask = 16'hA808;
defparam \instr~3 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y30_N4
cycloneive_lcell_comb \instr[26]~feeder (
// Equation(s):
// \instr[26]~feeder_combout  = \instr~3_combout 

	.dataa(gnd),
	.datab(\instr~3_combout ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\instr[26]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \instr[26]~feeder .lut_mask = 16'hCCCC;
defparam \instr[26]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y30_N30
cycloneive_lcell_comb \instr~4 (
// Equation(s):
// \instr~4_combout  = (\nRST~input_o  & ((ccifiwait_0 & ((instr_28))) # (!ccifiwait_0 & (ramiframload_28))))

	.dataa(ramiframload_28),
	.datab(ccifiwait_0),
	.datac(nRST),
	.datad(instr_28),
	.cin(gnd),
	.combout(\instr~4_combout ),
	.cout());
// synopsys translate_off
defparam \instr~4 .lut_mask = 16'hE020;
defparam \instr~4 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y30_N2
cycloneive_lcell_comb \instr~5 (
// Equation(s):
// \instr~5_combout  = (\nRST~input_o  & ((ccifiwait_0 & (instr_30)) # (!ccifiwait_0 & ((ramiframload_30)))))

	.dataa(ccifiwait_0),
	.datab(instr_30),
	.datac(nRST),
	.datad(ramiframload_30),
	.cin(gnd),
	.combout(\instr~5_combout ),
	.cout());
// synopsys translate_off
defparam \instr~5 .lut_mask = 16'hD080;
defparam \instr~5 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y30_N14
cycloneive_lcell_comb \instr[30]~feeder (
// Equation(s):
// \instr[30]~feeder_combout  = \instr~5_combout 

	.dataa(\instr~5_combout ),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\instr[30]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \instr[30]~feeder .lut_mask = 16'hAAAA;
defparam \instr[30]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y30_N20
cycloneive_lcell_comb \instr~6 (
// Equation(s):
// \instr~6_combout  = (\nRST~input_o  & ((ccifiwait_0 & ((instr_5))) # (!ccifiwait_0 & (ramiframload_5))))

	.dataa(ramiframload_5),
	.datab(instr_5),
	.datac(nRST),
	.datad(ccifiwait_0),
	.cin(gnd),
	.combout(\instr~6_combout ),
	.cout());
// synopsys translate_off
defparam \instr~6 .lut_mask = 16'hC0A0;
defparam \instr~6 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y30_N8
cycloneive_lcell_comb \instr[5]~feeder (
// Equation(s):
// \instr[5]~feeder_combout  = \instr~6_combout 

	.dataa(gnd),
	.datab(\instr~6_combout ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\instr[5]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \instr[5]~feeder .lut_mask = 16'hCCCC;
defparam \instr[5]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y30_N0
cycloneive_lcell_comb \instr~7 (
// Equation(s):
// \instr~7_combout  = (\nRST~input_o  & ((ccifiwait_0 & ((instr_1))) # (!ccifiwait_0 & (ramiframload_1))))

	.dataa(ccifiwait_0),
	.datab(ramiframload_1),
	.datac(instr_1),
	.datad(nRST),
	.cin(gnd),
	.combout(\instr~7_combout ),
	.cout());
// synopsys translate_off
defparam \instr~7 .lut_mask = 16'hE400;
defparam \instr~7 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y30_N8
cycloneive_lcell_comb \instr[1]~feeder (
// Equation(s):
// \instr[1]~feeder_combout  = \instr~7_combout 

	.dataa(gnd),
	.datab(\instr~7_combout ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\instr[1]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \instr[1]~feeder .lut_mask = 16'hCCCC;
defparam \instr[1]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y33_N2
cycloneive_lcell_comb \instr~8 (
// Equation(s):
// \instr~8_combout  = (\nRST~input_o  & ((ccifiwait_0 & (instr_0)) # (!ccifiwait_0 & ((ramiframload_0)))))

	.dataa(nRST),
	.datab(ccifiwait_0),
	.datac(instr_0),
	.datad(ramiframload_0),
	.cin(gnd),
	.combout(\instr~8_combout ),
	.cout());
// synopsys translate_off
defparam \instr~8 .lut_mask = 16'hA280;
defparam \instr~8 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y29_N18
cycloneive_lcell_comb \instr~9 (
// Equation(s):
// \instr~9_combout  = (\nRST~input_o  & ((ccifiwait_0 & ((instr_2))) # (!ccifiwait_0 & (ramiframload_2))))

	.dataa(nRST),
	.datab(ramiframload_2),
	.datac(instr_2),
	.datad(ccifiwait_0),
	.cin(gnd),
	.combout(\instr~9_combout ),
	.cout());
// synopsys translate_off
defparam \instr~9 .lut_mask = 16'hA088;
defparam \instr~9 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y29_N4
cycloneive_lcell_comb \instr[2]~feeder (
// Equation(s):
// \instr[2]~feeder_combout  = \instr~9_combout 

	.dataa(gnd),
	.datab(\instr~9_combout ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\instr[2]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \instr[2]~feeder .lut_mask = 16'hCCCC;
defparam \instr[2]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y30_N14
cycloneive_lcell_comb \instr~10 (
// Equation(s):
// \instr~10_combout  = (\nRST~input_o  & ((ccifiwait_0 & ((instr_3))) # (!ccifiwait_0 & (ramiframload_3))))

	.dataa(ramiframload_3),
	.datab(nRST),
	.datac(instr_3),
	.datad(ccifiwait_0),
	.cin(gnd),
	.combout(\instr~10_combout ),
	.cout());
// synopsys translate_off
defparam \instr~10 .lut_mask = 16'hC088;
defparam \instr~10 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y30_N30
cycloneive_lcell_comb \instr[3]~feeder (
// Equation(s):
// \instr[3]~feeder_combout  = \instr~10_combout 

	.dataa(gnd),
	.datab(\instr~10_combout ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\instr[3]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \instr[3]~feeder .lut_mask = 16'hCCCC;
defparam \instr[3]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y33_N28
cycloneive_lcell_comb \instr~11 (
// Equation(s):
// \instr~11_combout  = (\nRST~input_o  & ((ccifiwait_0 & (instr_4)) # (!ccifiwait_0 & ((ramiframload_4)))))

	.dataa(instr_4),
	.datab(nRST),
	.datac(ramiframload_4),
	.datad(ccifiwait_0),
	.cin(gnd),
	.combout(\instr~11_combout ),
	.cout());
// synopsys translate_off
defparam \instr~11 .lut_mask = 16'h88C0;
defparam \instr~11 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y32_N4
cycloneive_lcell_comb \instr~12 (
// Equation(s):
// \instr~12_combout  = (\nRST~input_o  & ((ccifiwait_0 & (instr_22)) # (!ccifiwait_0 & ((ramiframload_22)))))

	.dataa(nRST),
	.datab(instr_22),
	.datac(ramiframload_22),
	.datad(ccifiwait_0),
	.cin(gnd),
	.combout(\instr~12_combout ),
	.cout());
// synopsys translate_off
defparam \instr~12 .lut_mask = 16'h88A0;
defparam \instr~12 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y32_N6
cycloneive_lcell_comb \instr~13 (
// Equation(s):
// \instr~13_combout  = (\nRST~input_o  & ((ccifiwait_0 & (instr_21)) # (!ccifiwait_0 & ((ramiframload_21)))))

	.dataa(nRST),
	.datab(ccifiwait_0),
	.datac(instr_21),
	.datad(ramiframload_21),
	.cin(gnd),
	.combout(\instr~13_combout ),
	.cout());
// synopsys translate_off
defparam \instr~13 .lut_mask = 16'hA280;
defparam \instr~13 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y32_N8
cycloneive_lcell_comb \instr[21]~feeder (
// Equation(s):
// \instr[21]~feeder_combout  = \instr~13_combout 

	.dataa(\instr~13_combout ),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\instr[21]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \instr[21]~feeder .lut_mask = 16'hAAAA;
defparam \instr[21]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y32_N12
cycloneive_lcell_comb \instr~14 (
// Equation(s):
// \instr~14_combout  = (\nRST~input_o  & ((ccifiwait_0 & (instr_24)) # (!ccifiwait_0 & ((ramiframload_24)))))

	.dataa(nRST),
	.datab(instr_24),
	.datac(ramiframload_24),
	.datad(ccifiwait_0),
	.cin(gnd),
	.combout(\instr~14_combout ),
	.cout());
// synopsys translate_off
defparam \instr~14 .lut_mask = 16'h88A0;
defparam \instr~14 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y32_N2
cycloneive_lcell_comb \instr~15 (
// Equation(s):
// \instr~15_combout  = (\nRST~input_o  & ((ccifiwait_0 & ((instr_23))) # (!ccifiwait_0 & (ramiframload_23))))

	.dataa(nRST),
	.datab(ramiframload_23),
	.datac(instr_23),
	.datad(ccifiwait_0),
	.cin(gnd),
	.combout(\instr~15_combout ),
	.cout());
// synopsys translate_off
defparam \instr~15 .lut_mask = 16'hA088;
defparam \instr~15 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y32_N30
cycloneive_lcell_comb \instr[23]~feeder (
// Equation(s):
// \instr[23]~feeder_combout  = \instr~15_combout 

	.dataa(gnd),
	.datab(\instr~15_combout ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\instr[23]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \instr[23]~feeder .lut_mask = 16'hCCCC;
defparam \instr[23]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y33_N24
cycloneive_lcell_comb \instr~16 (
// Equation(s):
// \instr~16_combout  = (\nRST~input_o  & ((ccifiwait_0 & (instr_25)) # (!ccifiwait_0 & ((ramiframload_25)))))

	.dataa(nRST),
	.datab(instr_25),
	.datac(ramiframload_25),
	.datad(ccifiwait_0),
	.cin(gnd),
	.combout(\instr~16_combout ),
	.cout());
// synopsys translate_off
defparam \instr~16 .lut_mask = 16'h88A0;
defparam \instr~16 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y33_N4
cycloneive_lcell_comb \instr[25]~feeder (
// Equation(s):
// \instr[25]~feeder_combout  = \instr~16_combout 

	.dataa(gnd),
	.datab(\instr~16_combout ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\instr[25]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \instr[25]~feeder .lut_mask = 16'hCCCC;
defparam \instr[25]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y31_N2
cycloneive_lcell_comb \instr~17 (
// Equation(s):
// \instr~17_combout  = (\nRST~input_o  & ((ccifiwait_0 & (instr_17)) # (!ccifiwait_0 & ((ramiframload_17)))))

	.dataa(nRST),
	.datab(instr_17),
	.datac(ramiframload_17),
	.datad(ccifiwait_0),
	.cin(gnd),
	.combout(\instr~17_combout ),
	.cout());
// synopsys translate_off
defparam \instr~17 .lut_mask = 16'h88A0;
defparam \instr~17 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y31_N4
cycloneive_lcell_comb \instr[17]~feeder (
// Equation(s):
// \instr[17]~feeder_combout  = \instr~17_combout 

	.dataa(gnd),
	.datab(\instr~17_combout ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\instr[17]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \instr[17]~feeder .lut_mask = 16'hCCCC;
defparam \instr[17]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y31_N12
cycloneive_lcell_comb \instr~18 (
// Equation(s):
// \instr~18_combout  = (\nRST~input_o  & ((ccifiwait_0 & ((instr_16))) # (!ccifiwait_0 & (ramiframload_16))))

	.dataa(nRST),
	.datab(ramiframload_16),
	.datac(instr_16),
	.datad(ccifiwait_0),
	.cin(gnd),
	.combout(\instr~18_combout ),
	.cout());
// synopsys translate_off
defparam \instr~18 .lut_mask = 16'hA088;
defparam \instr~18 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y31_N26
cycloneive_lcell_comb \instr[16]~feeder (
// Equation(s):
// \instr[16]~feeder_combout  = \instr~18_combout 

	.dataa(\instr~18_combout ),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\instr[16]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \instr[16]~feeder .lut_mask = 16'hAAAA;
defparam \instr[16]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y33_N2
cycloneive_lcell_comb \instr~19 (
// Equation(s):
// \instr~19_combout  = (\nRST~input_o  & ((ccifiwait_0 & ((instr_19))) # (!ccifiwait_0 & (ramiframload_19))))

	.dataa(nRST),
	.datab(ramiframload_19),
	.datac(instr_19),
	.datad(ccifiwait_0),
	.cin(gnd),
	.combout(\instr~19_combout ),
	.cout());
// synopsys translate_off
defparam \instr~19 .lut_mask = 16'hA088;
defparam \instr~19 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y33_N26
cycloneive_lcell_comb \instr[19]~feeder (
// Equation(s):
// \instr[19]~feeder_combout  = \instr~19_combout 

	.dataa(gnd),
	.datab(\instr~19_combout ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\instr[19]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \instr[19]~feeder .lut_mask = 16'hCCCC;
defparam \instr[19]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y31_N22
cycloneive_lcell_comb \instr~20 (
// Equation(s):
// \instr~20_combout  = (\nRST~input_o  & ((ccifiwait_0 & (instr_18)) # (!ccifiwait_0 & ((ramiframload_18)))))

	.dataa(nRST),
	.datab(instr_18),
	.datac(ccifiwait_0),
	.datad(ramiframload_18),
	.cin(gnd),
	.combout(\instr~20_combout ),
	.cout());
// synopsys translate_off
defparam \instr~20 .lut_mask = 16'h8A80;
defparam \instr~20 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y33_N28
cycloneive_lcell_comb \instr~21 (
// Equation(s):
// \instr~21_combout  = (\nRST~input_o  & ((ccifiwait_0 & ((instr_20))) # (!ccifiwait_0 & (ramiframload_20))))

	.dataa(nRST),
	.datab(ramiframload_20),
	.datac(instr_20),
	.datad(ccifiwait_0),
	.cin(gnd),
	.combout(\instr~21_combout ),
	.cout());
// synopsys translate_off
defparam \instr~21 .lut_mask = 16'hA088;
defparam \instr~21 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y33_N8
cycloneive_lcell_comb \instr[20]~feeder (
// Equation(s):
// \instr[20]~feeder_combout  = \instr~21_combout 

	.dataa(gnd),
	.datab(\instr~21_combout ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\instr[20]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \instr[20]~feeder .lut_mask = 16'hCCCC;
defparam \instr[20]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y33_N10
cycloneive_lcell_comb \instr~22 (
// Equation(s):
// \instr~22_combout  = (\nRST~input_o  & ((ccifiwait_0 & ((instr_15))) # (!ccifiwait_0 & (ramiframload_15))))

	.dataa(nRST),
	.datab(ramiframload_15),
	.datac(instr_15),
	.datad(ccifiwait_0),
	.cin(gnd),
	.combout(\instr~22_combout ),
	.cout());
// synopsys translate_off
defparam \instr~22 .lut_mask = 16'hA088;
defparam \instr~22 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y33_N22
cycloneive_lcell_comb \instr[15]~feeder (
// Equation(s):
// \instr[15]~feeder_combout  = \instr~22_combout 

	.dataa(\instr~22_combout ),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\instr[15]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \instr[15]~feeder .lut_mask = 16'hAAAA;
defparam \instr[15]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y31_N26
cycloneive_lcell_comb \instr~23 (
// Equation(s):
// \instr~23_combout  = (\nRST~input_o  & ((ccifiwait_0 & (instr_14)) # (!ccifiwait_0 & ((ramiframload_14)))))

	.dataa(nRST),
	.datab(instr_14),
	.datac(ccifiwait_0),
	.datad(ramiframload_14),
	.cin(gnd),
	.combout(\instr~23_combout ),
	.cout());
// synopsys translate_off
defparam \instr~23 .lut_mask = 16'h8A80;
defparam \instr~23 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y31_N14
cycloneive_lcell_comb \instr[14]~feeder (
// Equation(s):
// \instr[14]~feeder_combout  = \instr~23_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(\instr~23_combout ),
	.datad(gnd),
	.cin(gnd),
	.combout(\instr[14]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \instr[14]~feeder .lut_mask = 16'hF0F0;
defparam \instr[14]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y33_N14
cycloneive_lcell_comb \instr~24 (
// Equation(s):
// \instr~24_combout  = (\nRST~input_o  & ((ccifiwait_0 & (instr_13)) # (!ccifiwait_0 & ((ramiframload_13)))))

	.dataa(nRST),
	.datab(ccifiwait_0),
	.datac(instr_13),
	.datad(ramiframload_13),
	.cin(gnd),
	.combout(\instr~24_combout ),
	.cout());
// synopsys translate_off
defparam \instr~24 .lut_mask = 16'hA280;
defparam \instr~24 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y31_N18
cycloneive_lcell_comb \instr~25 (
// Equation(s):
// \instr~25_combout  = (\nRST~input_o  & ((ccifiwait_0 & (instr_12)) # (!ccifiwait_0 & ((ramiframload_12)))))

	.dataa(nRST),
	.datab(instr_12),
	.datac(ccifiwait_0),
	.datad(ramiframload_12),
	.cin(gnd),
	.combout(\instr~25_combout ),
	.cout());
// synopsys translate_off
defparam \instr~25 .lut_mask = 16'h8A80;
defparam \instr~25 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y31_N8
cycloneive_lcell_comb \instr[12]~feeder (
// Equation(s):
// \instr[12]~feeder_combout  = \instr~25_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(\instr~25_combout ),
	.cin(gnd),
	.combout(\instr[12]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \instr[12]~feeder .lut_mask = 16'hFF00;
defparam \instr[12]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y29_N12
cycloneive_lcell_comb \instr~26 (
// Equation(s):
// \instr~26_combout  = (\nRST~input_o  & ((ccifiwait_0 & ((instr_11))) # (!ccifiwait_0 & (ramiframload_11))))

	.dataa(nRST),
	.datab(ramiframload_11),
	.datac(instr_11),
	.datad(ccifiwait_0),
	.cin(gnd),
	.combout(\instr~26_combout ),
	.cout());
// synopsys translate_off
defparam \instr~26 .lut_mask = 16'hA088;
defparam \instr~26 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y29_N6
cycloneive_lcell_comb \instr[11]~feeder (
// Equation(s):
// \instr[11]~feeder_combout  = \instr~26_combout 

	.dataa(\instr~26_combout ),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\instr[11]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \instr[11]~feeder .lut_mask = 16'hAAAA;
defparam \instr[11]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y30_N22
cycloneive_lcell_comb \instr~27 (
// Equation(s):
// \instr~27_combout  = (\nRST~input_o  & ((ccifiwait_0 & (instr_10)) # (!ccifiwait_0 & ((ramiframload_10)))))

	.dataa(instr_10),
	.datab(ccifiwait_0),
	.datac(nRST),
	.datad(ramiframload_10),
	.cin(gnd),
	.combout(\instr~27_combout ),
	.cout());
// synopsys translate_off
defparam \instr~27 .lut_mask = 16'hB080;
defparam \instr~27 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y31_N0
cycloneive_lcell_comb \instr~28 (
// Equation(s):
// \instr~28_combout  = (\nRST~input_o  & ((ccifiwait_0 & (instr_9)) # (!ccifiwait_0 & ((ramiframload_9)))))

	.dataa(instr_9),
	.datab(nRST),
	.datac(ccifiwait_0),
	.datad(ramiframload_9),
	.cin(gnd),
	.combout(\instr~28_combout ),
	.cout());
// synopsys translate_off
defparam \instr~28 .lut_mask = 16'h8C80;
defparam \instr~28 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y31_N30
cycloneive_lcell_comb \instr[9]~feeder (
// Equation(s):
// \instr[9]~feeder_combout  = \instr~28_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(\instr~28_combout ),
	.cin(gnd),
	.combout(\instr[9]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \instr[9]~feeder .lut_mask = 16'hFF00;
defparam \instr[9]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y29_N2
cycloneive_lcell_comb \instr~29 (
// Equation(s):
// \instr~29_combout  = (\nRST~input_o  & ((ccifiwait_0 & ((instr_8))) # (!ccifiwait_0 & (ramiframload_8))))

	.dataa(ramiframload_8),
	.datab(instr_8),
	.datac(nRST),
	.datad(ccifiwait_0),
	.cin(gnd),
	.combout(\instr~29_combout ),
	.cout());
// synopsys translate_off
defparam \instr~29 .lut_mask = 16'hC0A0;
defparam \instr~29 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y29_N16
cycloneive_lcell_comb \instr[8]~feeder (
// Equation(s):
// \instr[8]~feeder_combout  = \instr~29_combout 

	.dataa(gnd),
	.datab(\instr~29_combout ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\instr[8]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \instr[8]~feeder .lut_mask = 16'hCCCC;
defparam \instr[8]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y30_N12
cycloneive_lcell_comb \instr~30 (
// Equation(s):
// \instr~30_combout  = (\nRST~input_o  & ((ccifiwait_0 & (instr_7)) # (!ccifiwait_0 & ((ramiframload_7)))))

	.dataa(nRST),
	.datab(instr_7),
	.datac(ramiframload_7),
	.datad(ccifiwait_0),
	.cin(gnd),
	.combout(\instr~30_combout ),
	.cout());
// synopsys translate_off
defparam \instr~30 .lut_mask = 16'h88A0;
defparam \instr~30 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y30_N4
cycloneive_lcell_comb \instr[7]~feeder (
// Equation(s):
// \instr[7]~feeder_combout  = \instr~30_combout 

	.dataa(\instr~30_combout ),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\instr[7]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \instr[7]~feeder .lut_mask = 16'hAAAA;
defparam \instr[7]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y30_N18
cycloneive_lcell_comb \instr~31 (
// Equation(s):
// \instr~31_combout  = (\nRST~input_o  & ((ccifiwait_0 & ((instr_6))) # (!ccifiwait_0 & (ramiframload_6))))

	.dataa(nRST),
	.datab(ramiframload_6),
	.datac(instr_6),
	.datad(ccifiwait_0),
	.cin(gnd),
	.combout(\instr~31_combout ),
	.cout());
// synopsys translate_off
defparam \instr~31 .lut_mask = 16'hA088;
defparam \instr~31 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y30_N22
cycloneive_lcell_comb \instr[6]~feeder (
// Equation(s):
// \instr[6]~feeder_combout  = \instr~31_combout 

	.dataa(gnd),
	.datab(\instr~31_combout ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\instr[6]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \instr[6]~feeder .lut_mask = 16'hCCCC;
defparam \instr[6]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

endmodule

module datapath (
	PCreg_1,
	PCreg_0,
	plif_exmemhlt_l,
	plif_exmemporto_l_1,
	plif_exmemdmemWEN_l,
	plif_exmemdmemREN_l,
	plif_exmemporto_l_0,
	plif_exmemporto_l_3,
	PCreg_3,
	plif_exmemporto_l_2,
	PCreg_2,
	plif_exmemporto_l_5,
	PCreg_5,
	plif_exmemporto_l_4,
	PCreg_4,
	plif_exmemporto_l_7,
	PCreg_7,
	plif_exmemporto_l_6,
	PCreg_6,
	plif_exmemporto_l_9,
	PCreg_9,
	plif_exmemporto_l_8,
	PCreg_8,
	plif_exmemporto_l_11,
	PCreg_11,
	plif_exmemporto_l_10,
	PCreg_10,
	plif_exmemporto_l_13,
	PCreg_13,
	plif_exmemporto_l_12,
	PCreg_12,
	plif_exmemporto_l_15,
	PCreg_15,
	plif_exmemporto_l_14,
	PCreg_14,
	plif_exmemporto_l_17,
	PCreg_17,
	plif_exmemporto_l_16,
	PCreg_16,
	plif_exmemporto_l_19,
	PCreg_19,
	plif_exmemporto_l_18,
	PCreg_18,
	plif_exmemporto_l_21,
	PCreg_21,
	plif_exmemporto_l_20,
	PCreg_20,
	plif_exmemporto_l_23,
	PCreg_23,
	plif_exmemporto_l_22,
	PCreg_22,
	plif_exmemporto_l_25,
	PCreg_25,
	plif_exmemporto_l_24,
	PCreg_24,
	plif_exmemporto_l_27,
	PCreg_27,
	plif_exmemporto_l_26,
	PCreg_26,
	plif_exmemporto_l_29,
	PCreg_29,
	plif_exmemporto_l_28,
	PCreg_28,
	plif_exmemporto_l_31,
	PCreg_31,
	plif_exmemporto_l_30,
	PCreg_30,
	dpifimemREN,
	always1,
	ramiframload_0,
	ramiframload_1,
	ramiframload_2,
	ramiframload_3,
	ramiframload_4,
	ramiframload_5,
	ramiframload_6,
	ramiframload_7,
	ramiframload_8,
	ramiframload_9,
	ramiframload_10,
	ramiframload_11,
	ramiframload_12,
	ramiframload_13,
	ramiframload_14,
	ramiframload_15,
	ramiframload_16,
	ramiframload_17,
	ramiframload_18,
	ramiframload_19,
	ramiframload_20,
	ramiframload_21,
	ramiframload_22,
	ramiframload_23,
	ramiframload_24,
	ramiframload_25,
	ramiframload_26,
	ramiframload_27,
	ramiframload_28,
	ramiframload_29,
	ramiframload_30,
	ramiframload_31,
	always0,
	plif_exmemrdat2_l_0,
	plif_exmemrdat2_l_1,
	plif_exmemrdat2_l_2,
	plif_exmemrdat2_l_3,
	plif_exmemrdat2_l_4,
	plif_exmemrdat2_l_5,
	plif_exmemrdat2_l_6,
	plif_exmemrdat2_l_7,
	plif_exmemrdat2_l_8,
	plif_exmemrdat2_l_9,
	plif_exmemrdat2_l_10,
	plif_exmemrdat2_l_11,
	plif_exmemrdat2_l_12,
	plif_exmemrdat2_l_13,
	plif_exmemrdat2_l_14,
	plif_exmemrdat2_l_15,
	plif_exmemrdat2_l_16,
	plif_exmemrdat2_l_17,
	plif_exmemrdat2_l_18,
	plif_exmemrdat2_l_19,
	plif_exmemrdat2_l_20,
	plif_exmemrdat2_l_21,
	plif_exmemrdat2_l_22,
	plif_exmemrdat2_l_23,
	plif_exmemrdat2_l_24,
	plif_exmemrdat2_l_25,
	plif_exmemrdat2_l_26,
	plif_exmemrdat2_l_27,
	plif_exmemrdat2_l_28,
	plif_exmemrdat2_l_29,
	plif_exmemrdat2_l_30,
	plif_exmemrdat2_l_31,
	instr_31,
	instr_29,
	instr_27,
	instr_26,
	instr_28,
	instr_30,
	instr_5,
	instr_1,
	instr_0,
	instr_2,
	instr_3,
	instr_4,
	instr_22,
	instr_21,
	instr_24,
	instr_23,
	instr_25,
	instr_17,
	instr_16,
	instr_19,
	instr_18,
	instr_20,
	instr_15,
	instr_14,
	instr_13,
	instr_12,
	instr_11,
	instr_10,
	instr_9,
	instr_8,
	instr_7,
	instr_6,
	ccifiwait_0,
	CLK,
	nRST,
	devpor,
	devclrn,
	devoe);
output 	PCreg_1;
output 	PCreg_0;
output 	plif_exmemhlt_l;
output 	plif_exmemporto_l_1;
output 	plif_exmemdmemWEN_l;
output 	plif_exmemdmemREN_l;
output 	plif_exmemporto_l_0;
output 	plif_exmemporto_l_3;
output 	PCreg_3;
output 	plif_exmemporto_l_2;
output 	PCreg_2;
output 	plif_exmemporto_l_5;
output 	PCreg_5;
output 	plif_exmemporto_l_4;
output 	PCreg_4;
output 	plif_exmemporto_l_7;
output 	PCreg_7;
output 	plif_exmemporto_l_6;
output 	PCreg_6;
output 	plif_exmemporto_l_9;
output 	PCreg_9;
output 	plif_exmemporto_l_8;
output 	PCreg_8;
output 	plif_exmemporto_l_11;
output 	PCreg_11;
output 	plif_exmemporto_l_10;
output 	PCreg_10;
output 	plif_exmemporto_l_13;
output 	PCreg_13;
output 	plif_exmemporto_l_12;
output 	PCreg_12;
output 	plif_exmemporto_l_15;
output 	PCreg_15;
output 	plif_exmemporto_l_14;
output 	PCreg_14;
output 	plif_exmemporto_l_17;
output 	PCreg_17;
output 	plif_exmemporto_l_16;
output 	PCreg_16;
output 	plif_exmemporto_l_19;
output 	PCreg_19;
output 	plif_exmemporto_l_18;
output 	PCreg_18;
output 	plif_exmemporto_l_21;
output 	PCreg_21;
output 	plif_exmemporto_l_20;
output 	PCreg_20;
output 	plif_exmemporto_l_23;
output 	PCreg_23;
output 	plif_exmemporto_l_22;
output 	PCreg_22;
output 	plif_exmemporto_l_25;
output 	PCreg_25;
output 	plif_exmemporto_l_24;
output 	PCreg_24;
output 	plif_exmemporto_l_27;
output 	PCreg_27;
output 	plif_exmemporto_l_26;
output 	PCreg_26;
output 	plif_exmemporto_l_29;
output 	PCreg_29;
output 	plif_exmemporto_l_28;
output 	PCreg_28;
output 	plif_exmemporto_l_31;
output 	PCreg_31;
output 	plif_exmemporto_l_30;
output 	PCreg_30;
output 	dpifimemREN;
input 	always1;
input 	ramiframload_0;
input 	ramiframload_1;
input 	ramiframload_2;
input 	ramiframload_3;
input 	ramiframload_4;
input 	ramiframload_5;
input 	ramiframload_6;
input 	ramiframload_7;
input 	ramiframload_8;
input 	ramiframload_9;
input 	ramiframload_10;
input 	ramiframload_11;
input 	ramiframload_12;
input 	ramiframload_13;
input 	ramiframload_14;
input 	ramiframload_15;
input 	ramiframload_16;
input 	ramiframload_17;
input 	ramiframload_18;
input 	ramiframload_19;
input 	ramiframload_20;
input 	ramiframload_21;
input 	ramiframload_22;
input 	ramiframload_23;
input 	ramiframload_24;
input 	ramiframload_25;
input 	ramiframload_26;
input 	ramiframload_27;
input 	ramiframload_28;
input 	ramiframload_29;
input 	ramiframload_30;
input 	ramiframload_31;
input 	always0;
output 	plif_exmemrdat2_l_0;
output 	plif_exmemrdat2_l_1;
output 	plif_exmemrdat2_l_2;
output 	plif_exmemrdat2_l_3;
output 	plif_exmemrdat2_l_4;
output 	plif_exmemrdat2_l_5;
output 	plif_exmemrdat2_l_6;
output 	plif_exmemrdat2_l_7;
output 	plif_exmemrdat2_l_8;
output 	plif_exmemrdat2_l_9;
output 	plif_exmemrdat2_l_10;
output 	plif_exmemrdat2_l_11;
output 	plif_exmemrdat2_l_12;
output 	plif_exmemrdat2_l_13;
output 	plif_exmemrdat2_l_14;
output 	plif_exmemrdat2_l_15;
output 	plif_exmemrdat2_l_16;
output 	plif_exmemrdat2_l_17;
output 	plif_exmemrdat2_l_18;
output 	plif_exmemrdat2_l_19;
output 	plif_exmemrdat2_l_20;
output 	plif_exmemrdat2_l_21;
output 	plif_exmemrdat2_l_22;
output 	plif_exmemrdat2_l_23;
output 	plif_exmemrdat2_l_24;
output 	plif_exmemrdat2_l_25;
output 	plif_exmemrdat2_l_26;
output 	plif_exmemrdat2_l_27;
output 	plif_exmemrdat2_l_28;
output 	plif_exmemrdat2_l_29;
output 	plif_exmemrdat2_l_30;
output 	plif_exmemrdat2_l_31;
input 	instr_31;
input 	instr_29;
input 	instr_27;
input 	instr_26;
input 	instr_28;
input 	instr_30;
input 	instr_5;
input 	instr_1;
input 	instr_0;
input 	instr_2;
input 	instr_3;
input 	instr_4;
input 	instr_22;
input 	instr_21;
input 	instr_24;
input 	instr_23;
input 	instr_25;
input 	instr_17;
input 	instr_16;
input 	instr_19;
input 	instr_18;
input 	instr_20;
input 	instr_15;
input 	instr_14;
input 	instr_13;
input 	instr_12;
input 	instr_11;
input 	instr_10;
input 	instr_9;
input 	instr_8;
input 	instr_7;
input 	instr_6;
input 	ccifiwait_0;
input 	CLK;
input 	nRST;

// Design Ports Information

input 	devpor;
input 	devclrn;
input 	devoe;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
assign unknown = 1'bx;

wire \PC|pcif.rtnaddr[2]~0_combout ;
wire \PC|pcif.rtnaddr[3]~2_combout ;
wire \PC|pcif.rtnaddr[4]~4_combout ;
wire \PC|pcif.rtnaddr[5]~6_combout ;
wire \PC|pcif.rtnaddr[6]~8_combout ;
wire \PC|pcif.rtnaddr[7]~10_combout ;
wire \PC|pcif.rtnaddr[8]~12_combout ;
wire \PC|pcif.rtnaddr[9]~14_combout ;
wire \PC|pcif.rtnaddr[10]~16_combout ;
wire \PC|pcif.rtnaddr[11]~18_combout ;
wire \PC|pcif.rtnaddr[12]~20_combout ;
wire \PC|pcif.rtnaddr[13]~22_combout ;
wire \PC|pcif.rtnaddr[14]~24_combout ;
wire \PC|pcif.rtnaddr[15]~26_combout ;
wire \PC|pcif.rtnaddr[16]~28_combout ;
wire \PC|pcif.rtnaddr[17]~30_combout ;
wire \PC|pcif.rtnaddr[18]~32_combout ;
wire \PC|pcif.rtnaddr[19]~34_combout ;
wire \PC|pcif.rtnaddr[20]~36_combout ;
wire \PC|pcif.rtnaddr[21]~38_combout ;
wire \PC|pcif.rtnaddr[22]~40_combout ;
wire \PC|pcif.rtnaddr[23]~42_combout ;
wire \PC|pcif.rtnaddr[24]~44_combout ;
wire \PC|pcif.rtnaddr[25]~46_combout ;
wire \PC|pcif.rtnaddr[26]~48_combout ;
wire \PC|pcif.rtnaddr[27]~50_combout ;
wire \PC|pcif.rtnaddr[28]~52_combout ;
wire \PC|pcif.rtnaddr[29]~54_combout ;
wire \PC|pcif.rtnaddr[30]~56_combout ;
wire \PC|pcif.rtnaddr[31]~58_combout ;
wire \IDEX|plif_idex.hlt_l~q ;
wire \HU|ifid_sRST~2_combout ;
wire \HU|exmem_en~0_combout ;
wire \IDEX|plif_idex.alusrc_l~q ;
wire \EXMEM|plif_exmem.regen_l~q ;
wire \FU|always0~2_combout ;
wire \FU|always0~3_combout ;
wire \portb~0_combout ;
wire \portb~1_combout ;
wire \wdat[31]~0_combout ;
wire \wdat[31]~1_combout ;
wire \FU|always0~4_combout ;
wire \RF|Decoder0~20_combout ;
wire \FU|WideOr0~combout ;
wire \FU|fwdc~2_combout ;
wire \MEMWB|plif_memwb.regen_l~q ;
wire \portb~2_combout ;
wire \portb~3_combout ;
wire \portb~4_combout ;
wire \wdat[30]~2_combout ;
wire \wdat[30]~3_combout ;
wire \portb~5_combout ;
wire \portb~6_combout ;
wire \wdat[29]~4_combout ;
wire \wdat[29]~5_combout ;
wire \portb~7_combout ;
wire \portb~8_combout ;
wire \wdat[28]~6_combout ;
wire \wdat[28]~7_combout ;
wire \portb~9_combout ;
wire \portb~10_combout ;
wire \wdat[27]~8_combout ;
wire \wdat[27]~9_combout ;
wire \portb~11_combout ;
wire \portb~12_combout ;
wire \wdat[26]~10_combout ;
wire \wdat[26]~11_combout ;
wire \portb~13_combout ;
wire \portb~14_combout ;
wire \wdat[25]~12_combout ;
wire \wdat[25]~13_combout ;
wire \portb~15_combout ;
wire \portb~16_combout ;
wire \wdat[24]~14_combout ;
wire \wdat[24]~15_combout ;
wire \portb~17_combout ;
wire \portb~18_combout ;
wire \wdat[23]~16_combout ;
wire \wdat[23]~17_combout ;
wire \portb~19_combout ;
wire \portb~20_combout ;
wire \wdat[22]~18_combout ;
wire \wdat[22]~19_combout ;
wire \portb~21_combout ;
wire \portb~22_combout ;
wire \wdat[21]~20_combout ;
wire \wdat[21]~21_combout ;
wire \portb~23_combout ;
wire \portb~24_combout ;
wire \wdat[20]~22_combout ;
wire \wdat[20]~23_combout ;
wire \portb~25_combout ;
wire \portb~26_combout ;
wire \wdat[19]~24_combout ;
wire \wdat[19]~25_combout ;
wire \portb~27_combout ;
wire \portb~28_combout ;
wire \wdat[18]~26_combout ;
wire \wdat[18]~27_combout ;
wire \portb~29_combout ;
wire \portb~30_combout ;
wire \wdat[17]~28_combout ;
wire \wdat[17]~29_combout ;
wire \portb~31_combout ;
wire \portb~32_combout ;
wire \wdat[16]~30_combout ;
wire \wdat[16]~31_combout ;
wire \portb~33_combout ;
wire \portb~34_combout ;
wire \wdat[15]~32_combout ;
wire \wdat[15]~33_combout ;
wire \portb~35_combout ;
wire \portb~36_combout ;
wire \wdat[14]~34_combout ;
wire \wdat[14]~35_combout ;
wire \portb~37_combout ;
wire \portb~38_combout ;
wire \wdat[13]~36_combout ;
wire \wdat[13]~37_combout ;
wire \portb~39_combout ;
wire \portb~40_combout ;
wire \wdat[12]~38_combout ;
wire \wdat[12]~39_combout ;
wire \portb~41_combout ;
wire \portb~42_combout ;
wire \wdat[11]~40_combout ;
wire \wdat[11]~41_combout ;
wire \portb~43_combout ;
wire \portb~44_combout ;
wire \wdat[10]~42_combout ;
wire \wdat[10]~43_combout ;
wire \portb~45_combout ;
wire \portb~46_combout ;
wire \wdat[9]~44_combout ;
wire \wdat[9]~45_combout ;
wire \portb~47_combout ;
wire \portb~48_combout ;
wire \wdat[8]~46_combout ;
wire \wdat[8]~47_combout ;
wire \portb~49_combout ;
wire \portb~50_combout ;
wire \wdat[7]~48_combout ;
wire \wdat[7]~49_combout ;
wire \portb~51_combout ;
wire \portb~52_combout ;
wire \wdat[6]~50_combout ;
wire \wdat[6]~51_combout ;
wire \portb~53_combout ;
wire \portb~54_combout ;
wire \wdat[5]~52_combout ;
wire \wdat[5]~53_combout ;
wire \portb~55_combout ;
wire \portb~56_combout ;
wire \wdat[2]~54_combout ;
wire \wdat[2]~55_combout ;
wire \FU|fwda~3_combout ;
wire \FU|always0~8_combout ;
wire \porta~54_combout ;
wire \porta~55_combout ;
wire \wdat[1]~56_combout ;
wire \wdat[1]~57_combout ;
wire \porta~56_combout ;
wire \porta~57_combout ;
wire \wdat[0]~58_combout ;
wire \wdat[0]~59_combout ;
wire \portb~57_combout ;
wire \portb~58_combout ;
wire \portb~59_combout ;
wire \portb~60_combout ;
wire \wdat[4]~60_combout ;
wire \wdat[4]~61_combout ;
wire \porta~58_combout ;
wire \porta~59_combout ;
wire \wdat[3]~62_combout ;
wire \wdat[3]~63_combout ;
wire \porta~60_combout ;
wire \porta~61_combout ;
wire \portb~61_combout ;
wire \portb~62_combout ;
wire \porta~62_combout ;
wire \porta~63_combout ;
wire \porta~64_combout ;
wire \porta~65_combout ;
wire \porta~66_combout ;
wire \portb~63_combout ;
wire \portb~64_combout ;
wire \porta~67_combout ;
wire \porta~68_combout ;
wire \porta~69_combout ;
wire \porta~70_combout ;
wire \porta~71_combout ;
wire \porta~72_combout ;
wire \porta~73_combout ;
wire \porta~74_combout ;
wire \portb~65_combout ;
wire \portb~66_combout ;
wire \porta~75_combout ;
wire \porta~76_combout ;
wire \porta~77_combout ;
wire \porta~78_combout ;
wire \porta~79_combout ;
wire \porta~80_combout ;
wire \porta~81_combout ;
wire \porta~82_combout ;
wire \porta~83_combout ;
wire \porta~84_combout ;
wire \porta~85_combout ;
wire \porta~86_combout ;
wire \porta~87_combout ;
wire \porta~88_combout ;
wire \porta~89_combout ;
wire \porta~90_combout ;
wire \porta~91_combout ;
wire \ALU|Selector30~8_combout ;
wire \MEMWB|plif_memwb.btype_l~q ;
wire \MEMWB|plif_memwb.zero_l~q ;
wire \pcsrc~0_combout ;
wire \IDEX|plif_idex.dmemREN_l~q ;
wire \CU|Equal16~0_combout ;
wire \CU|Equal22~0_combout ;
wire \CU|WideNor0~2_combout ;
wire \CU|Equal11~0_combout ;
wire \CU|Equal26~0_combout ;
wire \CU|Equal21~0_combout ;
wire \CU|WideOr14~0_combout ;
wire \CU|Equal13~1_combout ;
wire \IDEX|aluop_l~0_combout ;
wire \CU|WideNor1~0_combout ;
wire \CU|Selector22~6_combout ;
wire \CU|Selector4~0_combout ;
wire \CU|Selector4~1_combout ;
wire \CU|Selector5~1_combout ;
wire \CU|Selector2~0_combout ;
wire \CU|Selector3~0_combout ;
wire \CU|Selector1~0_combout ;
wire \CU|Equal6~0_combout ;
wire \CU|Selector11~0_combout ;
wire \CU|Selector21~0_combout ;
wire \CU|Selector9~0_combout ;
wire \CU|Selector9~1_combout ;
wire \CU|Selector10~0_combout ;
wire \CU|Selector7~0_combout ;
wire \CU|Selector8~0_combout ;
wire \CU|Selector6~0_combout ;
wire \HU|ifid_en~0_combout ;
wire \IDEX|plif_idex.dmemWEN_l~q ;
wire \ALU|Selector31~8_combout ;
wire \ALU|Selector28~10_combout ;
wire \HU|rambusy~0_combout ;
wire \ALU|Selector29~8_combout ;
wire \ALU|Selector26~8_combout ;
wire \ALU|Selector27~8_combout ;
wire \ALU|Selector24~9_combout ;
wire \ALU|Selector25~7_combout ;
wire \ALU|Selector22~8_combout ;
wire \ALU|Selector23~9_combout ;
wire \ALU|Selector20~9_combout ;
wire \ALU|Selector21~8_combout ;
wire \ALU|Selector18~9_combout ;
wire \ALU|Selector19~8_combout ;
wire \ALU|Selector16~10_combout ;
wire \ALU|Selector17~7_combout ;
wire \ALU|Selector14~8_combout ;
wire \ALU|Selector15~8_combout ;
wire \ALU|Selector12~10_combout ;
wire \ALU|Selector13~8_combout ;
wire \ALU|Selector10~8_combout ;
wire \ALU|Selector11~9_combout ;
wire \ALU|Selector8~10_combout ;
wire \ALU|Selector9~8_combout ;
wire \ALU|Selector6~8_combout ;
wire \ALU|Selector7~11_combout ;
wire \ALU|Selector4~10_combout ;
wire \ALU|Selector5~8_combout ;
wire \ALU|Selector2~11_combout ;
wire \ALU|Selector3~11_combout ;
wire \ALU|Selector0~34_combout ;
wire \ALU|Selector1~20_combout ;
wire \CU|Equal23~0_combout ;
wire \HU|idex_sRST~3_combout ;
wire \HU|idex_sRST~4_combout ;
wire \CU|pcsrc~0_combout ;
wire \rdat2~64_combout ;
wire \CU|Equal1~0_combout ;
wire \CU|Equal20~0_combout ;
wire \CU|WideNor1~1_combout ;
wire \CU|Equal19~0_combout ;
wire \CU|Equal1~1_combout ;
wire \CU|Equal18~0_combout ;
wire \CU|Selector22~7_combout ;
wire \CU|WideOr14~combout ;
wire \CU|WideOr15~combout ;
wire \CU|WideOr16~0_combout ;
wire \IDEX|plif_idex.regen_l~q ;
wire \RF|Mux32~9_combout ;
wire \RF|Mux32~19_combout ;
wire \extimm[30]~0_combout ;
wire \Equal0~0_combout ;
wire \RF|Mux33~9_combout ;
wire \RF|Mux33~19_combout ;
wire \RF|Mux34~9_combout ;
wire \RF|Mux34~19_combout ;
wire \RF|Mux35~9_combout ;
wire \RF|Mux35~19_combout ;
wire \RF|Mux36~9_combout ;
wire \RF|Mux36~19_combout ;
wire \RF|Mux37~9_combout ;
wire \RF|Mux37~19_combout ;
wire \RF|Mux38~9_combout ;
wire \RF|Mux38~19_combout ;
wire \RF|Mux39~9_combout ;
wire \RF|Mux39~19_combout ;
wire \RF|Mux40~9_combout ;
wire \RF|Mux40~19_combout ;
wire \RF|Mux41~9_combout ;
wire \RF|Mux41~19_combout ;
wire \RF|Mux42~9_combout ;
wire \RF|Mux42~19_combout ;
wire \CU|Selector14~0_combout ;
wire \RF|Mux43~9_combout ;
wire \RF|Mux43~19_combout ;
wire \CU|Selector15~0_combout ;
wire \RF|Mux44~9_combout ;
wire \RF|Mux44~19_combout ;
wire \CU|Selector16~0_combout ;
wire \RF|Mux45~9_combout ;
wire \RF|Mux45~19_combout ;
wire \CU|Selector17~0_combout ;
wire \RF|Mux46~9_combout ;
wire \RF|Mux46~19_combout ;
wire \CU|Selector18~0_combout ;
wire \RF|Mux47~9_combout ;
wire \RF|Mux47~19_combout ;
wire \RF|Mux48~9_combout ;
wire \RF|Mux48~19_combout ;
wire \RF|Mux49~9_combout ;
wire \RF|Mux49~19_combout ;
wire \RF|Mux50~9_combout ;
wire \RF|Mux50~19_combout ;
wire \RF|Mux51~9_combout ;
wire \RF|Mux51~19_combout ;
wire \RF|Mux52~9_combout ;
wire \RF|Mux52~19_combout ;
wire \RF|Mux53~9_combout ;
wire \RF|Mux53~19_combout ;
wire \RF|Mux54~9_combout ;
wire \RF|Mux54~19_combout ;
wire \RF|Mux55~9_combout ;
wire \RF|Mux55~19_combout ;
wire \RF|Mux56~9_combout ;
wire \RF|Mux56~19_combout ;
wire \RF|Mux57~9_combout ;
wire \RF|Mux57~19_combout ;
wire \RF|Mux58~9_combout ;
wire \RF|Mux58~19_combout ;
wire \RF|Mux29~9_combout ;
wire \RF|Mux29~19_combout ;
wire \RF|Mux30~9_combout ;
wire \RF|Mux30~19_combout ;
wire \RF|Mux63~9_combout ;
wire \RF|Mux63~19_combout ;
wire \RF|Mux62~9_combout ;
wire \RF|Mux62~19_combout ;
wire \RF|Mux27~9_combout ;
wire \RF|Mux27~19_combout ;
wire \RF|Mux28~9_combout ;
wire \RF|Mux28~19_combout ;
wire \RF|Mux61~9_combout ;
wire \RF|Mux61~19_combout ;
wire \RF|Mux23~9_combout ;
wire \RF|Mux23~19_combout ;
wire \RF|Mux24~9_combout ;
wire \RF|Mux24~19_combout ;
wire \RF|Mux25~9_combout ;
wire \RF|Mux25~19_combout ;
wire \RF|Mux26~9_combout ;
wire \RF|Mux26~19_combout ;
wire \RF|Mux60~9_combout ;
wire \RF|Mux60~19_combout ;
wire \RF|Mux15~9_combout ;
wire \RF|Mux15~19_combout ;
wire \RF|Mux16~9_combout ;
wire \RF|Mux16~19_combout ;
wire \RF|Mux17~9_combout ;
wire \RF|Mux17~19_combout ;
wire \RF|Mux18~9_combout ;
wire \RF|Mux18~19_combout ;
wire \RF|Mux19~9_combout ;
wire \RF|Mux19~19_combout ;
wire \RF|Mux20~9_combout ;
wire \RF|Mux20~19_combout ;
wire \RF|Mux21~9_combout ;
wire \RF|Mux21~19_combout ;
wire \RF|Mux22~9_combout ;
wire \RF|Mux22~19_combout ;
wire \RF|Mux59~9_combout ;
wire \RF|Mux59~19_combout ;
wire \RF|Mux0~9_combout ;
wire \RF|Mux0~19_combout ;
wire \RF|Mux2~9_combout ;
wire \RF|Mux2~19_combout ;
wire \RF|Mux1~9_combout ;
wire \RF|Mux1~19_combout ;
wire \RF|Mux3~9_combout ;
wire \RF|Mux3~19_combout ;
wire \RF|Mux4~9_combout ;
wire \RF|Mux4~19_combout ;
wire \RF|Mux5~9_combout ;
wire \RF|Mux5~19_combout ;
wire \RF|Mux6~9_combout ;
wire \RF|Mux6~19_combout ;
wire \RF|Mux7~9_combout ;
wire \RF|Mux7~19_combout ;
wire \RF|Mux8~9_combout ;
wire \RF|Mux8~19_combout ;
wire \RF|Mux9~9_combout ;
wire \RF|Mux9~19_combout ;
wire \RF|Mux10~9_combout ;
wire \RF|Mux10~19_combout ;
wire \RF|Mux11~9_combout ;
wire \RF|Mux11~19_combout ;
wire \RF|Mux12~9_combout ;
wire \RF|Mux12~19_combout ;
wire \RF|Mux13~9_combout ;
wire \RF|Mux13~19_combout ;
wire \RF|Mux14~9_combout ;
wire \RF|Mux14~19_combout ;
wire \RF|Mux31~9_combout ;
wire \RF|Mux31~19_combout ;
wire \EXMEM|plif_exmem.btype_l~q ;
wire \EXMEM|plif_exmem.zero_l~q ;
wire \CU|Selector24~0_combout ;
wire \rdat2~65_combout ;
wire \rdat2~66_combout ;
wire \rdat2~67_combout ;
wire \rdat2~68_combout ;
wire \rdat2~69_combout ;
wire \rdat2~70_combout ;
wire \rdat2~71_combout ;
wire \rdat2~72_combout ;
wire \rdat2~73_combout ;
wire \rdat2~74_combout ;
wire \rdat2~75_combout ;
wire \rdat2~76_combout ;
wire \rdat2~77_combout ;
wire \rdat2~78_combout ;
wire \rdat2~79_combout ;
wire \rdat2~80_combout ;
wire \rdat2~81_combout ;
wire \rdat2~82_combout ;
wire \rdat2~83_combout ;
wire \rdat2~84_combout ;
wire \rdat2~85_combout ;
wire \rdat2~86_combout ;
wire \rdat2~87_combout ;
wire \rdat2~88_combout ;
wire \rdat2~89_combout ;
wire \rdat2~90_combout ;
wire \rdat2~91_combout ;
wire \rdat2~92_combout ;
wire \rdat2~93_combout ;
wire \rdat2~94_combout ;
wire \rdat2~95_combout ;
wire \IDEX|plif_idex.btype_l~q ;
wire \ALU|WideOr1~combout ;
wire \CU|Equal12~0_combout ;
wire \porta~92_combout ;
wire \porta~93_combout ;
wire \porta~94_combout ;
wire \porta~95_combout ;
wire \porta~96_combout ;
wire \porta~97_combout ;
wire \porta~98_combout ;
wire \porta~99_combout ;
wire \porta~100_combout ;
wire \porta~101_combout ;
wire \porta~102_combout ;
wire \porta~103_combout ;
wire \porta~104_combout ;
wire \porta~105_combout ;
wire \porta~106_combout ;
wire \porta~107_combout ;
wire \porta~108_combout ;
wire \porta~109_combout ;
wire \porta~110_combout ;
wire \porta~111_combout ;
wire \porta~112_combout ;
wire \porta~113_combout ;
wire \porta~114_combout ;
wire \porta~115_combout ;
wire \porta~116_combout ;
wire \porta~117_combout ;
wire \porta~118_combout ;
wire \HU|idex_sRST~5_combout ;
wire \rdat2~96_combout ;
wire \CU|Selector0~2_combout ;
wire \HU|ifid_sRST~3_combout ;
wire \rdat2~97_combout ;
wire \rdat2~98_combout ;
wire \rdat2~99_combout ;
wire \rdat2~100_combout ;
wire \rdat2~101_combout ;
wire \rdat2~102_combout ;
wire \rdat2~103_combout ;
wire \rdat2~104_combout ;
wire \rdat2~105_combout ;
wire \rdat2~106_combout ;
wire \rdat2~107_combout ;
wire \rdat2~108_combout ;
wire \rdat2~109_combout ;
wire \rdat2~110_combout ;
wire \rdat2~111_combout ;
wire \rdat2~112_combout ;
wire \rdat2~113_combout ;
wire \rdat2~114_combout ;
wire \rdat2~115_combout ;
wire \rdat2~116_combout ;
wire \rdat2~117_combout ;
wire \rdat2~118_combout ;
wire \rdat2~119_combout ;
wire \rdat2~120_combout ;
wire \rdat2~121_combout ;
wire \rdat2~122_combout ;
wire \rdat2~123_combout ;
wire \rdat2~124_combout ;
wire \rdat2~125_combout ;
wire \rdat2~126_combout ;
wire \rdat2~127_combout ;
wire \CU|Equal25~4_combout ;
wire \dpif.imemREN~0_combout ;
wire [31:0] \IFID|plif_ifid.rtnaddr_l ;
wire [31:0] \IFID|plif_ifid.instr_l ;
wire [4:0] \IDEX|plif_idex.wsel_l ;
wire [31:0] \IDEX|plif_idex.rtnaddr_l ;
wire [4:0] \IDEX|plif_idex.rsel2_l ;
wire [4:0] \IDEX|plif_idex.rsel1_l ;
wire [1:0] \IDEX|plif_idex.regsrc_l ;
wire [31:0] \IDEX|plif_idex.rdat2_l ;
wire [31:0] \IDEX|plif_idex.rdat1_l ;
wire [1:0] \IDEX|plif_idex.pcsrc_l ;
wire [25:0] \IDEX|plif_idex.jaddr_l ;
wire [31:0] \IDEX|plif_idex.extimm_l ;
wire [3:0] \IDEX|plif_idex.aluop_l ;
wire [4:0] \EXMEM|plif_exmem.wsel_l ;
wire [31:0] \EXMEM|plif_exmem.rtnaddr_l ;
wire [1:0] \EXMEM|plif_exmem.regsrc_l ;
wire [1:0] \EXMEM|plif_exmem.pcsrc_l ;
wire [25:0] \EXMEM|plif_exmem.jaddr_l ;
wire [31:0] \EXMEM|plif_exmem.extimm_l ;
wire [4:0] \MEMWB|plif_memwb.wsel_l ;
wire [31:0] \MEMWB|plif_memwb.rtnaddr_l ;
wire [1:0] \MEMWB|plif_memwb.regsrc_l ;
wire [31:0] \MEMWB|plif_memwb.porto_l ;
wire [1:0] \MEMWB|plif_memwb.pcsrc_l ;
wire [25:0] \MEMWB|plif_memwb.jaddr_l ;
wire [31:0] \MEMWB|plif_memwb.extimm_l ;
wire [31:0] \MEMWB|plif_memwb.dmemload_l ;


pipeline_memwb MEMWB(
	.plif_exmemporto_l_1(plif_exmemporto_l_1),
	.plif_exmemporto_l_0(plif_exmemporto_l_0),
	.plif_exmemporto_l_3(plif_exmemporto_l_3),
	.plif_exmemporto_l_2(plif_exmemporto_l_2),
	.plif_exmemporto_l_5(plif_exmemporto_l_5),
	.plif_exmemporto_l_4(plif_exmemporto_l_4),
	.plif_exmemporto_l_7(plif_exmemporto_l_7),
	.plif_exmemporto_l_6(plif_exmemporto_l_6),
	.plif_exmemporto_l_9(plif_exmemporto_l_9),
	.plif_exmemporto_l_8(plif_exmemporto_l_8),
	.plif_exmemporto_l_11(plif_exmemporto_l_11),
	.plif_exmemporto_l_10(plif_exmemporto_l_10),
	.plif_exmemporto_l_13(plif_exmemporto_l_13),
	.plif_exmemporto_l_12(plif_exmemporto_l_12),
	.plif_exmemporto_l_15(plif_exmemporto_l_15),
	.plif_exmemporto_l_14(plif_exmemporto_l_14),
	.plif_exmemporto_l_17(plif_exmemporto_l_17),
	.plif_exmemporto_l_16(plif_exmemporto_l_16),
	.plif_exmemporto_l_19(plif_exmemporto_l_19),
	.plif_exmemporto_l_18(plif_exmemporto_l_18),
	.plif_exmemporto_l_21(plif_exmemporto_l_21),
	.plif_exmemporto_l_20(plif_exmemporto_l_20),
	.plif_exmemporto_l_23(plif_exmemporto_l_23),
	.plif_exmemporto_l_22(plif_exmemporto_l_22),
	.plif_exmemporto_l_25(plif_exmemporto_l_25),
	.plif_exmemporto_l_24(plif_exmemporto_l_24),
	.plif_exmemporto_l_27(plif_exmemporto_l_27),
	.plif_exmemporto_l_26(plif_exmemporto_l_26),
	.plif_exmemporto_l_29(plif_exmemporto_l_29),
	.plif_exmemporto_l_28(plif_exmemporto_l_28),
	.plif_exmemporto_l_31(plif_exmemporto_l_31),
	.plif_exmemporto_l_30(plif_exmemporto_l_30),
	.ramiframload_0(ramiframload_0),
	.ramiframload_1(ramiframload_1),
	.ramiframload_2(ramiframload_2),
	.ramiframload_3(ramiframload_3),
	.ramiframload_4(ramiframload_4),
	.ramiframload_5(ramiframload_5),
	.ramiframload_6(ramiframload_6),
	.ramiframload_7(ramiframload_7),
	.ramiframload_8(ramiframload_8),
	.ramiframload_9(ramiframload_9),
	.ramiframload_10(ramiframload_10),
	.ramiframload_11(ramiframload_11),
	.ramiframload_12(ramiframload_12),
	.ramiframload_13(ramiframload_13),
	.ramiframload_14(ramiframload_14),
	.ramiframload_15(ramiframload_15),
	.ramiframload_16(ramiframload_16),
	.ramiframload_17(ramiframload_17),
	.ramiframload_18(ramiframload_18),
	.ramiframload_19(ramiframload_19),
	.ramiframload_20(ramiframload_20),
	.ramiframload_21(ramiframload_21),
	.ramiframload_22(ramiframload_22),
	.ramiframload_23(ramiframload_23),
	.ramiframload_24(ramiframload_24),
	.ramiframload_25(ramiframload_25),
	.ramiframload_26(ramiframload_26),
	.ramiframload_27(ramiframload_27),
	.ramiframload_28(ramiframload_28),
	.ramiframload_29(ramiframload_29),
	.ramiframload_30(ramiframload_30),
	.ramiframload_31(ramiframload_31),
	.plif_memwbpcsrc_l_1(\MEMWB|plif_memwb.pcsrc_l [1]),
	.plif_memwbpcsrc_l_0(\MEMWB|plif_memwb.pcsrc_l [0]),
	.plif_exmempcsrc_l_1(\EXMEM|plif_exmem.pcsrc_l [1]),
	.plif_exmempcsrc_l_0(\EXMEM|plif_exmem.pcsrc_l [0]),
	.plif_exmemregen_l(\EXMEM|plif_exmem.regen_l~q ),
	.plif_exmemwsel_l_0(\EXMEM|plif_exmem.wsel_l [0]),
	.plif_exmemwsel_l_1(\EXMEM|plif_exmem.wsel_l [1]),
	.plif_exmemwsel_l_4(\EXMEM|plif_exmem.wsel_l [4]),
	.plif_exmemwsel_l_3(\EXMEM|plif_exmem.wsel_l [3]),
	.plif_exmemwsel_l_2(\EXMEM|plif_exmem.wsel_l [2]),
	.plif_memwbdmemload_l_31(\MEMWB|plif_memwb.dmemload_l [31]),
	.plif_memwbporto_l_31(\MEMWB|plif_memwb.porto_l [31]),
	.plif_memwbregsrc_l_0(\MEMWB|plif_memwb.regsrc_l [0]),
	.plif_memwbregsrc_l_1(\MEMWB|plif_memwb.regsrc_l [1]),
	.plif_memwbrtnaddr_l_31(\MEMWB|plif_memwb.rtnaddr_l [31]),
	.plif_memwbwsel_l_4(\MEMWB|plif_memwb.wsel_l [4]),
	.plif_memwbwsel_l_3(\MEMWB|plif_memwb.wsel_l [3]),
	.plif_memwbwsel_l_0(\MEMWB|plif_memwb.wsel_l [0]),
	.plif_memwbwsel_l_2(\MEMWB|plif_memwb.wsel_l [2]),
	.plif_memwbwsel_l_1(\MEMWB|plif_memwb.wsel_l [1]),
	.plif_memwbregen_l(\MEMWB|plif_memwb.regen_l~q ),
	.plif_memwbdmemload_l_30(\MEMWB|plif_memwb.dmemload_l [30]),
	.plif_memwbporto_l_30(\MEMWB|plif_memwb.porto_l [30]),
	.plif_memwbrtnaddr_l_30(\MEMWB|plif_memwb.rtnaddr_l [30]),
	.plif_memwbdmemload_l_29(\MEMWB|plif_memwb.dmemload_l [29]),
	.plif_memwbporto_l_29(\MEMWB|plif_memwb.porto_l [29]),
	.plif_memwbrtnaddr_l_29(\MEMWB|plif_memwb.rtnaddr_l [29]),
	.plif_memwbdmemload_l_28(\MEMWB|plif_memwb.dmemload_l [28]),
	.plif_memwbporto_l_28(\MEMWB|plif_memwb.porto_l [28]),
	.plif_memwbrtnaddr_l_28(\MEMWB|plif_memwb.rtnaddr_l [28]),
	.plif_memwbdmemload_l_27(\MEMWB|plif_memwb.dmemload_l [27]),
	.plif_memwbporto_l_27(\MEMWB|plif_memwb.porto_l [27]),
	.plif_memwbrtnaddr_l_27(\MEMWB|plif_memwb.rtnaddr_l [27]),
	.plif_memwbdmemload_l_26(\MEMWB|plif_memwb.dmemload_l [26]),
	.plif_memwbporto_l_26(\MEMWB|plif_memwb.porto_l [26]),
	.plif_memwbrtnaddr_l_26(\MEMWB|plif_memwb.rtnaddr_l [26]),
	.plif_memwbdmemload_l_25(\MEMWB|plif_memwb.dmemload_l [25]),
	.plif_memwbporto_l_25(\MEMWB|plif_memwb.porto_l [25]),
	.plif_memwbrtnaddr_l_25(\MEMWB|plif_memwb.rtnaddr_l [25]),
	.plif_memwbdmemload_l_24(\MEMWB|plif_memwb.dmemload_l [24]),
	.plif_memwbporto_l_24(\MEMWB|plif_memwb.porto_l [24]),
	.plif_memwbrtnaddr_l_24(\MEMWB|plif_memwb.rtnaddr_l [24]),
	.plif_memwbdmemload_l_23(\MEMWB|plif_memwb.dmemload_l [23]),
	.plif_memwbporto_l_23(\MEMWB|plif_memwb.porto_l [23]),
	.plif_memwbrtnaddr_l_23(\MEMWB|plif_memwb.rtnaddr_l [23]),
	.plif_memwbdmemload_l_22(\MEMWB|plif_memwb.dmemload_l [22]),
	.plif_memwbporto_l_22(\MEMWB|plif_memwb.porto_l [22]),
	.plif_memwbrtnaddr_l_22(\MEMWB|plif_memwb.rtnaddr_l [22]),
	.plif_memwbdmemload_l_21(\MEMWB|plif_memwb.dmemload_l [21]),
	.plif_memwbporto_l_21(\MEMWB|plif_memwb.porto_l [21]),
	.plif_memwbrtnaddr_l_21(\MEMWB|plif_memwb.rtnaddr_l [21]),
	.plif_memwbdmemload_l_20(\MEMWB|plif_memwb.dmemload_l [20]),
	.plif_memwbporto_l_20(\MEMWB|plif_memwb.porto_l [20]),
	.plif_memwbrtnaddr_l_20(\MEMWB|plif_memwb.rtnaddr_l [20]),
	.plif_memwbdmemload_l_19(\MEMWB|plif_memwb.dmemload_l [19]),
	.plif_memwbporto_l_19(\MEMWB|plif_memwb.porto_l [19]),
	.plif_memwbrtnaddr_l_19(\MEMWB|plif_memwb.rtnaddr_l [19]),
	.plif_memwbdmemload_l_18(\MEMWB|plif_memwb.dmemload_l [18]),
	.plif_memwbporto_l_18(\MEMWB|plif_memwb.porto_l [18]),
	.plif_memwbrtnaddr_l_18(\MEMWB|plif_memwb.rtnaddr_l [18]),
	.plif_memwbdmemload_l_17(\MEMWB|plif_memwb.dmemload_l [17]),
	.plif_memwbporto_l_17(\MEMWB|plif_memwb.porto_l [17]),
	.plif_memwbrtnaddr_l_17(\MEMWB|plif_memwb.rtnaddr_l [17]),
	.plif_memwbdmemload_l_16(\MEMWB|plif_memwb.dmemload_l [16]),
	.plif_memwbporto_l_16(\MEMWB|plif_memwb.porto_l [16]),
	.plif_memwbrtnaddr_l_16(\MEMWB|plif_memwb.rtnaddr_l [16]),
	.plif_memwbdmemload_l_15(\MEMWB|plif_memwb.dmemload_l [15]),
	.plif_memwbporto_l_15(\MEMWB|plif_memwb.porto_l [15]),
	.plif_memwbrtnaddr_l_15(\MEMWB|plif_memwb.rtnaddr_l [15]),
	.plif_memwbdmemload_l_14(\MEMWB|plif_memwb.dmemload_l [14]),
	.plif_memwbporto_l_14(\MEMWB|plif_memwb.porto_l [14]),
	.plif_memwbrtnaddr_l_14(\MEMWB|plif_memwb.rtnaddr_l [14]),
	.plif_memwbdmemload_l_13(\MEMWB|plif_memwb.dmemload_l [13]),
	.plif_memwbporto_l_13(\MEMWB|plif_memwb.porto_l [13]),
	.plif_memwbrtnaddr_l_13(\MEMWB|plif_memwb.rtnaddr_l [13]),
	.plif_memwbdmemload_l_12(\MEMWB|plif_memwb.dmemload_l [12]),
	.plif_memwbporto_l_12(\MEMWB|plif_memwb.porto_l [12]),
	.plif_memwbrtnaddr_l_12(\MEMWB|plif_memwb.rtnaddr_l [12]),
	.plif_memwbdmemload_l_11(\MEMWB|plif_memwb.dmemload_l [11]),
	.plif_memwbporto_l_11(\MEMWB|plif_memwb.porto_l [11]),
	.plif_memwbrtnaddr_l_11(\MEMWB|plif_memwb.rtnaddr_l [11]),
	.plif_memwbdmemload_l_10(\MEMWB|plif_memwb.dmemload_l [10]),
	.plif_memwbporto_l_10(\MEMWB|plif_memwb.porto_l [10]),
	.plif_memwbrtnaddr_l_10(\MEMWB|plif_memwb.rtnaddr_l [10]),
	.plif_memwbdmemload_l_9(\MEMWB|plif_memwb.dmemload_l [9]),
	.plif_memwbporto_l_9(\MEMWB|plif_memwb.porto_l [9]),
	.plif_memwbrtnaddr_l_9(\MEMWB|plif_memwb.rtnaddr_l [9]),
	.plif_memwbdmemload_l_8(\MEMWB|plif_memwb.dmemload_l [8]),
	.plif_memwbporto_l_8(\MEMWB|plif_memwb.porto_l [8]),
	.plif_memwbrtnaddr_l_8(\MEMWB|plif_memwb.rtnaddr_l [8]),
	.plif_memwbdmemload_l_7(\MEMWB|plif_memwb.dmemload_l [7]),
	.plif_memwbporto_l_7(\MEMWB|plif_memwb.porto_l [7]),
	.plif_memwbrtnaddr_l_7(\MEMWB|plif_memwb.rtnaddr_l [7]),
	.plif_memwbdmemload_l_6(\MEMWB|plif_memwb.dmemload_l [6]),
	.plif_memwbporto_l_6(\MEMWB|plif_memwb.porto_l [6]),
	.plif_memwbrtnaddr_l_6(\MEMWB|plif_memwb.rtnaddr_l [6]),
	.plif_memwbdmemload_l_5(\MEMWB|plif_memwb.dmemload_l [5]),
	.plif_memwbporto_l_5(\MEMWB|plif_memwb.porto_l [5]),
	.plif_memwbrtnaddr_l_5(\MEMWB|plif_memwb.rtnaddr_l [5]),
	.plif_memwbdmemload_l_2(\MEMWB|plif_memwb.dmemload_l [2]),
	.plif_memwbporto_l_2(\MEMWB|plif_memwb.porto_l [2]),
	.plif_memwbrtnaddr_l_2(\MEMWB|plif_memwb.rtnaddr_l [2]),
	.plif_memwbdmemload_l_1(\MEMWB|plif_memwb.dmemload_l [1]),
	.plif_memwbporto_l_1(\MEMWB|plif_memwb.porto_l [1]),
	.plif_memwbrtnaddr_l_1(\MEMWB|plif_memwb.rtnaddr_l [1]),
	.plif_memwbdmemload_l_0(\MEMWB|plif_memwb.dmemload_l [0]),
	.plif_memwbporto_l_0(\MEMWB|plif_memwb.porto_l [0]),
	.plif_memwbrtnaddr_l_0(\MEMWB|plif_memwb.rtnaddr_l [0]),
	.plif_memwbdmemload_l_4(\MEMWB|plif_memwb.dmemload_l [4]),
	.plif_memwbporto_l_4(\MEMWB|plif_memwb.porto_l [4]),
	.plif_memwbrtnaddr_l_4(\MEMWB|plif_memwb.rtnaddr_l [4]),
	.plif_memwbdmemload_l_3(\MEMWB|plif_memwb.dmemload_l [3]),
	.plif_memwbporto_l_3(\MEMWB|plif_memwb.porto_l [3]),
	.plif_memwbrtnaddr_l_3(\MEMWB|plif_memwb.rtnaddr_l [3]),
	.plif_memwbbtype_l(\MEMWB|plif_memwb.btype_l~q ),
	.plif_memwbzero_l(\MEMWB|plif_memwb.zero_l~q ),
	.plif_memwbjaddr_l_1(\MEMWB|plif_memwb.jaddr_l [1]),
	.plif_memwbextimm_l_1(\MEMWB|plif_memwb.extimm_l [1]),
	.plif_memwbextimm_l_0(\MEMWB|plif_memwb.extimm_l [0]),
	.plif_memwbjaddr_l_0(\MEMWB|plif_memwb.jaddr_l [0]),
	.plif_memwbjaddr_l_3(\MEMWB|plif_memwb.jaddr_l [3]),
	.plif_memwbextimm_l_3(\MEMWB|plif_memwb.extimm_l [3]),
	.plif_memwbextimm_l_2(\MEMWB|plif_memwb.extimm_l [2]),
	.plif_memwbjaddr_l_2(\MEMWB|plif_memwb.jaddr_l [2]),
	.plif_memwbjaddr_l_5(\MEMWB|plif_memwb.jaddr_l [5]),
	.plif_memwbextimm_l_5(\MEMWB|plif_memwb.extimm_l [5]),
	.plif_memwbextimm_l_4(\MEMWB|plif_memwb.extimm_l [4]),
	.plif_memwbjaddr_l_4(\MEMWB|plif_memwb.jaddr_l [4]),
	.plif_memwbjaddr_l_7(\MEMWB|plif_memwb.jaddr_l [7]),
	.plif_memwbextimm_l_7(\MEMWB|plif_memwb.extimm_l [7]),
	.plif_memwbextimm_l_6(\MEMWB|plif_memwb.extimm_l [6]),
	.plif_memwbjaddr_l_6(\MEMWB|plif_memwb.jaddr_l [6]),
	.plif_memwbjaddr_l_9(\MEMWB|plif_memwb.jaddr_l [9]),
	.plif_memwbextimm_l_9(\MEMWB|plif_memwb.extimm_l [9]),
	.plif_memwbextimm_l_8(\MEMWB|plif_memwb.extimm_l [8]),
	.plif_memwbjaddr_l_8(\MEMWB|plif_memwb.jaddr_l [8]),
	.plif_memwbjaddr_l_11(\MEMWB|plif_memwb.jaddr_l [11]),
	.plif_memwbextimm_l_11(\MEMWB|plif_memwb.extimm_l [11]),
	.plif_memwbextimm_l_10(\MEMWB|plif_memwb.extimm_l [10]),
	.plif_memwbjaddr_l_10(\MEMWB|plif_memwb.jaddr_l [10]),
	.plif_memwbjaddr_l_13(\MEMWB|plif_memwb.jaddr_l [13]),
	.plif_memwbextimm_l_13(\MEMWB|plif_memwb.extimm_l [13]),
	.plif_memwbextimm_l_12(\MEMWB|plif_memwb.extimm_l [12]),
	.plif_memwbjaddr_l_12(\MEMWB|plif_memwb.jaddr_l [12]),
	.plif_memwbjaddr_l_15(\MEMWB|plif_memwb.jaddr_l [15]),
	.plif_memwbextimm_l_15(\MEMWB|plif_memwb.extimm_l [15]),
	.plif_memwbextimm_l_14(\MEMWB|plif_memwb.extimm_l [14]),
	.plif_memwbjaddr_l_14(\MEMWB|plif_memwb.jaddr_l [14]),
	.plif_memwbjaddr_l_17(\MEMWB|plif_memwb.jaddr_l [17]),
	.plif_memwbextimm_l_17(\MEMWB|plif_memwb.extimm_l [17]),
	.plif_memwbextimm_l_16(\MEMWB|plif_memwb.extimm_l [16]),
	.plif_memwbjaddr_l_16(\MEMWB|plif_memwb.jaddr_l [16]),
	.plif_memwbjaddr_l_19(\MEMWB|plif_memwb.jaddr_l [19]),
	.plif_memwbextimm_l_19(\MEMWB|plif_memwb.extimm_l [19]),
	.plif_memwbextimm_l_18(\MEMWB|plif_memwb.extimm_l [18]),
	.plif_memwbjaddr_l_18(\MEMWB|plif_memwb.jaddr_l [18]),
	.plif_memwbjaddr_l_21(\MEMWB|plif_memwb.jaddr_l [21]),
	.plif_memwbextimm_l_21(\MEMWB|plif_memwb.extimm_l [21]),
	.plif_memwbextimm_l_20(\MEMWB|plif_memwb.extimm_l [20]),
	.plif_memwbjaddr_l_20(\MEMWB|plif_memwb.jaddr_l [20]),
	.plif_memwbjaddr_l_23(\MEMWB|plif_memwb.jaddr_l [23]),
	.plif_memwbextimm_l_23(\MEMWB|plif_memwb.extimm_l [23]),
	.plif_memwbextimm_l_22(\MEMWB|plif_memwb.extimm_l [22]),
	.plif_memwbjaddr_l_22(\MEMWB|plif_memwb.jaddr_l [22]),
	.plif_memwbjaddr_l_25(\MEMWB|plif_memwb.jaddr_l [25]),
	.plif_memwbextimm_l_25(\MEMWB|plif_memwb.extimm_l [25]),
	.plif_memwbextimm_l_24(\MEMWB|plif_memwb.extimm_l [24]),
	.plif_memwbjaddr_l_24(\MEMWB|plif_memwb.jaddr_l [24]),
	.plif_memwbextimm_l_27(\MEMWB|plif_memwb.extimm_l [27]),
	.plif_memwbextimm_l_26(\MEMWB|plif_memwb.extimm_l [26]),
	.plif_memwbextimm_l_29(\MEMWB|plif_memwb.extimm_l [29]),
	.plif_memwbextimm_l_28(\MEMWB|plif_memwb.extimm_l [28]),
	.plif_exmemregsrc_l_0(\EXMEM|plif_exmem.regsrc_l [0]),
	.plif_exmemregsrc_l_1(\EXMEM|plif_exmem.regsrc_l [1]),
	.plif_exmemrtnaddr_l_31(\EXMEM|plif_exmem.rtnaddr_l [31]),
	.plif_exmemrtnaddr_l_30(\EXMEM|plif_exmem.rtnaddr_l [30]),
	.plif_exmemrtnaddr_l_29(\EXMEM|plif_exmem.rtnaddr_l [29]),
	.plif_exmemrtnaddr_l_28(\EXMEM|plif_exmem.rtnaddr_l [28]),
	.plif_exmemrtnaddr_l_27(\EXMEM|plif_exmem.rtnaddr_l [27]),
	.plif_exmemrtnaddr_l_26(\EXMEM|plif_exmem.rtnaddr_l [26]),
	.plif_exmemrtnaddr_l_25(\EXMEM|plif_exmem.rtnaddr_l [25]),
	.plif_exmemrtnaddr_l_24(\EXMEM|plif_exmem.rtnaddr_l [24]),
	.plif_exmemrtnaddr_l_23(\EXMEM|plif_exmem.rtnaddr_l [23]),
	.plif_exmemrtnaddr_l_22(\EXMEM|plif_exmem.rtnaddr_l [22]),
	.plif_exmemrtnaddr_l_21(\EXMEM|plif_exmem.rtnaddr_l [21]),
	.plif_exmemrtnaddr_l_20(\EXMEM|plif_exmem.rtnaddr_l [20]),
	.plif_exmemrtnaddr_l_19(\EXMEM|plif_exmem.rtnaddr_l [19]),
	.plif_exmemrtnaddr_l_18(\EXMEM|plif_exmem.rtnaddr_l [18]),
	.plif_exmemrtnaddr_l_17(\EXMEM|plif_exmem.rtnaddr_l [17]),
	.plif_exmemrtnaddr_l_16(\EXMEM|plif_exmem.rtnaddr_l [16]),
	.plif_exmemrtnaddr_l_15(\EXMEM|plif_exmem.rtnaddr_l [15]),
	.plif_exmemrtnaddr_l_14(\EXMEM|plif_exmem.rtnaddr_l [14]),
	.plif_exmemrtnaddr_l_13(\EXMEM|plif_exmem.rtnaddr_l [13]),
	.plif_exmemrtnaddr_l_12(\EXMEM|plif_exmem.rtnaddr_l [12]),
	.plif_exmemrtnaddr_l_11(\EXMEM|plif_exmem.rtnaddr_l [11]),
	.plif_exmemrtnaddr_l_10(\EXMEM|plif_exmem.rtnaddr_l [10]),
	.plif_exmemrtnaddr_l_9(\EXMEM|plif_exmem.rtnaddr_l [9]),
	.plif_exmemrtnaddr_l_8(\EXMEM|plif_exmem.rtnaddr_l [8]),
	.plif_exmemrtnaddr_l_7(\EXMEM|plif_exmem.rtnaddr_l [7]),
	.plif_exmemrtnaddr_l_6(\EXMEM|plif_exmem.rtnaddr_l [6]),
	.plif_exmemrtnaddr_l_5(\EXMEM|plif_exmem.rtnaddr_l [5]),
	.plif_exmemrtnaddr_l_2(\EXMEM|plif_exmem.rtnaddr_l [2]),
	.plif_exmemrtnaddr_l_1(\EXMEM|plif_exmem.rtnaddr_l [1]),
	.plif_exmemrtnaddr_l_0(\EXMEM|plif_exmem.rtnaddr_l [0]),
	.plif_exmemrtnaddr_l_4(\EXMEM|plif_exmem.rtnaddr_l [4]),
	.plif_exmemrtnaddr_l_3(\EXMEM|plif_exmem.rtnaddr_l [3]),
	.plif_exmembtype_l(\EXMEM|plif_exmem.btype_l~q ),
	.plif_exmemzero_l(\EXMEM|plif_exmem.zero_l~q ),
	.plif_exmemjaddr_l_1(\EXMEM|plif_exmem.jaddr_l [1]),
	.plif_exmemextimm_l_1(\EXMEM|plif_exmem.extimm_l [1]),
	.plif_exmemextimm_l_0(\EXMEM|plif_exmem.extimm_l [0]),
	.plif_exmemjaddr_l_0(\EXMEM|plif_exmem.jaddr_l [0]),
	.plif_exmemjaddr_l_3(\EXMEM|plif_exmem.jaddr_l [3]),
	.plif_exmemextimm_l_3(\EXMEM|plif_exmem.extimm_l [3]),
	.plif_exmemextimm_l_2(\EXMEM|plif_exmem.extimm_l [2]),
	.plif_exmemjaddr_l_2(\EXMEM|plif_exmem.jaddr_l [2]),
	.plif_exmemjaddr_l_5(\EXMEM|plif_exmem.jaddr_l [5]),
	.plif_exmemextimm_l_5(\EXMEM|plif_exmem.extimm_l [5]),
	.plif_exmemextimm_l_4(\EXMEM|plif_exmem.extimm_l [4]),
	.plif_exmemjaddr_l_4(\EXMEM|plif_exmem.jaddr_l [4]),
	.plif_exmemjaddr_l_7(\EXMEM|plif_exmem.jaddr_l [7]),
	.plif_exmemextimm_l_7(\EXMEM|plif_exmem.extimm_l [7]),
	.plif_exmemextimm_l_6(\EXMEM|plif_exmem.extimm_l [6]),
	.plif_exmemjaddr_l_6(\EXMEM|plif_exmem.jaddr_l [6]),
	.plif_exmemjaddr_l_9(\EXMEM|plif_exmem.jaddr_l [9]),
	.plif_exmemextimm_l_9(\EXMEM|plif_exmem.extimm_l [9]),
	.plif_exmemextimm_l_8(\EXMEM|plif_exmem.extimm_l [8]),
	.plif_exmemjaddr_l_8(\EXMEM|plif_exmem.jaddr_l [8]),
	.plif_exmemjaddr_l_11(\EXMEM|plif_exmem.jaddr_l [11]),
	.plif_exmemextimm_l_11(\EXMEM|plif_exmem.extimm_l [11]),
	.plif_exmemextimm_l_10(\EXMEM|plif_exmem.extimm_l [10]),
	.plif_exmemjaddr_l_10(\EXMEM|plif_exmem.jaddr_l [10]),
	.plif_exmemjaddr_l_13(\EXMEM|plif_exmem.jaddr_l [13]),
	.plif_exmemextimm_l_13(\EXMEM|plif_exmem.extimm_l [13]),
	.plif_exmemextimm_l_12(\EXMEM|plif_exmem.extimm_l [12]),
	.plif_exmemjaddr_l_12(\EXMEM|plif_exmem.jaddr_l [12]),
	.plif_exmemjaddr_l_15(\EXMEM|plif_exmem.jaddr_l [15]),
	.plif_exmemextimm_l_15(\EXMEM|plif_exmem.extimm_l [15]),
	.plif_exmemextimm_l_14(\EXMEM|plif_exmem.extimm_l [14]),
	.plif_exmemjaddr_l_14(\EXMEM|plif_exmem.jaddr_l [14]),
	.plif_exmemjaddr_l_17(\EXMEM|plif_exmem.jaddr_l [17]),
	.plif_exmemextimm_l_17(\EXMEM|plif_exmem.extimm_l [17]),
	.plif_exmemextimm_l_16(\EXMEM|plif_exmem.extimm_l [16]),
	.plif_exmemjaddr_l_16(\EXMEM|plif_exmem.jaddr_l [16]),
	.plif_exmemjaddr_l_19(\EXMEM|plif_exmem.jaddr_l [19]),
	.plif_exmemextimm_l_19(\EXMEM|plif_exmem.extimm_l [19]),
	.plif_exmemextimm_l_18(\EXMEM|plif_exmem.extimm_l [18]),
	.plif_exmemjaddr_l_18(\EXMEM|plif_exmem.jaddr_l [18]),
	.plif_exmemjaddr_l_21(\EXMEM|plif_exmem.jaddr_l [21]),
	.plif_exmemextimm_l_21(\EXMEM|plif_exmem.extimm_l [21]),
	.plif_exmemextimm_l_20(\EXMEM|plif_exmem.extimm_l [20]),
	.plif_exmemjaddr_l_20(\EXMEM|plif_exmem.jaddr_l [20]),
	.plif_exmemjaddr_l_23(\EXMEM|plif_exmem.jaddr_l [23]),
	.plif_exmemextimm_l_23(\EXMEM|plif_exmem.extimm_l [23]),
	.plif_exmemextimm_l_22(\EXMEM|plif_exmem.extimm_l [22]),
	.plif_exmemjaddr_l_22(\EXMEM|plif_exmem.jaddr_l [22]),
	.plif_exmemjaddr_l_25(\EXMEM|plif_exmem.jaddr_l [25]),
	.plif_exmemextimm_l_25(\EXMEM|plif_exmem.extimm_l [25]),
	.plif_exmemextimm_l_24(\EXMEM|plif_exmem.extimm_l [24]),
	.plif_exmemjaddr_l_24(\EXMEM|plif_exmem.jaddr_l [24]),
	.plif_exmemextimm_l_27(\EXMEM|plif_exmem.extimm_l [27]),
	.plif_exmemextimm_l_26(\EXMEM|plif_exmem.extimm_l [26]),
	.plif_exmemextimm_l_29(\EXMEM|plif_exmem.extimm_l [29]),
	.plif_exmemextimm_l_28(\EXMEM|plif_exmem.extimm_l [28]),
	.CPUCLK(CLK),
	.nRST(nRST),
	.devpor(devpor),
	.devclrn(devclrn),
	.devoe(devoe));

pipeline_exmem EXMEM(
	.plif_exmemhlt_l(plif_exmemhlt_l),
	.plif_exmemporto_l_1(plif_exmemporto_l_1),
	.plif_exmemdmemWEN_l(plif_exmemdmemWEN_l),
	.plif_exmemdmemREN_l(plif_exmemdmemREN_l),
	.plif_exmemporto_l_0(plif_exmemporto_l_0),
	.plif_exmemporto_l_3(plif_exmemporto_l_3),
	.plif_exmemporto_l_2(plif_exmemporto_l_2),
	.plif_exmemporto_l_5(plif_exmemporto_l_5),
	.plif_exmemporto_l_4(plif_exmemporto_l_4),
	.plif_exmemporto_l_7(plif_exmemporto_l_7),
	.plif_exmemporto_l_6(plif_exmemporto_l_6),
	.plif_exmemporto_l_9(plif_exmemporto_l_9),
	.plif_exmemporto_l_8(plif_exmemporto_l_8),
	.plif_exmemporto_l_11(plif_exmemporto_l_11),
	.plif_exmemporto_l_10(plif_exmemporto_l_10),
	.plif_exmemporto_l_13(plif_exmemporto_l_13),
	.plif_exmemporto_l_12(plif_exmemporto_l_12),
	.plif_exmemporto_l_15(plif_exmemporto_l_15),
	.plif_exmemporto_l_14(plif_exmemporto_l_14),
	.plif_exmemporto_l_17(plif_exmemporto_l_17),
	.plif_exmemporto_l_16(plif_exmemporto_l_16),
	.plif_exmemporto_l_19(plif_exmemporto_l_19),
	.plif_exmemporto_l_18(plif_exmemporto_l_18),
	.plif_exmemporto_l_21(plif_exmemporto_l_21),
	.plif_exmemporto_l_20(plif_exmemporto_l_20),
	.plif_exmemporto_l_23(plif_exmemporto_l_23),
	.plif_exmemporto_l_22(plif_exmemporto_l_22),
	.plif_exmemporto_l_25(plif_exmemporto_l_25),
	.plif_exmemporto_l_24(plif_exmemporto_l_24),
	.plif_exmemporto_l_27(plif_exmemporto_l_27),
	.plif_exmemporto_l_26(plif_exmemporto_l_26),
	.plif_exmemporto_l_29(plif_exmemporto_l_29),
	.plif_exmemporto_l_28(plif_exmemporto_l_28),
	.plif_exmemporto_l_31(plif_exmemporto_l_31),
	.plif_exmemporto_l_30(plif_exmemporto_l_30),
	.plif_idexhlt_l(\IDEX|plif_idex.hlt_l~q ),
	.plif_idexpcsrc_l_1(\IDEX|plif_idex.pcsrc_l [1]),
	.plif_idexpcsrc_l_0(\IDEX|plif_idex.pcsrc_l [0]),
	.plif_exmempcsrc_l_1(\EXMEM|plif_exmem.pcsrc_l [1]),
	.plif_exmempcsrc_l_0(\EXMEM|plif_exmem.pcsrc_l [0]),
	.exmem_en(\HU|exmem_en~0_combout ),
	.plif_exmemrdat2_l_0(plif_exmemrdat2_l_0),
	.plif_exmemregen_l(\EXMEM|plif_exmem.regen_l~q ),
	.plif_exmemwsel_l_0(\EXMEM|plif_exmem.wsel_l [0]),
	.plif_exmemwsel_l_1(\EXMEM|plif_exmem.wsel_l [1]),
	.plif_exmemwsel_l_4(\EXMEM|plif_exmem.wsel_l [4]),
	.plif_exmemwsel_l_3(\EXMEM|plif_exmem.wsel_l [3]),
	.plif_exmemwsel_l_2(\EXMEM|plif_exmem.wsel_l [2]),
	.plif_idexextimm_l_29(\IDEX|plif_idex.extimm_l [29]),
	.plif_idexextimm_l_28(\IDEX|plif_idex.extimm_l [28]),
	.plif_idexextimm_l_27(\IDEX|plif_idex.extimm_l [27]),
	.plif_idexextimm_l_26(\IDEX|plif_idex.extimm_l [26]),
	.plif_idexextimm_l_25(\IDEX|plif_idex.extimm_l [25]),
	.plif_idexextimm_l_24(\IDEX|plif_idex.extimm_l [24]),
	.plif_idexextimm_l_23(\IDEX|plif_idex.extimm_l [23]),
	.plif_idexextimm_l_22(\IDEX|plif_idex.extimm_l [22]),
	.plif_idexextimm_l_21(\IDEX|plif_idex.extimm_l [21]),
	.plif_idexextimm_l_20(\IDEX|plif_idex.extimm_l [20]),
	.plif_idexextimm_l_19(\IDEX|plif_idex.extimm_l [19]),
	.plif_idexextimm_l_18(\IDEX|plif_idex.extimm_l [18]),
	.plif_idexextimm_l_17(\IDEX|plif_idex.extimm_l [17]),
	.plif_idexextimm_l_16(\IDEX|plif_idex.extimm_l [16]),
	.plif_idexextimm_l_15(\IDEX|plif_idex.extimm_l [15]),
	.plif_idexextimm_l_14(\IDEX|plif_idex.extimm_l [14]),
	.plif_idexextimm_l_13(\IDEX|plif_idex.extimm_l [13]),
	.plif_idexextimm_l_12(\IDEX|plif_idex.extimm_l [12]),
	.plif_idexextimm_l_11(\IDEX|plif_idex.extimm_l [11]),
	.plif_idexextimm_l_10(\IDEX|plif_idex.extimm_l [10]),
	.plif_idexextimm_l_9(\IDEX|plif_idex.extimm_l [9]),
	.plif_idexextimm_l_8(\IDEX|plif_idex.extimm_l [8]),
	.plif_idexextimm_l_7(\IDEX|plif_idex.extimm_l [7]),
	.plif_idexextimm_l_6(\IDEX|plif_idex.extimm_l [6]),
	.plif_idexextimm_l_5(\IDEX|plif_idex.extimm_l [5]),
	.plif_idexextimm_l_0(\IDEX|plif_idex.extimm_l [0]),
	.plif_idexextimm_l_1(\IDEX|plif_idex.extimm_l [1]),
	.plif_idexextimm_l_2(\IDEX|plif_idex.extimm_l [2]),
	.plif_idexextimm_l_3(\IDEX|plif_idex.extimm_l [3]),
	.plif_idexextimm_l_4(\IDEX|plif_idex.extimm_l [4]),
	.Selector30(\ALU|Selector30~8_combout ),
	.plif_idexdmemREN_l(\IDEX|plif_idex.dmemREN_l~q ),
	.plif_idexwsel_l_0(\IDEX|plif_idex.wsel_l [0]),
	.plif_idexwsel_l_1(\IDEX|plif_idex.wsel_l [1]),
	.plif_idexwsel_l_2(\IDEX|plif_idex.wsel_l [2]),
	.plif_idexwsel_l_3(\IDEX|plif_idex.wsel_l [3]),
	.plif_idexwsel_l_4(\IDEX|plif_idex.wsel_l [4]),
	.plif_idexdmemWEN_l(\IDEX|plif_idex.dmemWEN_l~q ),
	.Selector31(\ALU|Selector31~8_combout ),
	.Selector28(\ALU|Selector28~10_combout ),
	.Selector29(\ALU|Selector29~8_combout ),
	.Selector26(\ALU|Selector26~8_combout ),
	.Selector27(\ALU|Selector27~8_combout ),
	.Selector24(\ALU|Selector24~9_combout ),
	.Selector25(\ALU|Selector25~7_combout ),
	.Selector22(\ALU|Selector22~8_combout ),
	.Selector23(\ALU|Selector23~9_combout ),
	.Selector20(\ALU|Selector20~9_combout ),
	.Selector21(\ALU|Selector21~8_combout ),
	.Selector18(\ALU|Selector18~9_combout ),
	.Selector19(\ALU|Selector19~8_combout ),
	.Selector16(\ALU|Selector16~10_combout ),
	.Selector17(\ALU|Selector17~7_combout ),
	.Selector14(\ALU|Selector14~8_combout ),
	.Selector15(\ALU|Selector15~8_combout ),
	.Selector12(\ALU|Selector12~10_combout ),
	.Selector13(\ALU|Selector13~8_combout ),
	.Selector10(\ALU|Selector10~8_combout ),
	.Selector11(\ALU|Selector11~9_combout ),
	.Selector8(\ALU|Selector8~10_combout ),
	.Selector9(\ALU|Selector9~8_combout ),
	.Selector6(\ALU|Selector6~8_combout ),
	.Selector7(\ALU|Selector7~11_combout ),
	.Selector4(\ALU|Selector4~10_combout ),
	.Selector5(\ALU|Selector5~8_combout ),
	.Selector2(\ALU|Selector2~11_combout ),
	.Selector3(\ALU|Selector3~11_combout ),
	.Selector0(\ALU|Selector0~34_combout ),
	.Selector1(\ALU|Selector1~20_combout ),
	.plif_exmemrdat2_l_1(plif_exmemrdat2_l_1),
	.plif_exmemrdat2_l_2(plif_exmemrdat2_l_2),
	.plif_exmemrdat2_l_3(plif_exmemrdat2_l_3),
	.plif_exmemrdat2_l_4(plif_exmemrdat2_l_4),
	.plif_exmemrdat2_l_5(plif_exmemrdat2_l_5),
	.plif_exmemrdat2_l_6(plif_exmemrdat2_l_6),
	.plif_exmemrdat2_l_7(plif_exmemrdat2_l_7),
	.plif_exmemrdat2_l_8(plif_exmemrdat2_l_8),
	.plif_exmemrdat2_l_9(plif_exmemrdat2_l_9),
	.plif_exmemrdat2_l_10(plif_exmemrdat2_l_10),
	.plif_exmemrdat2_l_11(plif_exmemrdat2_l_11),
	.plif_exmemrdat2_l_12(plif_exmemrdat2_l_12),
	.plif_exmemrdat2_l_13(plif_exmemrdat2_l_13),
	.plif_exmemrdat2_l_14(plif_exmemrdat2_l_14),
	.plif_exmemrdat2_l_15(plif_exmemrdat2_l_15),
	.plif_exmemrdat2_l_16(plif_exmemrdat2_l_16),
	.plif_exmemrdat2_l_17(plif_exmemrdat2_l_17),
	.plif_exmemrdat2_l_18(plif_exmemrdat2_l_18),
	.plif_exmemrdat2_l_19(plif_exmemrdat2_l_19),
	.plif_exmemrdat2_l_20(plif_exmemrdat2_l_20),
	.plif_exmemrdat2_l_21(plif_exmemrdat2_l_21),
	.plif_exmemrdat2_l_22(plif_exmemrdat2_l_22),
	.plif_exmemrdat2_l_23(plif_exmemrdat2_l_23),
	.plif_exmemrdat2_l_24(plif_exmemrdat2_l_24),
	.plif_exmemrdat2_l_25(plif_exmemrdat2_l_25),
	.plif_exmemrdat2_l_26(plif_exmemrdat2_l_26),
	.plif_exmemrdat2_l_27(plif_exmemrdat2_l_27),
	.plif_exmemrdat2_l_28(plif_exmemrdat2_l_28),
	.plif_exmemrdat2_l_29(plif_exmemrdat2_l_29),
	.plif_exmemrdat2_l_30(plif_exmemrdat2_l_30),
	.plif_exmemrdat2_l_31(plif_exmemrdat2_l_31),
	.plif_idexregen_l(\IDEX|plif_idex.regen_l~q ),
	.plif_exmemregsrc_l_0(\EXMEM|plif_exmem.regsrc_l [0]),
	.plif_exmemregsrc_l_1(\EXMEM|plif_exmem.regsrc_l [1]),
	.plif_exmemrtnaddr_l_31(\EXMEM|plif_exmem.rtnaddr_l [31]),
	.plif_exmemrtnaddr_l_30(\EXMEM|plif_exmem.rtnaddr_l [30]),
	.plif_exmemrtnaddr_l_29(\EXMEM|plif_exmem.rtnaddr_l [29]),
	.plif_exmemrtnaddr_l_28(\EXMEM|plif_exmem.rtnaddr_l [28]),
	.plif_exmemrtnaddr_l_27(\EXMEM|plif_exmem.rtnaddr_l [27]),
	.plif_exmemrtnaddr_l_26(\EXMEM|plif_exmem.rtnaddr_l [26]),
	.plif_exmemrtnaddr_l_25(\EXMEM|plif_exmem.rtnaddr_l [25]),
	.plif_exmemrtnaddr_l_24(\EXMEM|plif_exmem.rtnaddr_l [24]),
	.plif_exmemrtnaddr_l_23(\EXMEM|plif_exmem.rtnaddr_l [23]),
	.plif_exmemrtnaddr_l_22(\EXMEM|plif_exmem.rtnaddr_l [22]),
	.plif_exmemrtnaddr_l_21(\EXMEM|plif_exmem.rtnaddr_l [21]),
	.plif_exmemrtnaddr_l_20(\EXMEM|plif_exmem.rtnaddr_l [20]),
	.plif_exmemrtnaddr_l_19(\EXMEM|plif_exmem.rtnaddr_l [19]),
	.plif_exmemrtnaddr_l_18(\EXMEM|plif_exmem.rtnaddr_l [18]),
	.plif_exmemrtnaddr_l_17(\EXMEM|plif_exmem.rtnaddr_l [17]),
	.plif_exmemrtnaddr_l_16(\EXMEM|plif_exmem.rtnaddr_l [16]),
	.plif_exmemrtnaddr_l_15(\EXMEM|plif_exmem.rtnaddr_l [15]),
	.plif_exmemrtnaddr_l_14(\EXMEM|plif_exmem.rtnaddr_l [14]),
	.plif_exmemrtnaddr_l_13(\EXMEM|plif_exmem.rtnaddr_l [13]),
	.plif_exmemrtnaddr_l_12(\EXMEM|plif_exmem.rtnaddr_l [12]),
	.plif_exmemrtnaddr_l_11(\EXMEM|plif_exmem.rtnaddr_l [11]),
	.plif_exmemrtnaddr_l_10(\EXMEM|plif_exmem.rtnaddr_l [10]),
	.plif_exmemrtnaddr_l_9(\EXMEM|plif_exmem.rtnaddr_l [9]),
	.plif_exmemrtnaddr_l_8(\EXMEM|plif_exmem.rtnaddr_l [8]),
	.plif_exmemrtnaddr_l_7(\EXMEM|plif_exmem.rtnaddr_l [7]),
	.plif_exmemrtnaddr_l_6(\EXMEM|plif_exmem.rtnaddr_l [6]),
	.plif_exmemrtnaddr_l_5(\EXMEM|plif_exmem.rtnaddr_l [5]),
	.plif_exmemrtnaddr_l_2(\EXMEM|plif_exmem.rtnaddr_l [2]),
	.plif_exmemrtnaddr_l_1(\EXMEM|plif_exmem.rtnaddr_l [1]),
	.plif_exmemrtnaddr_l_0(\EXMEM|plif_exmem.rtnaddr_l [0]),
	.plif_exmemrtnaddr_l_4(\EXMEM|plif_exmem.rtnaddr_l [4]),
	.plif_exmemrtnaddr_l_3(\EXMEM|plif_exmem.rtnaddr_l [3]),
	.plif_exmembtype_l(\EXMEM|plif_exmem.btype_l~q ),
	.plif_exmemzero_l(\EXMEM|plif_exmem.zero_l~q ),
	.plif_exmemjaddr_l_1(\EXMEM|plif_exmem.jaddr_l [1]),
	.plif_exmemextimm_l_1(\EXMEM|plif_exmem.extimm_l [1]),
	.plif_exmemextimm_l_0(\EXMEM|plif_exmem.extimm_l [0]),
	.plif_exmemjaddr_l_0(\EXMEM|plif_exmem.jaddr_l [0]),
	.plif_exmemjaddr_l_3(\EXMEM|plif_exmem.jaddr_l [3]),
	.plif_exmemextimm_l_3(\EXMEM|plif_exmem.extimm_l [3]),
	.plif_exmemextimm_l_2(\EXMEM|plif_exmem.extimm_l [2]),
	.plif_exmemjaddr_l_2(\EXMEM|plif_exmem.jaddr_l [2]),
	.plif_exmemjaddr_l_5(\EXMEM|plif_exmem.jaddr_l [5]),
	.plif_exmemextimm_l_5(\EXMEM|plif_exmem.extimm_l [5]),
	.plif_exmemextimm_l_4(\EXMEM|plif_exmem.extimm_l [4]),
	.plif_exmemjaddr_l_4(\EXMEM|plif_exmem.jaddr_l [4]),
	.plif_exmemjaddr_l_7(\EXMEM|plif_exmem.jaddr_l [7]),
	.plif_exmemextimm_l_7(\EXMEM|plif_exmem.extimm_l [7]),
	.plif_exmemextimm_l_6(\EXMEM|plif_exmem.extimm_l [6]),
	.plif_exmemjaddr_l_6(\EXMEM|plif_exmem.jaddr_l [6]),
	.plif_exmemjaddr_l_9(\EXMEM|plif_exmem.jaddr_l [9]),
	.plif_exmemextimm_l_9(\EXMEM|plif_exmem.extimm_l [9]),
	.plif_exmemextimm_l_8(\EXMEM|plif_exmem.extimm_l [8]),
	.plif_exmemjaddr_l_8(\EXMEM|plif_exmem.jaddr_l [8]),
	.plif_exmemjaddr_l_11(\EXMEM|plif_exmem.jaddr_l [11]),
	.plif_exmemextimm_l_11(\EXMEM|plif_exmem.extimm_l [11]),
	.plif_exmemextimm_l_10(\EXMEM|plif_exmem.extimm_l [10]),
	.plif_exmemjaddr_l_10(\EXMEM|plif_exmem.jaddr_l [10]),
	.plif_exmemjaddr_l_13(\EXMEM|plif_exmem.jaddr_l [13]),
	.plif_exmemextimm_l_13(\EXMEM|plif_exmem.extimm_l [13]),
	.plif_exmemextimm_l_12(\EXMEM|plif_exmem.extimm_l [12]),
	.plif_exmemjaddr_l_12(\EXMEM|plif_exmem.jaddr_l [12]),
	.plif_exmemjaddr_l_15(\EXMEM|plif_exmem.jaddr_l [15]),
	.plif_exmemextimm_l_15(\EXMEM|plif_exmem.extimm_l [15]),
	.plif_exmemextimm_l_14(\EXMEM|plif_exmem.extimm_l [14]),
	.plif_exmemjaddr_l_14(\EXMEM|plif_exmem.jaddr_l [14]),
	.plif_exmemjaddr_l_17(\EXMEM|plif_exmem.jaddr_l [17]),
	.plif_exmemextimm_l_17(\EXMEM|plif_exmem.extimm_l [17]),
	.plif_exmemextimm_l_16(\EXMEM|plif_exmem.extimm_l [16]),
	.plif_exmemjaddr_l_16(\EXMEM|plif_exmem.jaddr_l [16]),
	.plif_exmemjaddr_l_19(\EXMEM|plif_exmem.jaddr_l [19]),
	.plif_exmemextimm_l_19(\EXMEM|plif_exmem.extimm_l [19]),
	.plif_exmemextimm_l_18(\EXMEM|plif_exmem.extimm_l [18]),
	.plif_exmemjaddr_l_18(\EXMEM|plif_exmem.jaddr_l [18]),
	.plif_exmemjaddr_l_21(\EXMEM|plif_exmem.jaddr_l [21]),
	.plif_exmemextimm_l_21(\EXMEM|plif_exmem.extimm_l [21]),
	.plif_exmemextimm_l_20(\EXMEM|plif_exmem.extimm_l [20]),
	.plif_exmemjaddr_l_20(\EXMEM|plif_exmem.jaddr_l [20]),
	.plif_exmemjaddr_l_23(\EXMEM|plif_exmem.jaddr_l [23]),
	.plif_exmemextimm_l_23(\EXMEM|plif_exmem.extimm_l [23]),
	.plif_exmemextimm_l_22(\EXMEM|plif_exmem.extimm_l [22]),
	.plif_exmemjaddr_l_22(\EXMEM|plif_exmem.jaddr_l [22]),
	.plif_exmemjaddr_l_25(\EXMEM|plif_exmem.jaddr_l [25]),
	.plif_exmemextimm_l_25(\EXMEM|plif_exmem.extimm_l [25]),
	.plif_exmemextimm_l_24(\EXMEM|plif_exmem.extimm_l [24]),
	.plif_exmemjaddr_l_24(\EXMEM|plif_exmem.jaddr_l [24]),
	.plif_exmemextimm_l_27(\EXMEM|plif_exmem.extimm_l [27]),
	.plif_exmemextimm_l_26(\EXMEM|plif_exmem.extimm_l [26]),
	.plif_exmemextimm_l_29(\EXMEM|plif_exmem.extimm_l [29]),
	.plif_exmemextimm_l_28(\EXMEM|plif_exmem.extimm_l [28]),
	.plif_idexregsrc_l_0(\IDEX|plif_idex.regsrc_l [0]),
	.plif_idexregsrc_l_1(\IDEX|plif_idex.regsrc_l [1]),
	.plif_idexrtnaddr_l_31(\IDEX|plif_idex.rtnaddr_l [31]),
	.plif_idexrtnaddr_l_30(\IDEX|plif_idex.rtnaddr_l [30]),
	.plif_idexrtnaddr_l_29(\IDEX|plif_idex.rtnaddr_l [29]),
	.plif_idexrtnaddr_l_28(\IDEX|plif_idex.rtnaddr_l [28]),
	.plif_idexrtnaddr_l_27(\IDEX|plif_idex.rtnaddr_l [27]),
	.plif_idexrtnaddr_l_26(\IDEX|plif_idex.rtnaddr_l [26]),
	.plif_idexrtnaddr_l_25(\IDEX|plif_idex.rtnaddr_l [25]),
	.plif_idexrtnaddr_l_24(\IDEX|plif_idex.rtnaddr_l [24]),
	.plif_idexrtnaddr_l_23(\IDEX|plif_idex.rtnaddr_l [23]),
	.plif_idexrtnaddr_l_22(\IDEX|plif_idex.rtnaddr_l [22]),
	.plif_idexrtnaddr_l_21(\IDEX|plif_idex.rtnaddr_l [21]),
	.plif_idexrtnaddr_l_20(\IDEX|plif_idex.rtnaddr_l [20]),
	.plif_idexrtnaddr_l_19(\IDEX|plif_idex.rtnaddr_l [19]),
	.plif_idexrtnaddr_l_18(\IDEX|plif_idex.rtnaddr_l [18]),
	.plif_idexrtnaddr_l_17(\IDEX|plif_idex.rtnaddr_l [17]),
	.plif_idexrtnaddr_l_16(\IDEX|plif_idex.rtnaddr_l [16]),
	.plif_idexrtnaddr_l_15(\IDEX|plif_idex.rtnaddr_l [15]),
	.plif_idexrtnaddr_l_14(\IDEX|plif_idex.rtnaddr_l [14]),
	.plif_idexrtnaddr_l_13(\IDEX|plif_idex.rtnaddr_l [13]),
	.plif_idexrtnaddr_l_12(\IDEX|plif_idex.rtnaddr_l [12]),
	.plif_idexrtnaddr_l_11(\IDEX|plif_idex.rtnaddr_l [11]),
	.plif_idexrtnaddr_l_10(\IDEX|plif_idex.rtnaddr_l [10]),
	.plif_idexrtnaddr_l_9(\IDEX|plif_idex.rtnaddr_l [9]),
	.plif_idexrtnaddr_l_8(\IDEX|plif_idex.rtnaddr_l [8]),
	.plif_idexrtnaddr_l_7(\IDEX|plif_idex.rtnaddr_l [7]),
	.plif_idexrtnaddr_l_6(\IDEX|plif_idex.rtnaddr_l [6]),
	.plif_idexrtnaddr_l_5(\IDEX|plif_idex.rtnaddr_l [5]),
	.plif_idexrtnaddr_l_2(\IDEX|plif_idex.rtnaddr_l [2]),
	.plif_idexrtnaddr_l_1(\IDEX|plif_idex.rtnaddr_l [1]),
	.plif_idexrtnaddr_l_0(\IDEX|plif_idex.rtnaddr_l [0]),
	.plif_idexrtnaddr_l_4(\IDEX|plif_idex.rtnaddr_l [4]),
	.plif_idexrtnaddr_l_3(\IDEX|plif_idex.rtnaddr_l [3]),
	.plif_idexbtype_l(\IDEX|plif_idex.btype_l~q ),
	.WideOr1(\ALU|WideOr1~combout ),
	.plif_idexjaddr_l_1(\IDEX|plif_idex.jaddr_l [1]),
	.plif_idexjaddr_l_0(\IDEX|plif_idex.jaddr_l [0]),
	.plif_idexjaddr_l_3(\IDEX|plif_idex.jaddr_l [3]),
	.plif_idexjaddr_l_2(\IDEX|plif_idex.jaddr_l [2]),
	.plif_idexjaddr_l_5(\IDEX|plif_idex.jaddr_l [5]),
	.plif_idexjaddr_l_4(\IDEX|plif_idex.jaddr_l [4]),
	.plif_idexjaddr_l_7(\IDEX|plif_idex.jaddr_l [7]),
	.plif_idexjaddr_l_6(\IDEX|plif_idex.jaddr_l [6]),
	.plif_idexjaddr_l_9(\IDEX|plif_idex.jaddr_l [9]),
	.plif_idexjaddr_l_8(\IDEX|plif_idex.jaddr_l [8]),
	.plif_idexjaddr_l_11(\IDEX|plif_idex.jaddr_l [11]),
	.plif_idexjaddr_l_10(\IDEX|plif_idex.jaddr_l [10]),
	.plif_idexjaddr_l_13(\IDEX|plif_idex.jaddr_l [13]),
	.plif_idexjaddr_l_12(\IDEX|plif_idex.jaddr_l [12]),
	.plif_idexjaddr_l_15(\IDEX|plif_idex.jaddr_l [15]),
	.plif_idexjaddr_l_14(\IDEX|plif_idex.jaddr_l [14]),
	.plif_idexjaddr_l_17(\IDEX|plif_idex.jaddr_l [17]),
	.plif_idexjaddr_l_16(\IDEX|plif_idex.jaddr_l [16]),
	.plif_idexjaddr_l_19(\IDEX|plif_idex.jaddr_l [19]),
	.plif_idexjaddr_l_18(\IDEX|plif_idex.jaddr_l [18]),
	.plif_idexjaddr_l_21(\IDEX|plif_idex.jaddr_l [21]),
	.plif_idexjaddr_l_20(\IDEX|plif_idex.jaddr_l [20]),
	.plif_idexjaddr_l_23(\IDEX|plif_idex.jaddr_l [23]),
	.plif_idexjaddr_l_22(\IDEX|plif_idex.jaddr_l [22]),
	.plif_idexjaddr_l_25(\IDEX|plif_idex.jaddr_l [25]),
	.plif_idexjaddr_l_24(\IDEX|plif_idex.jaddr_l [24]),
	.rdat2(\rdat2~96_combout ),
	.rdat21(\rdat2~97_combout ),
	.rdat22(\rdat2~98_combout ),
	.rdat23(\rdat2~99_combout ),
	.rdat24(\rdat2~100_combout ),
	.rdat25(\rdat2~101_combout ),
	.rdat26(\rdat2~102_combout ),
	.rdat27(\rdat2~103_combout ),
	.rdat28(\rdat2~104_combout ),
	.rdat29(\rdat2~105_combout ),
	.rdat210(\rdat2~106_combout ),
	.rdat211(\rdat2~107_combout ),
	.rdat212(\rdat2~108_combout ),
	.rdat213(\rdat2~109_combout ),
	.rdat214(\rdat2~110_combout ),
	.rdat215(\rdat2~111_combout ),
	.rdat216(\rdat2~112_combout ),
	.rdat217(\rdat2~113_combout ),
	.rdat218(\rdat2~114_combout ),
	.rdat219(\rdat2~115_combout ),
	.rdat220(\rdat2~116_combout ),
	.rdat221(\rdat2~117_combout ),
	.rdat222(\rdat2~118_combout ),
	.rdat223(\rdat2~119_combout ),
	.rdat224(\rdat2~120_combout ),
	.rdat225(\rdat2~121_combout ),
	.rdat226(\rdat2~122_combout ),
	.rdat227(\rdat2~123_combout ),
	.rdat228(\rdat2~124_combout ),
	.rdat229(\rdat2~125_combout ),
	.rdat230(\rdat2~126_combout ),
	.rdat231(\rdat2~127_combout ),
	.CPUCLK(CLK),
	.nRST(nRST),
	.devpor(devpor),
	.devclrn(devclrn),
	.devoe(devoe));

pipeline_idex IDEX(
	.plif_exmemdmemWEN_l(plif_exmemdmemWEN_l),
	.plif_exmemdmemREN_l(plif_exmemdmemREN_l),
	.always1(always1),
	.plif_idexhlt_l(\IDEX|plif_idex.hlt_l~q ),
	.plif_memwbpcsrc_l_1(\MEMWB|plif_memwb.pcsrc_l [1]),
	.plif_memwbpcsrc_l_0(\MEMWB|plif_memwb.pcsrc_l [0]),
	.plif_idexpcsrc_l_1(\IDEX|plif_idex.pcsrc_l [1]),
	.plif_idexpcsrc_l_0(\IDEX|plif_idex.pcsrc_l [0]),
	.ifid_sRST(\HU|ifid_sRST~2_combout ),
	.plif_idexaluop_l_3(\IDEX|plif_idex.aluop_l [3]),
	.plif_idexaluop_l_2(\IDEX|plif_idex.aluop_l [2]),
	.plif_idexaluop_l_1(\IDEX|plif_idex.aluop_l [1]),
	.plif_idexaluop_l_0(\IDEX|plif_idex.aluop_l [0]),
	.plif_idexextimm_l_31(\IDEX|plif_idex.extimm_l [31]),
	.plif_idexalusrc_l(\IDEX|plif_idex.alusrc_l~q ),
	.plif_idexrsel2_l_1(\IDEX|plif_idex.rsel2_l [1]),
	.plif_idexrsel2_l_0(\IDEX|plif_idex.rsel2_l [0]),
	.plif_idexrsel2_l_2(\IDEX|plif_idex.rsel2_l [2]),
	.plif_idexrsel2_l_3(\IDEX|plif_idex.rsel2_l [3]),
	.plif_idexrsel2_l_4(\IDEX|plif_idex.rsel2_l [4]),
	.plif_idexrdat2_l_31(\IDEX|plif_idex.rdat2_l [31]),
	.plif_idexextimm_l_30(\IDEX|plif_idex.extimm_l [30]),
	.plif_idexrdat2_l_30(\IDEX|plif_idex.rdat2_l [30]),
	.plif_idexextimm_l_29(\IDEX|plif_idex.extimm_l [29]),
	.plif_idexrdat2_l_29(\IDEX|plif_idex.rdat2_l [29]),
	.plif_idexextimm_l_28(\IDEX|plif_idex.extimm_l [28]),
	.plif_idexrdat2_l_28(\IDEX|plif_idex.rdat2_l [28]),
	.plif_idexextimm_l_27(\IDEX|plif_idex.extimm_l [27]),
	.plif_idexrdat2_l_27(\IDEX|plif_idex.rdat2_l [27]),
	.plif_idexextimm_l_26(\IDEX|plif_idex.extimm_l [26]),
	.plif_idexrdat2_l_26(\IDEX|plif_idex.rdat2_l [26]),
	.plif_idexextimm_l_25(\IDEX|plif_idex.extimm_l [25]),
	.plif_idexrdat2_l_25(\IDEX|plif_idex.rdat2_l [25]),
	.plif_idexextimm_l_24(\IDEX|plif_idex.extimm_l [24]),
	.plif_idexrdat2_l_24(\IDEX|plif_idex.rdat2_l [24]),
	.plif_idexextimm_l_23(\IDEX|plif_idex.extimm_l [23]),
	.plif_idexrdat2_l_23(\IDEX|plif_idex.rdat2_l [23]),
	.plif_idexextimm_l_22(\IDEX|plif_idex.extimm_l [22]),
	.plif_idexrdat2_l_22(\IDEX|plif_idex.rdat2_l [22]),
	.plif_idexextimm_l_21(\IDEX|plif_idex.extimm_l [21]),
	.plif_idexrdat2_l_21(\IDEX|plif_idex.rdat2_l [21]),
	.plif_idexextimm_l_20(\IDEX|plif_idex.extimm_l [20]),
	.plif_idexrdat2_l_20(\IDEX|plif_idex.rdat2_l [20]),
	.plif_idexextimm_l_19(\IDEX|plif_idex.extimm_l [19]),
	.plif_idexrdat2_l_19(\IDEX|plif_idex.rdat2_l [19]),
	.plif_idexextimm_l_18(\IDEX|plif_idex.extimm_l [18]),
	.plif_idexrdat2_l_18(\IDEX|plif_idex.rdat2_l [18]),
	.plif_idexextimm_l_17(\IDEX|plif_idex.extimm_l [17]),
	.plif_idexrdat2_l_17(\IDEX|plif_idex.rdat2_l [17]),
	.plif_idexextimm_l_16(\IDEX|plif_idex.extimm_l [16]),
	.plif_idexrdat2_l_16(\IDEX|plif_idex.rdat2_l [16]),
	.plif_idexextimm_l_15(\IDEX|plif_idex.extimm_l [15]),
	.plif_idexrdat2_l_15(\IDEX|plif_idex.rdat2_l [15]),
	.plif_idexrdat2_l_14(\IDEX|plif_idex.rdat2_l [14]),
	.plif_idexextimm_l_14(\IDEX|plif_idex.extimm_l [14]),
	.plif_idexextimm_l_13(\IDEX|plif_idex.extimm_l [13]),
	.plif_idexrdat2_l_13(\IDEX|plif_idex.rdat2_l [13]),
	.plif_idexrdat2_l_12(\IDEX|plif_idex.rdat2_l [12]),
	.plif_idexextimm_l_12(\IDEX|plif_idex.extimm_l [12]),
	.plif_idexextimm_l_11(\IDEX|plif_idex.extimm_l [11]),
	.plif_idexrdat2_l_11(\IDEX|plif_idex.rdat2_l [11]),
	.plif_idexrdat2_l_10(\IDEX|plif_idex.rdat2_l [10]),
	.plif_idexextimm_l_10(\IDEX|plif_idex.extimm_l [10]),
	.plif_idexextimm_l_9(\IDEX|plif_idex.extimm_l [9]),
	.plif_idexrdat2_l_9(\IDEX|plif_idex.rdat2_l [9]),
	.plif_idexrdat2_l_8(\IDEX|plif_idex.rdat2_l [8]),
	.plif_idexextimm_l_8(\IDEX|plif_idex.extimm_l [8]),
	.plif_idexextimm_l_7(\IDEX|plif_idex.extimm_l [7]),
	.plif_idexrdat2_l_7(\IDEX|plif_idex.rdat2_l [7]),
	.plif_idexrdat2_l_6(\IDEX|plif_idex.rdat2_l [6]),
	.plif_idexextimm_l_6(\IDEX|plif_idex.extimm_l [6]),
	.plif_idexextimm_l_5(\IDEX|plif_idex.extimm_l [5]),
	.plif_idexrdat2_l_5(\IDEX|plif_idex.rdat2_l [5]),
	.plif_idexrsel1_l_4(\IDEX|plif_idex.rsel1_l [4]),
	.plif_idexrsel1_l_1(\IDEX|plif_idex.rsel1_l [1]),
	.plif_idexrsel1_l_0(\IDEX|plif_idex.rsel1_l [0]),
	.plif_idexrsel1_l_2(\IDEX|plif_idex.rsel1_l [2]),
	.plif_idexrsel1_l_3(\IDEX|plif_idex.rsel1_l [3]),
	.plif_idexrdat1_l_2(\IDEX|plif_idex.rdat1_l [2]),
	.plif_idexrdat1_l_1(\IDEX|plif_idex.rdat1_l [1]),
	.plif_idexrdat2_l_0(\IDEX|plif_idex.rdat2_l [0]),
	.plif_idexextimm_l_0(\IDEX|plif_idex.extimm_l [0]),
	.plif_idexextimm_l_1(\IDEX|plif_idex.extimm_l [1]),
	.plif_idexrdat2_l_1(\IDEX|plif_idex.rdat2_l [1]),
	.plif_idexrdat1_l_4(\IDEX|plif_idex.rdat1_l [4]),
	.plif_idexrdat1_l_3(\IDEX|plif_idex.rdat1_l [3]),
	.plif_idexrdat2_l_2(\IDEX|plif_idex.rdat2_l [2]),
	.plif_idexextimm_l_2(\IDEX|plif_idex.extimm_l [2]),
	.plif_idexrdat1_l_8(\IDEX|plif_idex.rdat1_l [8]),
	.plif_idexrdat1_l_7(\IDEX|plif_idex.rdat1_l [7]),
	.plif_idexrdat1_l_6(\IDEX|plif_idex.rdat1_l [6]),
	.plif_idexrdat1_l_5(\IDEX|plif_idex.rdat1_l [5]),
	.plif_idexextimm_l_3(\IDEX|plif_idex.extimm_l [3]),
	.plif_idexrdat2_l_3(\IDEX|plif_idex.rdat2_l [3]),
	.plif_idexrdat1_l_16(\IDEX|plif_idex.rdat1_l [16]),
	.plif_idexrdat1_l_15(\IDEX|plif_idex.rdat1_l [15]),
	.plif_idexrdat1_l_14(\IDEX|plif_idex.rdat1_l [14]),
	.plif_idexrdat1_l_13(\IDEX|plif_idex.rdat1_l [13]),
	.plif_idexrdat1_l_12(\IDEX|plif_idex.rdat1_l [12]),
	.plif_idexrdat1_l_11(\IDEX|plif_idex.rdat1_l [11]),
	.plif_idexrdat1_l_10(\IDEX|plif_idex.rdat1_l [10]),
	.plif_idexrdat1_l_9(\IDEX|plif_idex.rdat1_l [9]),
	.plif_idexrdat2_l_4(\IDEX|plif_idex.rdat2_l [4]),
	.plif_idexextimm_l_4(\IDEX|plif_idex.extimm_l [4]),
	.plif_idexrdat1_l_31(\IDEX|plif_idex.rdat1_l [31]),
	.plif_idexrdat1_l_29(\IDEX|plif_idex.rdat1_l [29]),
	.plif_idexrdat1_l_30(\IDEX|plif_idex.rdat1_l [30]),
	.plif_idexrdat1_l_28(\IDEX|plif_idex.rdat1_l [28]),
	.plif_idexrdat1_l_27(\IDEX|plif_idex.rdat1_l [27]),
	.plif_idexrdat1_l_26(\IDEX|plif_idex.rdat1_l [26]),
	.plif_idexrdat1_l_25(\IDEX|plif_idex.rdat1_l [25]),
	.plif_idexrdat1_l_24(\IDEX|plif_idex.rdat1_l [24]),
	.plif_idexrdat1_l_23(\IDEX|plif_idex.rdat1_l [23]),
	.plif_idexrdat1_l_22(\IDEX|plif_idex.rdat1_l [22]),
	.plif_idexrdat1_l_21(\IDEX|plif_idex.rdat1_l [21]),
	.plif_idexrdat1_l_20(\IDEX|plif_idex.rdat1_l [20]),
	.plif_idexrdat1_l_19(\IDEX|plif_idex.rdat1_l [19]),
	.plif_idexrdat1_l_18(\IDEX|plif_idex.rdat1_l [18]),
	.plif_idexrdat1_l_17(\IDEX|plif_idex.rdat1_l [17]),
	.plif_idexrdat1_l_0(\IDEX|plif_idex.rdat1_l [0]),
	.plif_idexdmemREN_l(\IDEX|plif_idex.dmemREN_l~q ),
	.plif_idexwsel_l_0(\IDEX|plif_idex.wsel_l [0]),
	.plif_idexwsel_l_1(\IDEX|plif_idex.wsel_l [1]),
	.plif_ifidinstr_l_31(\IFID|plif_ifid.instr_l [31]),
	.plif_ifidinstr_l_29(\IFID|plif_ifid.instr_l [29]),
	.plif_ifidinstr_l_27(\IFID|plif_ifid.instr_l [27]),
	.plif_ifidinstr_l_26(\IFID|plif_ifid.instr_l [26]),
	.plif_ifidinstr_l_28(\IFID|plif_ifid.instr_l [28]),
	.Equal16(\CU|Equal16~0_combout ),
	.plif_ifidinstr_l_30(\IFID|plif_ifid.instr_l [30]),
	.Equal22(\CU|Equal22~0_combout ),
	.plif_ifidinstr_l_5(\IFID|plif_ifid.instr_l [5]),
	.plif_ifidinstr_l_1(\IFID|plif_ifid.instr_l [1]),
	.plif_ifidinstr_l_0(\IFID|plif_ifid.instr_l [0]),
	.plif_ifidinstr_l_2(\IFID|plif_ifid.instr_l [2]),
	.plif_ifidinstr_l_3(\IFID|plif_ifid.instr_l [3]),
	.WideNor0(\CU|WideNor0~2_combout ),
	.Equal11(\CU|Equal11~0_combout ),
	.Equal26(\CU|Equal26~0_combout ),
	.plif_ifidinstr_l_4(\IFID|plif_ifid.instr_l [4]),
	.Equal21(\CU|Equal21~0_combout ),
	.WideOr14(\CU|WideOr14~0_combout ),
	.Equal13(\CU|Equal13~1_combout ),
	.aluop_l(\IDEX|aluop_l~0_combout ),
	.WideNor1(\CU|WideNor1~0_combout ),
	.Selector22(\CU|Selector22~6_combout ),
	.Selector4(\CU|Selector4~0_combout ),
	.plif_ifidinstr_l_22(\IFID|plif_ifid.instr_l [22]),
	.plif_ifidinstr_l_21(\IFID|plif_ifid.instr_l [21]),
	.plif_idexwsel_l_2(\IDEX|plif_idex.wsel_l [2]),
	.plif_idexwsel_l_3(\IDEX|plif_idex.wsel_l [3]),
	.plif_ifidinstr_l_24(\IFID|plif_ifid.instr_l [24]),
	.plif_ifidinstr_l_23(\IFID|plif_ifid.instr_l [23]),
	.plif_idexwsel_l_4(\IDEX|plif_idex.wsel_l [4]),
	.plif_ifidinstr_l_25(\IFID|plif_ifid.instr_l [25]),
	.Selector1(\CU|Selector1~0_combout ),
	.Equal6(\CU|Equal6~0_combout ),
	.Selector11(\CU|Selector11~0_combout ),
	.Selector21(\CU|Selector21~0_combout ),
	.Selector9(\CU|Selector9~0_combout ),
	.plif_ifidinstr_l_17(\IFID|plif_ifid.instr_l [17]),
	.plif_ifidinstr_l_16(\IFID|plif_ifid.instr_l [16]),
	.plif_ifidinstr_l_19(\IFID|plif_ifid.instr_l [19]),
	.plif_ifidinstr_l_18(\IFID|plif_ifid.instr_l [18]),
	.plif_ifidinstr_l_20(\IFID|plif_ifid.instr_l [20]),
	.Selector6(\CU|Selector6~0_combout ),
	.plif_idexdmemWEN_l(\IDEX|plif_idex.dmemWEN_l~q ),
	.Equal23(\CU|Equal23~0_combout ),
	.idex_sRST(\HU|idex_sRST~3_combout ),
	.idex_sRST1(\HU|idex_sRST~4_combout ),
	.pcsrc(\CU|pcsrc~0_combout ),
	.Equal1(\CU|Equal1~0_combout ),
	.Equal20(\CU|Equal20~0_combout ),
	.WideNor11(\CU|WideNor1~1_combout ),
	.Equal19(\CU|Equal19~0_combout ),
	.Equal12(\CU|Equal1~1_combout ),
	.Equal18(\CU|Equal18~0_combout ),
	.Selector221(\CU|Selector22~7_combout ),
	.plif_ifidinstr_l_15(\IFID|plif_ifid.instr_l [15]),
	.WideOr141(\CU|WideOr14~combout ),
	.WideOr15(\CU|WideOr15~combout ),
	.WideOr16(\CU|WideOr16~0_combout ),
	.plif_idexregen_l(\IDEX|plif_idex.regen_l~q ),
	.Mux32(\RF|Mux32~9_combout ),
	.Mux321(\RF|Mux32~19_combout ),
	.extimm_30(\extimm[30]~0_combout ),
	.plif_ifidinstr_l_14(\IFID|plif_ifid.instr_l [14]),
	.Equal0(\Equal0~0_combout ),
	.Mux33(\RF|Mux33~9_combout ),
	.Mux331(\RF|Mux33~19_combout ),
	.plif_ifidinstr_l_13(\IFID|plif_ifid.instr_l [13]),
	.Mux34(\RF|Mux34~9_combout ),
	.Mux341(\RF|Mux34~19_combout ),
	.plif_ifidinstr_l_12(\IFID|plif_ifid.instr_l [12]),
	.Mux35(\RF|Mux35~9_combout ),
	.Mux351(\RF|Mux35~19_combout ),
	.plif_ifidinstr_l_11(\IFID|plif_ifid.instr_l [11]),
	.Mux36(\RF|Mux36~9_combout ),
	.Mux361(\RF|Mux36~19_combout ),
	.plif_ifidinstr_l_10(\IFID|plif_ifid.instr_l [10]),
	.Mux37(\RF|Mux37~9_combout ),
	.Mux371(\RF|Mux37~19_combout ),
	.plif_ifidinstr_l_9(\IFID|plif_ifid.instr_l [9]),
	.Mux38(\RF|Mux38~9_combout ),
	.Mux381(\RF|Mux38~19_combout ),
	.plif_ifidinstr_l_8(\IFID|plif_ifid.instr_l [8]),
	.Mux39(\RF|Mux39~9_combout ),
	.Mux391(\RF|Mux39~19_combout ),
	.plif_ifidinstr_l_7(\IFID|plif_ifid.instr_l [7]),
	.Mux40(\RF|Mux40~9_combout ),
	.Mux401(\RF|Mux40~19_combout ),
	.plif_ifidinstr_l_6(\IFID|plif_ifid.instr_l [6]),
	.Mux41(\RF|Mux41~9_combout ),
	.Mux411(\RF|Mux41~19_combout ),
	.Mux42(\RF|Mux42~9_combout ),
	.Mux421(\RF|Mux42~19_combout ),
	.Selector14(\CU|Selector14~0_combout ),
	.Mux43(\RF|Mux43~9_combout ),
	.Mux431(\RF|Mux43~19_combout ),
	.Selector15(\CU|Selector15~0_combout ),
	.Mux44(\RF|Mux44~9_combout ),
	.Mux441(\RF|Mux44~19_combout ),
	.Selector16(\CU|Selector16~0_combout ),
	.Mux45(\RF|Mux45~9_combout ),
	.Mux451(\RF|Mux45~19_combout ),
	.Selector17(\CU|Selector17~0_combout ),
	.Mux46(\RF|Mux46~9_combout ),
	.Mux461(\RF|Mux46~19_combout ),
	.Selector18(\CU|Selector18~0_combout ),
	.Mux47(\RF|Mux47~9_combout ),
	.Mux471(\RF|Mux47~19_combout ),
	.Mux48(\RF|Mux48~9_combout ),
	.Mux481(\RF|Mux48~19_combout ),
	.Mux49(\RF|Mux49~9_combout ),
	.Mux491(\RF|Mux49~19_combout ),
	.Mux50(\RF|Mux50~9_combout ),
	.Mux501(\RF|Mux50~19_combout ),
	.Mux51(\RF|Mux51~9_combout ),
	.Mux511(\RF|Mux51~19_combout ),
	.Mux52(\RF|Mux52~9_combout ),
	.Mux521(\RF|Mux52~19_combout ),
	.Mux53(\RF|Mux53~9_combout ),
	.Mux531(\RF|Mux53~19_combout ),
	.Mux54(\RF|Mux54~9_combout ),
	.Mux541(\RF|Mux54~19_combout ),
	.Mux55(\RF|Mux55~9_combout ),
	.Mux551(\RF|Mux55~19_combout ),
	.Mux56(\RF|Mux56~9_combout ),
	.Mux561(\RF|Mux56~19_combout ),
	.Mux57(\RF|Mux57~9_combout ),
	.Mux571(\RF|Mux57~19_combout ),
	.Mux58(\RF|Mux58~9_combout ),
	.Mux581(\RF|Mux58~19_combout ),
	.Mux29(\RF|Mux29~9_combout ),
	.Mux291(\RF|Mux29~19_combout ),
	.Mux30(\RF|Mux30~9_combout ),
	.Mux301(\RF|Mux30~19_combout ),
	.Mux63(\RF|Mux63~9_combout ),
	.Mux631(\RF|Mux63~19_combout ),
	.Mux62(\RF|Mux62~9_combout ),
	.Mux621(\RF|Mux62~19_combout ),
	.Mux27(\RF|Mux27~9_combout ),
	.Mux271(\RF|Mux27~19_combout ),
	.Mux28(\RF|Mux28~9_combout ),
	.Mux281(\RF|Mux28~19_combout ),
	.Mux61(\RF|Mux61~9_combout ),
	.Mux611(\RF|Mux61~19_combout ),
	.Mux23(\RF|Mux23~9_combout ),
	.Mux231(\RF|Mux23~19_combout ),
	.Mux24(\RF|Mux24~9_combout ),
	.Mux241(\RF|Mux24~19_combout ),
	.Mux25(\RF|Mux25~9_combout ),
	.Mux251(\RF|Mux25~19_combout ),
	.Mux26(\RF|Mux26~9_combout ),
	.Mux261(\RF|Mux26~19_combout ),
	.Mux60(\RF|Mux60~9_combout ),
	.Mux601(\RF|Mux60~19_combout ),
	.Mux15(\RF|Mux15~9_combout ),
	.Mux151(\RF|Mux15~19_combout ),
	.Mux16(\RF|Mux16~9_combout ),
	.Mux161(\RF|Mux16~19_combout ),
	.Mux17(\RF|Mux17~9_combout ),
	.Mux171(\RF|Mux17~19_combout ),
	.Mux18(\RF|Mux18~9_combout ),
	.Mux181(\RF|Mux18~19_combout ),
	.Mux19(\RF|Mux19~9_combout ),
	.Mux191(\RF|Mux19~19_combout ),
	.Mux20(\RF|Mux20~9_combout ),
	.Mux201(\RF|Mux20~19_combout ),
	.Mux21(\RF|Mux21~9_combout ),
	.Mux211(\RF|Mux21~19_combout ),
	.Mux22(\RF|Mux22~9_combout ),
	.Mux221(\RF|Mux22~19_combout ),
	.Mux59(\RF|Mux59~9_combout ),
	.Mux591(\RF|Mux59~19_combout ),
	.Mux0(\RF|Mux0~9_combout ),
	.Mux01(\RF|Mux0~19_combout ),
	.Mux2(\RF|Mux2~9_combout ),
	.Mux210(\RF|Mux2~19_combout ),
	.Mux1(\RF|Mux1~9_combout ),
	.Mux11(\RF|Mux1~19_combout ),
	.Mux3(\RF|Mux3~9_combout ),
	.Mux31(\RF|Mux3~19_combout ),
	.Mux4(\RF|Mux4~9_combout ),
	.Mux410(\RF|Mux4~19_combout ),
	.Mux5(\RF|Mux5~9_combout ),
	.Mux510(\RF|Mux5~19_combout ),
	.Mux6(\RF|Mux6~9_combout ),
	.Mux64(\RF|Mux6~19_combout ),
	.Mux7(\RF|Mux7~9_combout ),
	.Mux71(\RF|Mux7~19_combout ),
	.Mux8(\RF|Mux8~9_combout ),
	.Mux81(\RF|Mux8~19_combout ),
	.Mux9(\RF|Mux9~9_combout ),
	.Mux91(\RF|Mux9~19_combout ),
	.Mux10(\RF|Mux10~9_combout ),
	.Mux101(\RF|Mux10~19_combout ),
	.Mux111(\RF|Mux11~9_combout ),
	.Mux112(\RF|Mux11~19_combout ),
	.Mux12(\RF|Mux12~9_combout ),
	.Mux121(\RF|Mux12~19_combout ),
	.Mux13(\RF|Mux13~9_combout ),
	.Mux131(\RF|Mux13~19_combout ),
	.Mux14(\RF|Mux14~9_combout ),
	.Mux141(\RF|Mux14~19_combout ),
	.Mux311(\RF|Mux31~9_combout ),
	.Mux312(\RF|Mux31~19_combout ),
	.Selector24(\CU|Selector24~0_combout ),
	.plif_idexregsrc_l_0(\IDEX|plif_idex.regsrc_l [0]),
	.plif_idexregsrc_l_1(\IDEX|plif_idex.regsrc_l [1]),
	.plif_idexrtnaddr_l_31(\IDEX|plif_idex.rtnaddr_l [31]),
	.plif_idexrtnaddr_l_30(\IDEX|plif_idex.rtnaddr_l [30]),
	.plif_idexrtnaddr_l_29(\IDEX|plif_idex.rtnaddr_l [29]),
	.plif_idexrtnaddr_l_28(\IDEX|plif_idex.rtnaddr_l [28]),
	.plif_idexrtnaddr_l_27(\IDEX|plif_idex.rtnaddr_l [27]),
	.plif_idexrtnaddr_l_26(\IDEX|plif_idex.rtnaddr_l [26]),
	.plif_idexrtnaddr_l_25(\IDEX|plif_idex.rtnaddr_l [25]),
	.plif_idexrtnaddr_l_24(\IDEX|plif_idex.rtnaddr_l [24]),
	.plif_idexrtnaddr_l_23(\IDEX|plif_idex.rtnaddr_l [23]),
	.plif_idexrtnaddr_l_22(\IDEX|plif_idex.rtnaddr_l [22]),
	.plif_idexrtnaddr_l_21(\IDEX|plif_idex.rtnaddr_l [21]),
	.plif_idexrtnaddr_l_20(\IDEX|plif_idex.rtnaddr_l [20]),
	.plif_idexrtnaddr_l_19(\IDEX|plif_idex.rtnaddr_l [19]),
	.plif_idexrtnaddr_l_18(\IDEX|plif_idex.rtnaddr_l [18]),
	.plif_idexrtnaddr_l_17(\IDEX|plif_idex.rtnaddr_l [17]),
	.plif_idexrtnaddr_l_16(\IDEX|plif_idex.rtnaddr_l [16]),
	.plif_idexrtnaddr_l_15(\IDEX|plif_idex.rtnaddr_l [15]),
	.plif_idexrtnaddr_l_14(\IDEX|plif_idex.rtnaddr_l [14]),
	.plif_idexrtnaddr_l_13(\IDEX|plif_idex.rtnaddr_l [13]),
	.plif_idexrtnaddr_l_12(\IDEX|plif_idex.rtnaddr_l [12]),
	.plif_idexrtnaddr_l_11(\IDEX|plif_idex.rtnaddr_l [11]),
	.plif_idexrtnaddr_l_10(\IDEX|plif_idex.rtnaddr_l [10]),
	.plif_idexrtnaddr_l_9(\IDEX|plif_idex.rtnaddr_l [9]),
	.plif_idexrtnaddr_l_8(\IDEX|plif_idex.rtnaddr_l [8]),
	.plif_idexrtnaddr_l_7(\IDEX|plif_idex.rtnaddr_l [7]),
	.plif_idexrtnaddr_l_6(\IDEX|plif_idex.rtnaddr_l [6]),
	.plif_idexrtnaddr_l_5(\IDEX|plif_idex.rtnaddr_l [5]),
	.plif_idexrtnaddr_l_2(\IDEX|plif_idex.rtnaddr_l [2]),
	.plif_idexrtnaddr_l_1(\IDEX|plif_idex.rtnaddr_l [1]),
	.plif_idexrtnaddr_l_0(\IDEX|plif_idex.rtnaddr_l [0]),
	.plif_idexrtnaddr_l_4(\IDEX|plif_idex.rtnaddr_l [4]),
	.plif_idexrtnaddr_l_3(\IDEX|plif_idex.rtnaddr_l [3]),
	.plif_idexbtype_l(\IDEX|plif_idex.btype_l~q ),
	.plif_idexjaddr_l_1(\IDEX|plif_idex.jaddr_l [1]),
	.plif_idexjaddr_l_0(\IDEX|plif_idex.jaddr_l [0]),
	.plif_idexjaddr_l_3(\IDEX|plif_idex.jaddr_l [3]),
	.plif_idexjaddr_l_2(\IDEX|plif_idex.jaddr_l [2]),
	.plif_idexjaddr_l_5(\IDEX|plif_idex.jaddr_l [5]),
	.plif_idexjaddr_l_4(\IDEX|plif_idex.jaddr_l [4]),
	.plif_idexjaddr_l_7(\IDEX|plif_idex.jaddr_l [7]),
	.plif_idexjaddr_l_6(\IDEX|plif_idex.jaddr_l [6]),
	.plif_idexjaddr_l_9(\IDEX|plif_idex.jaddr_l [9]),
	.plif_idexjaddr_l_8(\IDEX|plif_idex.jaddr_l [8]),
	.plif_idexjaddr_l_11(\IDEX|plif_idex.jaddr_l [11]),
	.plif_idexjaddr_l_10(\IDEX|plif_idex.jaddr_l [10]),
	.plif_idexjaddr_l_13(\IDEX|plif_idex.jaddr_l [13]),
	.plif_idexjaddr_l_12(\IDEX|plif_idex.jaddr_l [12]),
	.plif_idexjaddr_l_15(\IDEX|plif_idex.jaddr_l [15]),
	.plif_idexjaddr_l_14(\IDEX|plif_idex.jaddr_l [14]),
	.plif_idexjaddr_l_17(\IDEX|plif_idex.jaddr_l [17]),
	.plif_idexjaddr_l_16(\IDEX|plif_idex.jaddr_l [16]),
	.plif_idexjaddr_l_19(\IDEX|plif_idex.jaddr_l [19]),
	.plif_idexjaddr_l_18(\IDEX|plif_idex.jaddr_l [18]),
	.plif_idexjaddr_l_21(\IDEX|plif_idex.jaddr_l [21]),
	.plif_idexjaddr_l_20(\IDEX|plif_idex.jaddr_l [20]),
	.plif_idexjaddr_l_23(\IDEX|plif_idex.jaddr_l [23]),
	.plif_idexjaddr_l_22(\IDEX|plif_idex.jaddr_l [22]),
	.plif_idexjaddr_l_25(\IDEX|plif_idex.jaddr_l [25]),
	.plif_idexjaddr_l_24(\IDEX|plif_idex.jaddr_l [24]),
	.plif_ifidrtnaddr_l_31(\IFID|plif_ifid.rtnaddr_l [31]),
	.plif_ifidrtnaddr_l_30(\IFID|plif_ifid.rtnaddr_l [30]),
	.plif_ifidrtnaddr_l_29(\IFID|plif_ifid.rtnaddr_l [29]),
	.plif_ifidrtnaddr_l_28(\IFID|plif_ifid.rtnaddr_l [28]),
	.plif_ifidrtnaddr_l_27(\IFID|plif_ifid.rtnaddr_l [27]),
	.plif_ifidrtnaddr_l_26(\IFID|plif_ifid.rtnaddr_l [26]),
	.plif_ifidrtnaddr_l_25(\IFID|plif_ifid.rtnaddr_l [25]),
	.plif_ifidrtnaddr_l_24(\IFID|plif_ifid.rtnaddr_l [24]),
	.plif_ifidrtnaddr_l_23(\IFID|plif_ifid.rtnaddr_l [23]),
	.plif_ifidrtnaddr_l_22(\IFID|plif_ifid.rtnaddr_l [22]),
	.plif_ifidrtnaddr_l_21(\IFID|plif_ifid.rtnaddr_l [21]),
	.plif_ifidrtnaddr_l_20(\IFID|plif_ifid.rtnaddr_l [20]),
	.plif_ifidrtnaddr_l_19(\IFID|plif_ifid.rtnaddr_l [19]),
	.plif_ifidrtnaddr_l_18(\IFID|plif_ifid.rtnaddr_l [18]),
	.plif_ifidrtnaddr_l_17(\IFID|plif_ifid.rtnaddr_l [17]),
	.plif_ifidrtnaddr_l_16(\IFID|plif_ifid.rtnaddr_l [16]),
	.plif_ifidrtnaddr_l_15(\IFID|plif_ifid.rtnaddr_l [15]),
	.plif_ifidrtnaddr_l_14(\IFID|plif_ifid.rtnaddr_l [14]),
	.plif_ifidrtnaddr_l_13(\IFID|plif_ifid.rtnaddr_l [13]),
	.plif_ifidrtnaddr_l_12(\IFID|plif_ifid.rtnaddr_l [12]),
	.plif_ifidrtnaddr_l_11(\IFID|plif_ifid.rtnaddr_l [11]),
	.plif_ifidrtnaddr_l_10(\IFID|plif_ifid.rtnaddr_l [10]),
	.plif_ifidrtnaddr_l_9(\IFID|plif_ifid.rtnaddr_l [9]),
	.plif_ifidrtnaddr_l_8(\IFID|plif_ifid.rtnaddr_l [8]),
	.plif_ifidrtnaddr_l_7(\IFID|plif_ifid.rtnaddr_l [7]),
	.plif_ifidrtnaddr_l_6(\IFID|plif_ifid.rtnaddr_l [6]),
	.plif_ifidrtnaddr_l_5(\IFID|plif_ifid.rtnaddr_l [5]),
	.plif_ifidrtnaddr_l_2(\IFID|plif_ifid.rtnaddr_l [2]),
	.plif_ifidrtnaddr_l_1(\IFID|plif_ifid.rtnaddr_l [1]),
	.plif_ifidrtnaddr_l_0(\IFID|plif_ifid.rtnaddr_l [0]),
	.plif_ifidrtnaddr_l_4(\IFID|plif_ifid.rtnaddr_l [4]),
	.plif_ifidrtnaddr_l_3(\IFID|plif_ifid.rtnaddr_l [3]),
	.Equal121(\CU|Equal12~0_combout ),
	.idex_sRST2(\HU|idex_sRST~5_combout ),
	.Selector0(\CU|Selector0~2_combout ),
	.Equal25(\CU|Equal25~4_combout ),
	.CPUCLK(CLK),
	.nRST(nRST),
	.devpor(devpor),
	.devclrn(devclrn),
	.devoe(devoe));

pipeline_ifid IFID(
	.PCreg_1(PCreg_1),
	.PCreg_0(PCreg_0),
	.pcifrtnaddr_2(\PC|pcif.rtnaddr[2]~0_combout ),
	.pcifrtnaddr_3(\PC|pcif.rtnaddr[3]~2_combout ),
	.pcifrtnaddr_4(\PC|pcif.rtnaddr[4]~4_combout ),
	.pcifrtnaddr_5(\PC|pcif.rtnaddr[5]~6_combout ),
	.pcifrtnaddr_6(\PC|pcif.rtnaddr[6]~8_combout ),
	.pcifrtnaddr_7(\PC|pcif.rtnaddr[7]~10_combout ),
	.pcifrtnaddr_8(\PC|pcif.rtnaddr[8]~12_combout ),
	.pcifrtnaddr_9(\PC|pcif.rtnaddr[9]~14_combout ),
	.pcifrtnaddr_10(\PC|pcif.rtnaddr[10]~16_combout ),
	.pcifrtnaddr_11(\PC|pcif.rtnaddr[11]~18_combout ),
	.pcifrtnaddr_12(\PC|pcif.rtnaddr[12]~20_combout ),
	.pcifrtnaddr_13(\PC|pcif.rtnaddr[13]~22_combout ),
	.pcifrtnaddr_14(\PC|pcif.rtnaddr[14]~24_combout ),
	.pcifrtnaddr_15(\PC|pcif.rtnaddr[15]~26_combout ),
	.pcifrtnaddr_16(\PC|pcif.rtnaddr[16]~28_combout ),
	.pcifrtnaddr_17(\PC|pcif.rtnaddr[17]~30_combout ),
	.pcifrtnaddr_18(\PC|pcif.rtnaddr[18]~32_combout ),
	.pcifrtnaddr_19(\PC|pcif.rtnaddr[19]~34_combout ),
	.pcifrtnaddr_20(\PC|pcif.rtnaddr[20]~36_combout ),
	.pcifrtnaddr_21(\PC|pcif.rtnaddr[21]~38_combout ),
	.pcifrtnaddr_22(\PC|pcif.rtnaddr[22]~40_combout ),
	.pcifrtnaddr_23(\PC|pcif.rtnaddr[23]~42_combout ),
	.pcifrtnaddr_24(\PC|pcif.rtnaddr[24]~44_combout ),
	.pcifrtnaddr_25(\PC|pcif.rtnaddr[25]~46_combout ),
	.pcifrtnaddr_26(\PC|pcif.rtnaddr[26]~48_combout ),
	.pcifrtnaddr_27(\PC|pcif.rtnaddr[27]~50_combout ),
	.pcifrtnaddr_28(\PC|pcif.rtnaddr[28]~52_combout ),
	.pcifrtnaddr_29(\PC|pcif.rtnaddr[29]~54_combout ),
	.pcifrtnaddr_30(\PC|pcif.rtnaddr[30]~56_combout ),
	.pcifrtnaddr_31(\PC|pcif.rtnaddr[31]~58_combout ),
	.ramiframload_0(ramiframload_0),
	.ramiframload_1(ramiframload_1),
	.ramiframload_2(ramiframload_2),
	.ramiframload_3(ramiframload_3),
	.ramiframload_4(ramiframload_4),
	.ramiframload_5(ramiframload_5),
	.ramiframload_6(ramiframload_6),
	.ramiframload_7(ramiframload_7),
	.ramiframload_8(ramiframload_8),
	.ramiframload_9(ramiframload_9),
	.ramiframload_10(ramiframload_10),
	.ramiframload_11(ramiframload_11),
	.ramiframload_12(ramiframload_12),
	.ramiframload_13(ramiframload_13),
	.ramiframload_14(ramiframload_14),
	.ramiframload_15(ramiframload_15),
	.ramiframload_16(ramiframload_16),
	.ramiframload_17(ramiframload_17),
	.ramiframload_18(ramiframload_18),
	.ramiframload_19(ramiframload_19),
	.ramiframload_20(ramiframload_20),
	.ramiframload_21(ramiframload_21),
	.ramiframload_22(ramiframload_22),
	.ramiframload_23(ramiframload_23),
	.ramiframload_24(ramiframload_24),
	.ramiframload_25(ramiframload_25),
	.ramiframload_26(ramiframload_26),
	.ramiframload_27(ramiframload_27),
	.ramiframload_28(ramiframload_28),
	.ramiframload_29(ramiframload_29),
	.ramiframload_30(ramiframload_30),
	.ramiframload_31(ramiframload_31),
	.plif_ifidinstr_l_31(\IFID|plif_ifid.instr_l [31]),
	.plif_ifidinstr_l_29(\IFID|plif_ifid.instr_l [29]),
	.plif_ifidinstr_l_27(\IFID|plif_ifid.instr_l [27]),
	.plif_ifidinstr_l_26(\IFID|plif_ifid.instr_l [26]),
	.plif_ifidinstr_l_28(\IFID|plif_ifid.instr_l [28]),
	.plif_ifidinstr_l_30(\IFID|plif_ifid.instr_l [30]),
	.plif_ifidinstr_l_5(\IFID|plif_ifid.instr_l [5]),
	.plif_ifidinstr_l_1(\IFID|plif_ifid.instr_l [1]),
	.plif_ifidinstr_l_0(\IFID|plif_ifid.instr_l [0]),
	.plif_ifidinstr_l_2(\IFID|plif_ifid.instr_l [2]),
	.plif_ifidinstr_l_3(\IFID|plif_ifid.instr_l [3]),
	.plif_ifidinstr_l_4(\IFID|plif_ifid.instr_l [4]),
	.plif_ifidinstr_l_22(\IFID|plif_ifid.instr_l [22]),
	.plif_ifidinstr_l_21(\IFID|plif_ifid.instr_l [21]),
	.plif_ifidinstr_l_24(\IFID|plif_ifid.instr_l [24]),
	.plif_ifidinstr_l_23(\IFID|plif_ifid.instr_l [23]),
	.plif_ifidinstr_l_25(\IFID|plif_ifid.instr_l [25]),
	.plif_ifidinstr_l_17(\IFID|plif_ifid.instr_l [17]),
	.plif_ifidinstr_l_16(\IFID|plif_ifid.instr_l [16]),
	.plif_ifidinstr_l_19(\IFID|plif_ifid.instr_l [19]),
	.plif_ifidinstr_l_18(\IFID|plif_ifid.instr_l [18]),
	.plif_ifidinstr_l_20(\IFID|plif_ifid.instr_l [20]),
	.ifid_en(\HU|ifid_en~0_combout ),
	.plif_ifidinstr_l_15(\IFID|plif_ifid.instr_l [15]),
	.plif_ifidinstr_l_14(\IFID|plif_ifid.instr_l [14]),
	.plif_ifidinstr_l_13(\IFID|plif_ifid.instr_l [13]),
	.plif_ifidinstr_l_12(\IFID|plif_ifid.instr_l [12]),
	.plif_ifidinstr_l_11(\IFID|plif_ifid.instr_l [11]),
	.plif_ifidinstr_l_10(\IFID|plif_ifid.instr_l [10]),
	.plif_ifidinstr_l_9(\IFID|plif_ifid.instr_l [9]),
	.plif_ifidinstr_l_8(\IFID|plif_ifid.instr_l [8]),
	.plif_ifidinstr_l_7(\IFID|plif_ifid.instr_l [7]),
	.plif_ifidinstr_l_6(\IFID|plif_ifid.instr_l [6]),
	.instr_31(instr_31),
	.instr_29(instr_29),
	.instr_27(instr_27),
	.instr_26(instr_26),
	.instr_28(instr_28),
	.instr_30(instr_30),
	.instr_5(instr_5),
	.instr_1(instr_1),
	.instr_0(instr_0),
	.instr_2(instr_2),
	.instr_3(instr_3),
	.instr_4(instr_4),
	.instr_22(instr_22),
	.instr_21(instr_21),
	.instr_24(instr_24),
	.instr_23(instr_23),
	.instr_25(instr_25),
	.instr_17(instr_17),
	.instr_16(instr_16),
	.instr_19(instr_19),
	.instr_18(instr_18),
	.instr_20(instr_20),
	.instr_15(instr_15),
	.instr_14(instr_14),
	.instr_13(instr_13),
	.instr_12(instr_12),
	.instr_11(instr_11),
	.instr_10(instr_10),
	.instr_9(instr_9),
	.instr_8(instr_8),
	.instr_7(instr_7),
	.instr_6(instr_6),
	.plif_ifidrtnaddr_l_31(\IFID|plif_ifid.rtnaddr_l [31]),
	.plif_ifidrtnaddr_l_30(\IFID|plif_ifid.rtnaddr_l [30]),
	.plif_ifidrtnaddr_l_29(\IFID|plif_ifid.rtnaddr_l [29]),
	.plif_ifidrtnaddr_l_28(\IFID|plif_ifid.rtnaddr_l [28]),
	.plif_ifidrtnaddr_l_27(\IFID|plif_ifid.rtnaddr_l [27]),
	.plif_ifidrtnaddr_l_26(\IFID|plif_ifid.rtnaddr_l [26]),
	.plif_ifidrtnaddr_l_25(\IFID|plif_ifid.rtnaddr_l [25]),
	.plif_ifidrtnaddr_l_24(\IFID|plif_ifid.rtnaddr_l [24]),
	.plif_ifidrtnaddr_l_23(\IFID|plif_ifid.rtnaddr_l [23]),
	.plif_ifidrtnaddr_l_22(\IFID|plif_ifid.rtnaddr_l [22]),
	.plif_ifidrtnaddr_l_21(\IFID|plif_ifid.rtnaddr_l [21]),
	.plif_ifidrtnaddr_l_20(\IFID|plif_ifid.rtnaddr_l [20]),
	.plif_ifidrtnaddr_l_19(\IFID|plif_ifid.rtnaddr_l [19]),
	.plif_ifidrtnaddr_l_18(\IFID|plif_ifid.rtnaddr_l [18]),
	.plif_ifidrtnaddr_l_17(\IFID|plif_ifid.rtnaddr_l [17]),
	.plif_ifidrtnaddr_l_16(\IFID|plif_ifid.rtnaddr_l [16]),
	.plif_ifidrtnaddr_l_15(\IFID|plif_ifid.rtnaddr_l [15]),
	.plif_ifidrtnaddr_l_14(\IFID|plif_ifid.rtnaddr_l [14]),
	.plif_ifidrtnaddr_l_13(\IFID|plif_ifid.rtnaddr_l [13]),
	.plif_ifidrtnaddr_l_12(\IFID|plif_ifid.rtnaddr_l [12]),
	.plif_ifidrtnaddr_l_11(\IFID|plif_ifid.rtnaddr_l [11]),
	.plif_ifidrtnaddr_l_10(\IFID|plif_ifid.rtnaddr_l [10]),
	.plif_ifidrtnaddr_l_9(\IFID|plif_ifid.rtnaddr_l [9]),
	.plif_ifidrtnaddr_l_8(\IFID|plif_ifid.rtnaddr_l [8]),
	.plif_ifidrtnaddr_l_7(\IFID|plif_ifid.rtnaddr_l [7]),
	.plif_ifidrtnaddr_l_6(\IFID|plif_ifid.rtnaddr_l [6]),
	.plif_ifidrtnaddr_l_5(\IFID|plif_ifid.rtnaddr_l [5]),
	.plif_ifidrtnaddr_l_2(\IFID|plif_ifid.rtnaddr_l [2]),
	.plif_ifidrtnaddr_l_1(\IFID|plif_ifid.rtnaddr_l [1]),
	.plif_ifidrtnaddr_l_0(\IFID|plif_ifid.rtnaddr_l [0]),
	.plif_ifidrtnaddr_l_4(\IFID|plif_ifid.rtnaddr_l [4]),
	.plif_ifidrtnaddr_l_3(\IFID|plif_ifid.rtnaddr_l [3]),
	.ccifiwait_0(ccifiwait_0),
	.ifid_sRST(\HU|ifid_sRST~3_combout ),
	.CPUCLK(CLK),
	.nRST(nRST),
	.devpor(devpor),
	.devclrn(devclrn),
	.devoe(devoe));

pc PC(
	.PCreg_1(PCreg_1),
	.PCreg_0(PCreg_0),
	.pcifrtnaddr_2(\PC|pcif.rtnaddr[2]~0_combout ),
	.pcifrtnaddr_3(\PC|pcif.rtnaddr[3]~2_combout ),
	.pcifrtnaddr_4(\PC|pcif.rtnaddr[4]~4_combout ),
	.pcifrtnaddr_5(\PC|pcif.rtnaddr[5]~6_combout ),
	.pcifrtnaddr_6(\PC|pcif.rtnaddr[6]~8_combout ),
	.pcifrtnaddr_7(\PC|pcif.rtnaddr[7]~10_combout ),
	.pcifrtnaddr_8(\PC|pcif.rtnaddr[8]~12_combout ),
	.pcifrtnaddr_9(\PC|pcif.rtnaddr[9]~14_combout ),
	.pcifrtnaddr_10(\PC|pcif.rtnaddr[10]~16_combout ),
	.pcifrtnaddr_11(\PC|pcif.rtnaddr[11]~18_combout ),
	.pcifrtnaddr_12(\PC|pcif.rtnaddr[12]~20_combout ),
	.pcifrtnaddr_13(\PC|pcif.rtnaddr[13]~22_combout ),
	.pcifrtnaddr_14(\PC|pcif.rtnaddr[14]~24_combout ),
	.pcifrtnaddr_15(\PC|pcif.rtnaddr[15]~26_combout ),
	.pcifrtnaddr_16(\PC|pcif.rtnaddr[16]~28_combout ),
	.pcifrtnaddr_17(\PC|pcif.rtnaddr[17]~30_combout ),
	.pcifrtnaddr_18(\PC|pcif.rtnaddr[18]~32_combout ),
	.pcifrtnaddr_19(\PC|pcif.rtnaddr[19]~34_combout ),
	.pcifrtnaddr_20(\PC|pcif.rtnaddr[20]~36_combout ),
	.pcifrtnaddr_21(\PC|pcif.rtnaddr[21]~38_combout ),
	.pcifrtnaddr_22(\PC|pcif.rtnaddr[22]~40_combout ),
	.pcifrtnaddr_23(\PC|pcif.rtnaddr[23]~42_combout ),
	.pcifrtnaddr_24(\PC|pcif.rtnaddr[24]~44_combout ),
	.pcifrtnaddr_25(\PC|pcif.rtnaddr[25]~46_combout ),
	.pcifrtnaddr_26(\PC|pcif.rtnaddr[26]~48_combout ),
	.pcifrtnaddr_27(\PC|pcif.rtnaddr[27]~50_combout ),
	.pcifrtnaddr_28(\PC|pcif.rtnaddr[28]~52_combout ),
	.pcifrtnaddr_29(\PC|pcif.rtnaddr[29]~54_combout ),
	.pcifrtnaddr_30(\PC|pcif.rtnaddr[30]~56_combout ),
	.pcifrtnaddr_31(\PC|pcif.rtnaddr[31]~58_combout ),
	.PCreg_3(PCreg_3),
	.PCreg_2(PCreg_2),
	.PCreg_5(PCreg_5),
	.PCreg_4(PCreg_4),
	.PCreg_7(PCreg_7),
	.PCreg_6(PCreg_6),
	.PCreg_9(PCreg_9),
	.PCreg_8(PCreg_8),
	.PCreg_11(PCreg_11),
	.PCreg_10(PCreg_10),
	.PCreg_13(PCreg_13),
	.PCreg_12(PCreg_12),
	.PCreg_15(PCreg_15),
	.PCreg_14(PCreg_14),
	.PCreg_17(PCreg_17),
	.PCreg_16(PCreg_16),
	.PCreg_19(PCreg_19),
	.PCreg_18(PCreg_18),
	.PCreg_21(PCreg_21),
	.PCreg_20(PCreg_20),
	.PCreg_23(PCreg_23),
	.PCreg_22(PCreg_22),
	.PCreg_25(PCreg_25),
	.PCreg_24(PCreg_24),
	.PCreg_27(PCreg_27),
	.PCreg_26(PCreg_26),
	.PCreg_29(PCreg_29),
	.PCreg_28(PCreg_28),
	.PCreg_31(PCreg_31),
	.PCreg_30(PCreg_30),
	.plif_memwbpcsrc_l_1(\MEMWB|plif_memwb.pcsrc_l [1]),
	.always0(always0),
	.plif_memwbporto_l_31(\MEMWB|plif_memwb.porto_l [31]),
	.plif_memwbrtnaddr_l_31(\MEMWB|plif_memwb.rtnaddr_l [31]),
	.plif_memwbporto_l_30(\MEMWB|plif_memwb.porto_l [30]),
	.plif_memwbrtnaddr_l_30(\MEMWB|plif_memwb.rtnaddr_l [30]),
	.plif_memwbporto_l_29(\MEMWB|plif_memwb.porto_l [29]),
	.plif_memwbrtnaddr_l_29(\MEMWB|plif_memwb.rtnaddr_l [29]),
	.plif_memwbporto_l_28(\MEMWB|plif_memwb.porto_l [28]),
	.plif_memwbrtnaddr_l_28(\MEMWB|plif_memwb.rtnaddr_l [28]),
	.plif_memwbporto_l_27(\MEMWB|plif_memwb.porto_l [27]),
	.plif_memwbrtnaddr_l_27(\MEMWB|plif_memwb.rtnaddr_l [27]),
	.plif_memwbporto_l_26(\MEMWB|plif_memwb.porto_l [26]),
	.plif_memwbrtnaddr_l_26(\MEMWB|plif_memwb.rtnaddr_l [26]),
	.plif_memwbporto_l_25(\MEMWB|plif_memwb.porto_l [25]),
	.plif_memwbrtnaddr_l_25(\MEMWB|plif_memwb.rtnaddr_l [25]),
	.plif_memwbporto_l_24(\MEMWB|plif_memwb.porto_l [24]),
	.plif_memwbrtnaddr_l_24(\MEMWB|plif_memwb.rtnaddr_l [24]),
	.plif_memwbporto_l_23(\MEMWB|plif_memwb.porto_l [23]),
	.plif_memwbrtnaddr_l_23(\MEMWB|plif_memwb.rtnaddr_l [23]),
	.plif_memwbporto_l_22(\MEMWB|plif_memwb.porto_l [22]),
	.plif_memwbrtnaddr_l_22(\MEMWB|plif_memwb.rtnaddr_l [22]),
	.plif_memwbporto_l_21(\MEMWB|plif_memwb.porto_l [21]),
	.plif_memwbrtnaddr_l_21(\MEMWB|plif_memwb.rtnaddr_l [21]),
	.plif_memwbporto_l_20(\MEMWB|plif_memwb.porto_l [20]),
	.plif_memwbrtnaddr_l_20(\MEMWB|plif_memwb.rtnaddr_l [20]),
	.plif_memwbporto_l_19(\MEMWB|plif_memwb.porto_l [19]),
	.plif_memwbrtnaddr_l_19(\MEMWB|plif_memwb.rtnaddr_l [19]),
	.plif_memwbporto_l_18(\MEMWB|plif_memwb.porto_l [18]),
	.plif_memwbrtnaddr_l_18(\MEMWB|plif_memwb.rtnaddr_l [18]),
	.plif_memwbporto_l_17(\MEMWB|plif_memwb.porto_l [17]),
	.plif_memwbrtnaddr_l_17(\MEMWB|plif_memwb.rtnaddr_l [17]),
	.plif_memwbporto_l_16(\MEMWB|plif_memwb.porto_l [16]),
	.plif_memwbrtnaddr_l_16(\MEMWB|plif_memwb.rtnaddr_l [16]),
	.plif_memwbporto_l_15(\MEMWB|plif_memwb.porto_l [15]),
	.plif_memwbrtnaddr_l_15(\MEMWB|plif_memwb.rtnaddr_l [15]),
	.plif_memwbporto_l_14(\MEMWB|plif_memwb.porto_l [14]),
	.plif_memwbrtnaddr_l_14(\MEMWB|plif_memwb.rtnaddr_l [14]),
	.plif_memwbporto_l_13(\MEMWB|plif_memwb.porto_l [13]),
	.plif_memwbrtnaddr_l_13(\MEMWB|plif_memwb.rtnaddr_l [13]),
	.plif_memwbporto_l_12(\MEMWB|plif_memwb.porto_l [12]),
	.plif_memwbrtnaddr_l_12(\MEMWB|plif_memwb.rtnaddr_l [12]),
	.plif_memwbporto_l_11(\MEMWB|plif_memwb.porto_l [11]),
	.plif_memwbrtnaddr_l_11(\MEMWB|plif_memwb.rtnaddr_l [11]),
	.plif_memwbporto_l_10(\MEMWB|plif_memwb.porto_l [10]),
	.plif_memwbrtnaddr_l_10(\MEMWB|plif_memwb.rtnaddr_l [10]),
	.plif_memwbporto_l_9(\MEMWB|plif_memwb.porto_l [9]),
	.plif_memwbrtnaddr_l_9(\MEMWB|plif_memwb.rtnaddr_l [9]),
	.plif_memwbporto_l_8(\MEMWB|plif_memwb.porto_l [8]),
	.plif_memwbrtnaddr_l_8(\MEMWB|plif_memwb.rtnaddr_l [8]),
	.plif_memwbporto_l_7(\MEMWB|plif_memwb.porto_l [7]),
	.plif_memwbrtnaddr_l_7(\MEMWB|plif_memwb.rtnaddr_l [7]),
	.plif_memwbporto_l_6(\MEMWB|plif_memwb.porto_l [6]),
	.plif_memwbrtnaddr_l_6(\MEMWB|plif_memwb.rtnaddr_l [6]),
	.plif_memwbporto_l_5(\MEMWB|plif_memwb.porto_l [5]),
	.plif_memwbrtnaddr_l_5(\MEMWB|plif_memwb.rtnaddr_l [5]),
	.plif_memwbporto_l_2(\MEMWB|plif_memwb.porto_l [2]),
	.plif_memwbrtnaddr_l_2(\MEMWB|plif_memwb.rtnaddr_l [2]),
	.plif_memwbporto_l_1(\MEMWB|plif_memwb.porto_l [1]),
	.plif_memwbrtnaddr_l_1(\MEMWB|plif_memwb.rtnaddr_l [1]),
	.plif_memwbporto_l_0(\MEMWB|plif_memwb.porto_l [0]),
	.plif_memwbrtnaddr_l_0(\MEMWB|plif_memwb.rtnaddr_l [0]),
	.plif_memwbporto_l_4(\MEMWB|plif_memwb.porto_l [4]),
	.plif_memwbrtnaddr_l_4(\MEMWB|plif_memwb.rtnaddr_l [4]),
	.plif_memwbporto_l_3(\MEMWB|plif_memwb.porto_l [3]),
	.plif_memwbrtnaddr_l_3(\MEMWB|plif_memwb.rtnaddr_l [3]),
	.pcsrc(\pcsrc~0_combout ),
	.ifid_en(\HU|ifid_en~0_combout ),
	.plif_memwbjaddr_l_1(\MEMWB|plif_memwb.jaddr_l [1]),
	.plif_memwbextimm_l_1(\MEMWB|plif_memwb.extimm_l [1]),
	.plif_memwbextimm_l_0(\MEMWB|plif_memwb.extimm_l [0]),
	.\pcif.rambusy (\HU|rambusy~0_combout ),
	.plif_memwbjaddr_l_0(\MEMWB|plif_memwb.jaddr_l [0]),
	.plif_memwbjaddr_l_3(\MEMWB|plif_memwb.jaddr_l [3]),
	.plif_memwbextimm_l_3(\MEMWB|plif_memwb.extimm_l [3]),
	.plif_memwbextimm_l_2(\MEMWB|plif_memwb.extimm_l [2]),
	.plif_memwbjaddr_l_2(\MEMWB|plif_memwb.jaddr_l [2]),
	.plif_memwbjaddr_l_5(\MEMWB|plif_memwb.jaddr_l [5]),
	.plif_memwbextimm_l_5(\MEMWB|plif_memwb.extimm_l [5]),
	.plif_memwbextimm_l_4(\MEMWB|plif_memwb.extimm_l [4]),
	.plif_memwbjaddr_l_4(\MEMWB|plif_memwb.jaddr_l [4]),
	.plif_memwbjaddr_l_7(\MEMWB|plif_memwb.jaddr_l [7]),
	.plif_memwbextimm_l_7(\MEMWB|plif_memwb.extimm_l [7]),
	.plif_memwbextimm_l_6(\MEMWB|plif_memwb.extimm_l [6]),
	.plif_memwbjaddr_l_6(\MEMWB|plif_memwb.jaddr_l [6]),
	.plif_memwbjaddr_l_9(\MEMWB|plif_memwb.jaddr_l [9]),
	.plif_memwbextimm_l_9(\MEMWB|plif_memwb.extimm_l [9]),
	.plif_memwbextimm_l_8(\MEMWB|plif_memwb.extimm_l [8]),
	.plif_memwbjaddr_l_8(\MEMWB|plif_memwb.jaddr_l [8]),
	.plif_memwbjaddr_l_11(\MEMWB|plif_memwb.jaddr_l [11]),
	.plif_memwbextimm_l_11(\MEMWB|plif_memwb.extimm_l [11]),
	.plif_memwbextimm_l_10(\MEMWB|plif_memwb.extimm_l [10]),
	.plif_memwbjaddr_l_10(\MEMWB|plif_memwb.jaddr_l [10]),
	.plif_memwbjaddr_l_13(\MEMWB|plif_memwb.jaddr_l [13]),
	.plif_memwbextimm_l_13(\MEMWB|plif_memwb.extimm_l [13]),
	.plif_memwbextimm_l_12(\MEMWB|plif_memwb.extimm_l [12]),
	.plif_memwbjaddr_l_12(\MEMWB|plif_memwb.jaddr_l [12]),
	.plif_memwbjaddr_l_15(\MEMWB|plif_memwb.jaddr_l [15]),
	.plif_memwbextimm_l_15(\MEMWB|plif_memwb.extimm_l [15]),
	.plif_memwbextimm_l_14(\MEMWB|plif_memwb.extimm_l [14]),
	.plif_memwbjaddr_l_14(\MEMWB|plif_memwb.jaddr_l [14]),
	.plif_memwbjaddr_l_17(\MEMWB|plif_memwb.jaddr_l [17]),
	.plif_memwbextimm_l_17(\MEMWB|plif_memwb.extimm_l [17]),
	.plif_memwbextimm_l_16(\MEMWB|plif_memwb.extimm_l [16]),
	.plif_memwbjaddr_l_16(\MEMWB|plif_memwb.jaddr_l [16]),
	.plif_memwbjaddr_l_19(\MEMWB|plif_memwb.jaddr_l [19]),
	.plif_memwbextimm_l_19(\MEMWB|plif_memwb.extimm_l [19]),
	.plif_memwbextimm_l_18(\MEMWB|plif_memwb.extimm_l [18]),
	.plif_memwbjaddr_l_18(\MEMWB|plif_memwb.jaddr_l [18]),
	.plif_memwbjaddr_l_21(\MEMWB|plif_memwb.jaddr_l [21]),
	.plif_memwbextimm_l_21(\MEMWB|plif_memwb.extimm_l [21]),
	.plif_memwbextimm_l_20(\MEMWB|plif_memwb.extimm_l [20]),
	.plif_memwbjaddr_l_20(\MEMWB|plif_memwb.jaddr_l [20]),
	.plif_memwbjaddr_l_23(\MEMWB|plif_memwb.jaddr_l [23]),
	.plif_memwbextimm_l_23(\MEMWB|plif_memwb.extimm_l [23]),
	.plif_memwbextimm_l_22(\MEMWB|plif_memwb.extimm_l [22]),
	.plif_memwbjaddr_l_22(\MEMWB|plif_memwb.jaddr_l [22]),
	.plif_memwbjaddr_l_25(\MEMWB|plif_memwb.jaddr_l [25]),
	.plif_memwbextimm_l_25(\MEMWB|plif_memwb.extimm_l [25]),
	.plif_memwbextimm_l_24(\MEMWB|plif_memwb.extimm_l [24]),
	.plif_memwbjaddr_l_24(\MEMWB|plif_memwb.jaddr_l [24]),
	.plif_memwbextimm_l_27(\MEMWB|plif_memwb.extimm_l [27]),
	.plif_memwbextimm_l_26(\MEMWB|plif_memwb.extimm_l [26]),
	.plif_memwbextimm_l_29(\MEMWB|plif_memwb.extimm_l [29]),
	.plif_memwbextimm_l_28(\MEMWB|plif_memwb.extimm_l [28]),
	.CLK(CLK),
	.nRST(nRST),
	.devpor(devpor),
	.devclrn(devclrn),
	.devoe(devoe));

alu ALU(
	.plif_idexaluop_l_3(\IDEX|plif_idex.aluop_l [3]),
	.plif_idexaluop_l_2(\IDEX|plif_idex.aluop_l [2]),
	.plif_idexaluop_l_1(\IDEX|plif_idex.aluop_l [1]),
	.plif_idexaluop_l_0(\IDEX|plif_idex.aluop_l [0]),
	.portb(\portb~4_combout ),
	.portb1(\portb~6_combout ),
	.portb2(\portb~8_combout ),
	.portb3(\portb~10_combout ),
	.portb4(\portb~12_combout ),
	.portb5(\portb~14_combout ),
	.portb6(\portb~16_combout ),
	.portb7(\portb~18_combout ),
	.portb8(\portb~20_combout ),
	.portb9(\portb~22_combout ),
	.portb10(\portb~24_combout ),
	.portb11(\portb~26_combout ),
	.portb12(\portb~28_combout ),
	.portb13(\portb~30_combout ),
	.portb14(\portb~32_combout ),
	.portb15(\portb~34_combout ),
	.portb16(\portb~36_combout ),
	.portb17(\portb~38_combout ),
	.portb18(\portb~40_combout ),
	.portb19(\portb~42_combout ),
	.portb20(\portb~44_combout ),
	.portb21(\portb~46_combout ),
	.portb22(\portb~48_combout ),
	.portb23(\portb~50_combout ),
	.portb24(\portb~52_combout ),
	.portb25(\portb~54_combout ),
	.portb26(\portb~56_combout ),
	.porta(\porta~55_combout ),
	.porta1(\porta~57_combout ),
	.portb27(\portb~58_combout ),
	.portb28(\portb~60_combout ),
	.porta2(\porta~59_combout ),
	.porta3(\porta~61_combout ),
	.portb29(\portb~62_combout ),
	.porta4(\porta~63_combout ),
	.portb30(\portb~64_combout ),
	.portb31(\portb~66_combout ),
	.porta5(\porta~76_combout ),
	.plif_idexrdat1_l_29(\IDEX|plif_idex.rdat1_l [29]),
	.porta6(\porta~81_combout ),
	.plif_idexrdat1_l_25(\IDEX|plif_idex.rdat1_l [25]),
	.porta7(\porta~91_combout ),
	.Selector30(\ALU|Selector30~8_combout ),
	.Selector31(\ALU|Selector31~8_combout ),
	.Selector28(\ALU|Selector28~10_combout ),
	.Selector29(\ALU|Selector29~8_combout ),
	.Selector26(\ALU|Selector26~8_combout ),
	.Selector27(\ALU|Selector27~8_combout ),
	.Selector24(\ALU|Selector24~9_combout ),
	.Selector25(\ALU|Selector25~7_combout ),
	.Selector22(\ALU|Selector22~8_combout ),
	.Selector23(\ALU|Selector23~9_combout ),
	.Selector20(\ALU|Selector20~9_combout ),
	.Selector21(\ALU|Selector21~8_combout ),
	.Selector18(\ALU|Selector18~9_combout ),
	.Selector19(\ALU|Selector19~8_combout ),
	.Selector16(\ALU|Selector16~10_combout ),
	.Selector17(\ALU|Selector17~7_combout ),
	.Selector14(\ALU|Selector14~8_combout ),
	.Selector15(\ALU|Selector15~8_combout ),
	.Selector12(\ALU|Selector12~10_combout ),
	.Selector13(\ALU|Selector13~8_combout ),
	.Selector10(\ALU|Selector10~8_combout ),
	.Selector11(\ALU|Selector11~9_combout ),
	.Selector8(\ALU|Selector8~10_combout ),
	.Selector9(\ALU|Selector9~8_combout ),
	.Selector6(\ALU|Selector6~8_combout ),
	.Selector7(\ALU|Selector7~11_combout ),
	.Selector4(\ALU|Selector4~10_combout ),
	.Selector5(\ALU|Selector5~8_combout ),
	.Selector2(\ALU|Selector2~11_combout ),
	.Selector3(\ALU|Selector3~11_combout ),
	.Selector0(\ALU|Selector0~34_combout ),
	.Selector1(\ALU|Selector1~20_combout ),
	.WideOr11(\ALU|WideOr1~combout ),
	.porta8(\porta~92_combout ),
	.porta9(\porta~93_combout ),
	.porta10(\porta~94_combout ),
	.porta11(\porta~95_combout ),
	.porta12(\porta~96_combout ),
	.porta13(\porta~97_combout ),
	.porta14(\porta~98_combout ),
	.porta15(\porta~99_combout ),
	.porta16(\porta~100_combout ),
	.porta17(\porta~101_combout ),
	.porta18(\porta~102_combout ),
	.porta19(\porta~103_combout ),
	.porta20(\porta~104_combout ),
	.porta21(\porta~105_combout ),
	.porta22(\porta~106_combout ),
	.porta23(\porta~107_combout ),
	.porta24(\porta~108_combout ),
	.porta25(\porta~109_combout ),
	.porta26(\porta~110_combout ),
	.porta27(\porta~111_combout ),
	.porta28(\porta~112_combout ),
	.porta29(\porta~113_combout ),
	.porta30(\porta~114_combout ),
	.porta31(\porta~115_combout ),
	.porta32(\porta~116_combout ),
	.porta33(\porta~117_combout ),
	.porta34(\porta~118_combout ),
	.devpor(devpor),
	.devclrn(devclrn),
	.devoe(devoe));

forwarding_unit FU(
	.plif_exmemregen_l(\EXMEM|plif_exmem.regen_l~q ),
	.plif_exmemwsel_l_0(\EXMEM|plif_exmem.wsel_l [0]),
	.plif_exmemwsel_l_1(\EXMEM|plif_exmem.wsel_l [1]),
	.plif_idexrsel2_l_1(\IDEX|plif_idex.rsel2_l [1]),
	.plif_idexrsel2_l_0(\IDEX|plif_idex.rsel2_l [0]),
	.plif_exmemwsel_l_4(\EXMEM|plif_exmem.wsel_l [4]),
	.plif_exmemwsel_l_3(\EXMEM|plif_exmem.wsel_l [3]),
	.plif_exmemwsel_l_2(\EXMEM|plif_exmem.wsel_l [2]),
	.always0(\FU|always0~2_combout ),
	.plif_idexrsel2_l_2(\IDEX|plif_idex.rsel2_l [2]),
	.plif_idexrsel2_l_3(\IDEX|plif_idex.rsel2_l [3]),
	.always01(\FU|always0~3_combout ),
	.plif_idexrsel2_l_4(\IDEX|plif_idex.rsel2_l [4]),
	.always02(\FU|always0~4_combout ),
	.plif_memwbwsel_l_4(\MEMWB|plif_memwb.wsel_l [4]),
	.plif_memwbwsel_l_3(\MEMWB|plif_memwb.wsel_l [3]),
	.plif_memwbwsel_l_0(\MEMWB|plif_memwb.wsel_l [0]),
	.plif_memwbwsel_l_2(\MEMWB|plif_memwb.wsel_l [2]),
	.plif_memwbwsel_l_1(\MEMWB|plif_memwb.wsel_l [1]),
	.Decoder0(\RF|Decoder0~20_combout ),
	.WideOr01(\FU|WideOr0~combout ),
	.fwdc(\FU|fwdc~2_combout ),
	.plif_memwbregen_l(\MEMWB|plif_memwb.regen_l~q ),
	.plif_idexrsel1_l_4(\IDEX|plif_idex.rsel1_l [4]),
	.plif_idexrsel1_l_1(\IDEX|plif_idex.rsel1_l [1]),
	.plif_idexrsel1_l_0(\IDEX|plif_idex.rsel1_l [0]),
	.plif_idexrsel1_l_2(\IDEX|plif_idex.rsel1_l [2]),
	.plif_idexrsel1_l_3(\IDEX|plif_idex.rsel1_l [3]),
	.fwda(\FU|fwda~3_combout ),
	.always03(\FU|always0~8_combout ),
	.devpor(devpor),
	.devclrn(devclrn),
	.devoe(devoe));

hazard_unit HU(
	.always1(always1),
	.plif_memwbpcsrc_l_1(\MEMWB|plif_memwb.pcsrc_l [1]),
	.plif_memwbpcsrc_l_0(\MEMWB|plif_memwb.pcsrc_l [0]),
	.always0(always0),
	.plif_idexpcsrc_l_1(\IDEX|plif_idex.pcsrc_l [1]),
	.plif_idexpcsrc_l_0(\IDEX|plif_idex.pcsrc_l [0]),
	.plif_exmempcsrc_l_1(\EXMEM|plif_exmem.pcsrc_l [1]),
	.plif_exmempcsrc_l_0(\EXMEM|plif_exmem.pcsrc_l [0]),
	.ifid_sRST(\HU|ifid_sRST~2_combout ),
	.exmem_en(\HU|exmem_en~0_combout ),
	.pcsrc(\pcsrc~0_combout ),
	.plif_idexdmemREN_l(\IDEX|plif_idex.dmemREN_l~q ),
	.plif_idexwsel_l_0(\IDEX|plif_idex.wsel_l [0]),
	.plif_idexwsel_l_1(\IDEX|plif_idex.wsel_l [1]),
	.Selector4(\CU|Selector4~1_combout ),
	.Selector5(\CU|Selector5~1_combout ),
	.plif_idexwsel_l_2(\IDEX|plif_idex.wsel_l [2]),
	.plif_idexwsel_l_3(\IDEX|plif_idex.wsel_l [3]),
	.Selector2(\CU|Selector2~0_combout ),
	.Selector3(\CU|Selector3~0_combout ),
	.plif_idexwsel_l_4(\IDEX|plif_idex.wsel_l [4]),
	.Selector1(\CU|Selector1~0_combout ),
	.Selector9(\CU|Selector9~1_combout ),
	.Selector10(\CU|Selector10~0_combout ),
	.Selector7(\CU|Selector7~0_combout ),
	.Selector8(\CU|Selector8~0_combout ),
	.Selector6(\CU|Selector6~0_combout ),
	.ifid_en(\HU|ifid_en~0_combout ),
	.rambusy(\HU|rambusy~0_combout ),
	.idex_sRST(\HU|idex_sRST~3_combout ),
	.idex_sRST1(\HU|idex_sRST~4_combout ),
	.idex_sRST2(\HU|idex_sRST~5_combout ),
	.ifid_sRST1(\HU|ifid_sRST~3_combout ),
	.devpor(devpor),
	.devclrn(devclrn),
	.devoe(devoe));

control_unit CU(
	.plif_ifidinstr_l_31(\IFID|plif_ifid.instr_l [31]),
	.plif_ifidinstr_l_29(\IFID|plif_ifid.instr_l [29]),
	.plif_ifidinstr_l_27(\IFID|plif_ifid.instr_l [27]),
	.plif_ifidinstr_l_26(\IFID|plif_ifid.instr_l [26]),
	.plif_ifidinstr_l_28(\IFID|plif_ifid.instr_l [28]),
	.Equal16(\CU|Equal16~0_combout ),
	.plif_ifidinstr_l_30(\IFID|plif_ifid.instr_l [30]),
	.Equal22(\CU|Equal22~0_combout ),
	.plif_ifidinstr_l_5(\IFID|plif_ifid.instr_l [5]),
	.plif_ifidinstr_l_1(\IFID|plif_ifid.instr_l [1]),
	.plif_ifidinstr_l_0(\IFID|plif_ifid.instr_l [0]),
	.plif_ifidinstr_l_2(\IFID|plif_ifid.instr_l [2]),
	.plif_ifidinstr_l_3(\IFID|plif_ifid.instr_l [3]),
	.WideNor0(\CU|WideNor0~2_combout ),
	.Equal11(\CU|Equal11~0_combout ),
	.Equal26(\CU|Equal26~0_combout ),
	.plif_ifidinstr_l_4(\IFID|plif_ifid.instr_l [4]),
	.Equal21(\CU|Equal21~0_combout ),
	.WideOr141(\CU|WideOr14~0_combout ),
	.Equal13(\CU|Equal13~1_combout ),
	.aluop_l(\IDEX|aluop_l~0_combout ),
	.WideNor1(\CU|WideNor1~0_combout ),
	.Selector22(\CU|Selector22~6_combout ),
	.Selector4(\CU|Selector4~0_combout ),
	.plif_ifidinstr_l_22(\IFID|plif_ifid.instr_l [22]),
	.Selector41(\CU|Selector4~1_combout ),
	.plif_ifidinstr_l_21(\IFID|plif_ifid.instr_l [21]),
	.Selector5(\CU|Selector5~1_combout ),
	.plif_ifidinstr_l_24(\IFID|plif_ifid.instr_l [24]),
	.Selector2(\CU|Selector2~0_combout ),
	.plif_ifidinstr_l_23(\IFID|plif_ifid.instr_l [23]),
	.Selector3(\CU|Selector3~0_combout ),
	.plif_ifidinstr_l_25(\IFID|plif_ifid.instr_l [25]),
	.Selector1(\CU|Selector1~0_combout ),
	.Equal6(\CU|Equal6~0_combout ),
	.Selector11(\CU|Selector11~0_combout ),
	.Selector21(\CU|Selector21~0_combout ),
	.Selector9(\CU|Selector9~0_combout ),
	.plif_ifidinstr_l_17(\IFID|plif_ifid.instr_l [17]),
	.Selector91(\CU|Selector9~1_combout ),
	.plif_ifidinstr_l_16(\IFID|plif_ifid.instr_l [16]),
	.Selector10(\CU|Selector10~0_combout ),
	.plif_ifidinstr_l_19(\IFID|plif_ifid.instr_l [19]),
	.Selector7(\CU|Selector7~0_combout ),
	.plif_ifidinstr_l_18(\IFID|plif_ifid.instr_l [18]),
	.Selector8(\CU|Selector8~0_combout ),
	.plif_ifidinstr_l_20(\IFID|plif_ifid.instr_l [20]),
	.Selector6(\CU|Selector6~0_combout ),
	.Equal23(\CU|Equal23~0_combout ),
	.pcsrc(\CU|pcsrc~0_combout ),
	.Equal1(\CU|Equal1~0_combout ),
	.Equal20(\CU|Equal20~0_combout ),
	.WideNor11(\CU|WideNor1~1_combout ),
	.Equal19(\CU|Equal19~0_combout ),
	.Equal12(\CU|Equal1~1_combout ),
	.Equal18(\CU|Equal18~0_combout ),
	.Selector221(\CU|Selector22~7_combout ),
	.WideOr142(\CU|WideOr14~combout ),
	.WideOr151(\CU|WideOr15~combout ),
	.WideOr161(\CU|WideOr16~0_combout ),
	.plif_ifidinstr_l_10(\IFID|plif_ifid.instr_l [10]),
	.plif_ifidinstr_l_9(\IFID|plif_ifid.instr_l [9]),
	.plif_ifidinstr_l_8(\IFID|plif_ifid.instr_l [8]),
	.plif_ifidinstr_l_7(\IFID|plif_ifid.instr_l [7]),
	.plif_ifidinstr_l_6(\IFID|plif_ifid.instr_l [6]),
	.Selector14(\CU|Selector14~0_combout ),
	.Selector15(\CU|Selector15~0_combout ),
	.Selector16(\CU|Selector16~0_combout ),
	.Selector17(\CU|Selector17~0_combout ),
	.Selector18(\CU|Selector18~0_combout ),
	.Selector24(\CU|Selector24~0_combout ),
	.Equal121(\CU|Equal12~0_combout ),
	.Selector0(\CU|Selector0~2_combout ),
	.Equal25(\CU|Equal25~4_combout ),
	.devpor(devpor),
	.devclrn(devclrn),
	.devoe(devoe));

register_file RF(
	.plif_memwbregsrc_l_1(\MEMWB|plif_memwb.regsrc_l [1]),
	.wdat_31(\wdat[31]~0_combout ),
	.plif_memwbrtnaddr_l_31(\MEMWB|plif_memwb.rtnaddr_l [31]),
	.plif_memwbwsel_l_4(\MEMWB|plif_memwb.wsel_l [4]),
	.plif_memwbwsel_l_3(\MEMWB|plif_memwb.wsel_l [3]),
	.plif_memwbwsel_l_0(\MEMWB|plif_memwb.wsel_l [0]),
	.plif_memwbwsel_l_2(\MEMWB|plif_memwb.wsel_l [2]),
	.plif_memwbwsel_l_1(\MEMWB|plif_memwb.wsel_l [1]),
	.Decoder0(\RF|Decoder0~20_combout ),
	.WideOr0(\FU|WideOr0~combout ),
	.plif_memwbregen_l(\MEMWB|plif_memwb.regen_l~q ),
	.wdat_30(\wdat[30]~2_combout ),
	.plif_memwbrtnaddr_l_30(\MEMWB|plif_memwb.rtnaddr_l [30]),
	.wdat_29(\wdat[29]~4_combout ),
	.plif_memwbrtnaddr_l_29(\MEMWB|plif_memwb.rtnaddr_l [29]),
	.wdat_28(\wdat[28]~6_combout ),
	.plif_memwbrtnaddr_l_28(\MEMWB|plif_memwb.rtnaddr_l [28]),
	.wdat_27(\wdat[27]~8_combout ),
	.plif_memwbrtnaddr_l_27(\MEMWB|plif_memwb.rtnaddr_l [27]),
	.wdat_26(\wdat[26]~10_combout ),
	.plif_memwbrtnaddr_l_26(\MEMWB|plif_memwb.rtnaddr_l [26]),
	.wdat_25(\wdat[25]~12_combout ),
	.plif_memwbrtnaddr_l_25(\MEMWB|plif_memwb.rtnaddr_l [25]),
	.wdat_24(\wdat[24]~14_combout ),
	.plif_memwbrtnaddr_l_24(\MEMWB|plif_memwb.rtnaddr_l [24]),
	.wdat_23(\wdat[23]~16_combout ),
	.plif_memwbrtnaddr_l_23(\MEMWB|plif_memwb.rtnaddr_l [23]),
	.wdat_22(\wdat[22]~18_combout ),
	.plif_memwbrtnaddr_l_22(\MEMWB|plif_memwb.rtnaddr_l [22]),
	.wdat_21(\wdat[21]~20_combout ),
	.plif_memwbrtnaddr_l_21(\MEMWB|plif_memwb.rtnaddr_l [21]),
	.wdat_20(\wdat[20]~22_combout ),
	.plif_memwbrtnaddr_l_20(\MEMWB|plif_memwb.rtnaddr_l [20]),
	.wdat_19(\wdat[19]~24_combout ),
	.plif_memwbrtnaddr_l_19(\MEMWB|plif_memwb.rtnaddr_l [19]),
	.wdat_18(\wdat[18]~26_combout ),
	.plif_memwbrtnaddr_l_18(\MEMWB|plif_memwb.rtnaddr_l [18]),
	.wdat_17(\wdat[17]~28_combout ),
	.plif_memwbrtnaddr_l_17(\MEMWB|plif_memwb.rtnaddr_l [17]),
	.wdat_16(\wdat[16]~30_combout ),
	.plif_memwbrtnaddr_l_16(\MEMWB|plif_memwb.rtnaddr_l [16]),
	.wdat_15(\wdat[15]~32_combout ),
	.plif_memwbrtnaddr_l_15(\MEMWB|plif_memwb.rtnaddr_l [15]),
	.wdat_14(\wdat[14]~34_combout ),
	.plif_memwbrtnaddr_l_14(\MEMWB|plif_memwb.rtnaddr_l [14]),
	.wdat_13(\wdat[13]~36_combout ),
	.plif_memwbrtnaddr_l_13(\MEMWB|plif_memwb.rtnaddr_l [13]),
	.wdat_12(\wdat[12]~38_combout ),
	.plif_memwbrtnaddr_l_12(\MEMWB|plif_memwb.rtnaddr_l [12]),
	.wdat_11(\wdat[11]~40_combout ),
	.plif_memwbrtnaddr_l_11(\MEMWB|plif_memwb.rtnaddr_l [11]),
	.wdat_10(\wdat[10]~42_combout ),
	.plif_memwbrtnaddr_l_10(\MEMWB|plif_memwb.rtnaddr_l [10]),
	.wdat_9(\wdat[9]~44_combout ),
	.plif_memwbrtnaddr_l_9(\MEMWB|plif_memwb.rtnaddr_l [9]),
	.wdat_8(\wdat[8]~46_combout ),
	.plif_memwbrtnaddr_l_8(\MEMWB|plif_memwb.rtnaddr_l [8]),
	.wdat_7(\wdat[7]~48_combout ),
	.plif_memwbrtnaddr_l_7(\MEMWB|plif_memwb.rtnaddr_l [7]),
	.wdat_6(\wdat[6]~50_combout ),
	.plif_memwbrtnaddr_l_6(\MEMWB|plif_memwb.rtnaddr_l [6]),
	.wdat_5(\wdat[5]~52_combout ),
	.plif_memwbrtnaddr_l_5(\MEMWB|plif_memwb.rtnaddr_l [5]),
	.wdat_2(\wdat[2]~54_combout ),
	.plif_memwbrtnaddr_l_2(\MEMWB|plif_memwb.rtnaddr_l [2]),
	.wdat_1(\wdat[1]~56_combout ),
	.plif_memwbrtnaddr_l_1(\MEMWB|plif_memwb.rtnaddr_l [1]),
	.wdat_0(\wdat[0]~58_combout ),
	.plif_memwbrtnaddr_l_0(\MEMWB|plif_memwb.rtnaddr_l [0]),
	.wdat_4(\wdat[4]~60_combout ),
	.plif_memwbrtnaddr_l_4(\MEMWB|plif_memwb.rtnaddr_l [4]),
	.wdat_3(\wdat[3]~62_combout ),
	.plif_memwbrtnaddr_l_3(\MEMWB|plif_memwb.rtnaddr_l [3]),
	.Selector4(\CU|Selector4~0_combout ),
	.plif_ifidinstr_l_22(\IFID|plif_ifid.instr_l [22]),
	.Selector41(\CU|Selector4~1_combout ),
	.Selector5(\CU|Selector5~1_combout ),
	.Selector2(\CU|Selector2~0_combout ),
	.Selector3(\CU|Selector3~0_combout ),
	.Selector9(\CU|Selector9~0_combout ),
	.plif_ifidinstr_l_17(\IFID|plif_ifid.instr_l [17]),
	.Selector91(\CU|Selector9~1_combout ),
	.Selector10(\CU|Selector10~0_combout ),
	.Selector7(\CU|Selector7~0_combout ),
	.Selector8(\CU|Selector8~0_combout ),
	.Mux32(\RF|Mux32~9_combout ),
	.Mux321(\RF|Mux32~19_combout ),
	.Mux33(\RF|Mux33~9_combout ),
	.Mux331(\RF|Mux33~19_combout ),
	.Mux34(\RF|Mux34~9_combout ),
	.Mux341(\RF|Mux34~19_combout ),
	.Mux35(\RF|Mux35~9_combout ),
	.Mux351(\RF|Mux35~19_combout ),
	.Mux36(\RF|Mux36~9_combout ),
	.Mux361(\RF|Mux36~19_combout ),
	.Mux37(\RF|Mux37~9_combout ),
	.Mux371(\RF|Mux37~19_combout ),
	.Mux38(\RF|Mux38~9_combout ),
	.Mux381(\RF|Mux38~19_combout ),
	.Mux39(\RF|Mux39~9_combout ),
	.Mux391(\RF|Mux39~19_combout ),
	.Mux40(\RF|Mux40~9_combout ),
	.Mux401(\RF|Mux40~19_combout ),
	.Mux41(\RF|Mux41~9_combout ),
	.Mux411(\RF|Mux41~19_combout ),
	.Mux42(\RF|Mux42~9_combout ),
	.Mux421(\RF|Mux42~19_combout ),
	.Mux43(\RF|Mux43~9_combout ),
	.Mux431(\RF|Mux43~19_combout ),
	.Mux44(\RF|Mux44~9_combout ),
	.Mux441(\RF|Mux44~19_combout ),
	.Mux45(\RF|Mux45~9_combout ),
	.Mux451(\RF|Mux45~19_combout ),
	.Mux46(\RF|Mux46~9_combout ),
	.Mux461(\RF|Mux46~19_combout ),
	.Mux47(\RF|Mux47~9_combout ),
	.Mux471(\RF|Mux47~19_combout ),
	.Mux48(\RF|Mux48~9_combout ),
	.Mux481(\RF|Mux48~19_combout ),
	.Mux49(\RF|Mux49~9_combout ),
	.Mux491(\RF|Mux49~19_combout ),
	.Mux50(\RF|Mux50~9_combout ),
	.Mux501(\RF|Mux50~19_combout ),
	.Mux51(\RF|Mux51~9_combout ),
	.Mux511(\RF|Mux51~19_combout ),
	.Mux52(\RF|Mux52~9_combout ),
	.Mux521(\RF|Mux52~19_combout ),
	.Mux53(\RF|Mux53~9_combout ),
	.Mux531(\RF|Mux53~19_combout ),
	.Mux54(\RF|Mux54~9_combout ),
	.Mux541(\RF|Mux54~19_combout ),
	.Mux55(\RF|Mux55~9_combout ),
	.Mux551(\RF|Mux55~19_combout ),
	.Mux56(\RF|Mux56~9_combout ),
	.Mux561(\RF|Mux56~19_combout ),
	.Mux57(\RF|Mux57~9_combout ),
	.Mux571(\RF|Mux57~19_combout ),
	.Mux58(\RF|Mux58~9_combout ),
	.Mux581(\RF|Mux58~19_combout ),
	.Mux29(\RF|Mux29~9_combout ),
	.Mux291(\RF|Mux29~19_combout ),
	.Mux30(\RF|Mux30~9_combout ),
	.Mux301(\RF|Mux30~19_combout ),
	.Mux63(\RF|Mux63~9_combout ),
	.Mux631(\RF|Mux63~19_combout ),
	.Mux62(\RF|Mux62~9_combout ),
	.Mux621(\RF|Mux62~19_combout ),
	.Mux27(\RF|Mux27~9_combout ),
	.Mux271(\RF|Mux27~19_combout ),
	.Mux28(\RF|Mux28~9_combout ),
	.Mux281(\RF|Mux28~19_combout ),
	.Mux61(\RF|Mux61~9_combout ),
	.Mux611(\RF|Mux61~19_combout ),
	.Mux23(\RF|Mux23~9_combout ),
	.Mux231(\RF|Mux23~19_combout ),
	.Mux24(\RF|Mux24~9_combout ),
	.Mux241(\RF|Mux24~19_combout ),
	.Mux25(\RF|Mux25~9_combout ),
	.Mux251(\RF|Mux25~19_combout ),
	.Mux26(\RF|Mux26~9_combout ),
	.Mux261(\RF|Mux26~19_combout ),
	.Mux60(\RF|Mux60~9_combout ),
	.Mux601(\RF|Mux60~19_combout ),
	.Mux15(\RF|Mux15~9_combout ),
	.Mux151(\RF|Mux15~19_combout ),
	.Mux16(\RF|Mux16~9_combout ),
	.Mux161(\RF|Mux16~19_combout ),
	.Mux17(\RF|Mux17~9_combout ),
	.Mux171(\RF|Mux17~19_combout ),
	.Mux18(\RF|Mux18~9_combout ),
	.Mux181(\RF|Mux18~19_combout ),
	.Mux19(\RF|Mux19~9_combout ),
	.Mux191(\RF|Mux19~19_combout ),
	.Mux20(\RF|Mux20~9_combout ),
	.Mux201(\RF|Mux20~19_combout ),
	.Mux21(\RF|Mux21~9_combout ),
	.Mux211(\RF|Mux21~19_combout ),
	.Mux22(\RF|Mux22~9_combout ),
	.Mux221(\RF|Mux22~19_combout ),
	.Mux59(\RF|Mux59~9_combout ),
	.Mux591(\RF|Mux59~19_combout ),
	.Mux0(\RF|Mux0~9_combout ),
	.Mux01(\RF|Mux0~19_combout ),
	.Mux2(\RF|Mux2~9_combout ),
	.Mux210(\RF|Mux2~19_combout ),
	.Mux1(\RF|Mux1~9_combout ),
	.Mux11(\RF|Mux1~19_combout ),
	.Mux3(\RF|Mux3~9_combout ),
	.Mux31(\RF|Mux3~19_combout ),
	.Mux4(\RF|Mux4~9_combout ),
	.Mux410(\RF|Mux4~19_combout ),
	.Mux5(\RF|Mux5~9_combout ),
	.Mux510(\RF|Mux5~19_combout ),
	.Mux6(\RF|Mux6~9_combout ),
	.Mux64(\RF|Mux6~19_combout ),
	.Mux7(\RF|Mux7~9_combout ),
	.Mux71(\RF|Mux7~19_combout ),
	.Mux8(\RF|Mux8~9_combout ),
	.Mux81(\RF|Mux8~19_combout ),
	.Mux9(\RF|Mux9~9_combout ),
	.Mux91(\RF|Mux9~19_combout ),
	.Mux10(\RF|Mux10~9_combout ),
	.Mux101(\RF|Mux10~19_combout ),
	.Mux111(\RF|Mux11~9_combout ),
	.Mux112(\RF|Mux11~19_combout ),
	.Mux12(\RF|Mux12~9_combout ),
	.Mux121(\RF|Mux12~19_combout ),
	.Mux13(\RF|Mux13~9_combout ),
	.Mux131(\RF|Mux13~19_combout ),
	.Mux14(\RF|Mux14~9_combout ),
	.Mux141(\RF|Mux14~19_combout ),
	.Mux311(\RF|Mux31~9_combout ),
	.Mux312(\RF|Mux31~19_combout ),
	.CLK(CLK),
	.nRST(nRST),
	.devpor(devpor),
	.devclrn(devclrn),
	.devoe(devoe));

// Location: LCCOMB_X57_Y37_N18
cycloneive_lcell_comb \portb~0 (
// Equation(s):
// \portb~0_combout  = plif_exmemwsel_l_4 $ (!plif_idexrsel2_l_4)

	.dataa(gnd),
	.datab(\EXMEM|plif_exmem.wsel_l [4]),
	.datac(gnd),
	.datad(\IDEX|plif_idex.rsel2_l [4]),
	.cin(gnd),
	.combout(\portb~0_combout ),
	.cout());
// synopsys translate_off
defparam \portb~0 .lut_mask = 16'hCC33;
defparam \portb~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y37_N2
cycloneive_lcell_comb \portb~1 (
// Equation(s):
// \portb~1_combout  = (plif_idexalusrc_l) # ((\portb~0_combout  & (always01 & always0)))

	.dataa(\IDEX|plif_idex.alusrc_l~q ),
	.datab(\portb~0_combout ),
	.datac(\FU|always0~3_combout ),
	.datad(\FU|always0~2_combout ),
	.cin(gnd),
	.combout(\portb~1_combout ),
	.cout());
// synopsys translate_off
defparam \portb~1 .lut_mask = 16'hEAAA;
defparam \portb~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y41_N0
cycloneive_lcell_comb \wdat[31]~0 (
// Equation(s):
// \wdat[31]~0_combout  = (!plif_memwbregsrc_l_1 & ((plif_memwbregsrc_l_0 & ((plif_memwbdmemload_l_31))) # (!plif_memwbregsrc_l_0 & (plif_memwbporto_l_31))))

	.dataa(\MEMWB|plif_memwb.regsrc_l [0]),
	.datab(\MEMWB|plif_memwb.porto_l [31]),
	.datac(\MEMWB|plif_memwb.dmemload_l [31]),
	.datad(\MEMWB|plif_memwb.regsrc_l [1]),
	.cin(gnd),
	.combout(\wdat[31]~0_combout ),
	.cout());
// synopsys translate_off
defparam \wdat[31]~0 .lut_mask = 16'h00E4;
defparam \wdat[31]~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y41_N10
cycloneive_lcell_comb \wdat[31]~1 (
// Equation(s):
// \wdat[31]~1_combout  = (\wdat[31]~0_combout ) # ((plif_memwbrtnaddr_l_31 & plif_memwbregsrc_l_1))

	.dataa(\MEMWB|plif_memwb.rtnaddr_l [31]),
	.datab(\MEMWB|plif_memwb.regsrc_l [1]),
	.datac(gnd),
	.datad(\wdat[31]~0_combout ),
	.cin(gnd),
	.combout(\wdat[31]~1_combout ),
	.cout());
// synopsys translate_off
defparam \wdat[31]~1 .lut_mask = 16'hFF88;
defparam \wdat[31]~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y37_N24
cycloneive_lcell_comb \portb~2 (
// Equation(s):
// \portb~2_combout  = (!plif_idexalusrc_l & ((always02) # ((plif_memwbregen_l & fwdc))))

	.dataa(\FU|always0~4_combout ),
	.datab(\IDEX|plif_idex.alusrc_l~q ),
	.datac(\MEMWB|plif_memwb.regen_l~q ),
	.datad(\FU|fwdc~2_combout ),
	.cin(gnd),
	.combout(\portb~2_combout ),
	.cout());
// synopsys translate_off
defparam \portb~2 .lut_mask = 16'h3222;
defparam \portb~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y41_N20
cycloneive_lcell_comb \portb~3 (
// Equation(s):
// \portb~3_combout  = (\portb~2_combout  & ((\wdat[31]~1_combout ) # ((\portb~1_combout )))) # (!\portb~2_combout  & (((plif_idexrdat2_l_31 & !\portb~1_combout ))))

	.dataa(\wdat[31]~1_combout ),
	.datab(\IDEX|plif_idex.rdat2_l [31]),
	.datac(\portb~2_combout ),
	.datad(\portb~1_combout ),
	.cin(gnd),
	.combout(\portb~3_combout ),
	.cout());
// synopsys translate_off
defparam \portb~3 .lut_mask = 16'hF0AC;
defparam \portb~3 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y41_N26
cycloneive_lcell_comb \portb~4 (
// Equation(s):
// \portb~4_combout  = (\portb~1_combout  & ((\portb~3_combout  & (plif_exmemporto_l_31)) # (!\portb~3_combout  & ((plif_idexextimm_l_31))))) # (!\portb~1_combout  & (((\portb~3_combout ))))

	.dataa(\portb~1_combout ),
	.datab(plif_exmemporto_l_31),
	.datac(\IDEX|plif_idex.extimm_l [31]),
	.datad(\portb~3_combout ),
	.cin(gnd),
	.combout(\portb~4_combout ),
	.cout());
// synopsys translate_off
defparam \portb~4 .lut_mask = 16'hDDA0;
defparam \portb~4 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y42_N10
cycloneive_lcell_comb \wdat[30]~2 (
// Equation(s):
// \wdat[30]~2_combout  = (!plif_memwbregsrc_l_1 & ((plif_memwbregsrc_l_0 & ((plif_memwbdmemload_l_30))) # (!plif_memwbregsrc_l_0 & (plif_memwbporto_l_30))))

	.dataa(\MEMWB|plif_memwb.regsrc_l [0]),
	.datab(\MEMWB|plif_memwb.porto_l [30]),
	.datac(\MEMWB|plif_memwb.dmemload_l [30]),
	.datad(\MEMWB|plif_memwb.regsrc_l [1]),
	.cin(gnd),
	.combout(\wdat[30]~2_combout ),
	.cout());
// synopsys translate_off
defparam \wdat[30]~2 .lut_mask = 16'h00E4;
defparam \wdat[30]~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y42_N22
cycloneive_lcell_comb \wdat[30]~3 (
// Equation(s):
// \wdat[30]~3_combout  = (\wdat[30]~2_combout ) # ((plif_memwbrtnaddr_l_30 & plif_memwbregsrc_l_1))

	.dataa(\wdat[30]~2_combout ),
	.datab(\MEMWB|plif_memwb.rtnaddr_l [30]),
	.datac(gnd),
	.datad(\MEMWB|plif_memwb.regsrc_l [1]),
	.cin(gnd),
	.combout(\wdat[30]~3_combout ),
	.cout());
// synopsys translate_off
defparam \wdat[30]~3 .lut_mask = 16'hEEAA;
defparam \wdat[30]~3 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y42_N24
cycloneive_lcell_comb \portb~5 (
// Equation(s):
// \portb~5_combout  = (\portb~1_combout  & ((plif_idexextimm_l_30) # ((\portb~2_combout )))) # (!\portb~1_combout  & (((plif_idexrdat2_l_30 & !\portb~2_combout ))))

	.dataa(\IDEX|plif_idex.extimm_l [30]),
	.datab(\IDEX|plif_idex.rdat2_l [30]),
	.datac(\portb~1_combout ),
	.datad(\portb~2_combout ),
	.cin(gnd),
	.combout(\portb~5_combout ),
	.cout());
// synopsys translate_off
defparam \portb~5 .lut_mask = 16'hF0AC;
defparam \portb~5 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y42_N8
cycloneive_lcell_comb \portb~6 (
// Equation(s):
// \portb~6_combout  = (\portb~2_combout  & ((\portb~5_combout  & ((plif_exmemporto_l_30))) # (!\portb~5_combout  & (\wdat[30]~3_combout )))) # (!\portb~2_combout  & (((\portb~5_combout ))))

	.dataa(\wdat[30]~3_combout ),
	.datab(\portb~2_combout ),
	.datac(plif_exmemporto_l_30),
	.datad(\portb~5_combout ),
	.cin(gnd),
	.combout(\portb~6_combout ),
	.cout());
// synopsys translate_off
defparam \portb~6 .lut_mask = 16'hF388;
defparam \portb~6 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y35_N28
cycloneive_lcell_comb \wdat[29]~4 (
// Equation(s):
// \wdat[29]~4_combout  = (!plif_memwbregsrc_l_1 & ((plif_memwbregsrc_l_0 & (plif_memwbdmemload_l_29)) # (!plif_memwbregsrc_l_0 & ((plif_memwbporto_l_29)))))

	.dataa(\MEMWB|plif_memwb.regsrc_l [1]),
	.datab(\MEMWB|plif_memwb.regsrc_l [0]),
	.datac(\MEMWB|plif_memwb.dmemload_l [29]),
	.datad(\MEMWB|plif_memwb.porto_l [29]),
	.cin(gnd),
	.combout(\wdat[29]~4_combout ),
	.cout());
// synopsys translate_off
defparam \wdat[29]~4 .lut_mask = 16'h5140;
defparam \wdat[29]~4 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y35_N24
cycloneive_lcell_comb \wdat[29]~5 (
// Equation(s):
// \wdat[29]~5_combout  = (\wdat[29]~4_combout ) # ((plif_memwbregsrc_l_1 & plif_memwbrtnaddr_l_29))

	.dataa(\MEMWB|plif_memwb.regsrc_l [1]),
	.datab(\MEMWB|plif_memwb.rtnaddr_l [29]),
	.datac(gnd),
	.datad(\wdat[29]~4_combout ),
	.cin(gnd),
	.combout(\wdat[29]~5_combout ),
	.cout());
// synopsys translate_off
defparam \wdat[29]~5 .lut_mask = 16'hFF88;
defparam \wdat[29]~5 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y35_N26
cycloneive_lcell_comb \portb~7 (
// Equation(s):
// \portb~7_combout  = (\portb~1_combout  & (((\portb~2_combout )))) # (!\portb~1_combout  & ((\portb~2_combout  & ((\wdat[29]~5_combout ))) # (!\portb~2_combout  & (plif_idexrdat2_l_29))))

	.dataa(\IDEX|plif_idex.rdat2_l [29]),
	.datab(\portb~1_combout ),
	.datac(\wdat[29]~5_combout ),
	.datad(\portb~2_combout ),
	.cin(gnd),
	.combout(\portb~7_combout ),
	.cout());
// synopsys translate_off
defparam \portb~7 .lut_mask = 16'hFC22;
defparam \portb~7 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y35_N16
cycloneive_lcell_comb \portb~8 (
// Equation(s):
// \portb~8_combout  = (\portb~1_combout  & ((\portb~7_combout  & ((plif_exmemporto_l_29))) # (!\portb~7_combout  & (plif_idexextimm_l_29)))) # (!\portb~1_combout  & (((\portb~7_combout ))))

	.dataa(\IDEX|plif_idex.extimm_l [29]),
	.datab(\portb~1_combout ),
	.datac(\portb~7_combout ),
	.datad(plif_exmemporto_l_29),
	.cin(gnd),
	.combout(\portb~8_combout ),
	.cout());
// synopsys translate_off
defparam \portb~8 .lut_mask = 16'hF838;
defparam \portb~8 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y35_N20
cycloneive_lcell_comb \wdat[28]~6 (
// Equation(s):
// \wdat[28]~6_combout  = (!plif_memwbregsrc_l_1 & ((plif_memwbregsrc_l_0 & (plif_memwbdmemload_l_28)) # (!plif_memwbregsrc_l_0 & ((plif_memwbporto_l_28)))))

	.dataa(\MEMWB|plif_memwb.regsrc_l [1]),
	.datab(\MEMWB|plif_memwb.regsrc_l [0]),
	.datac(\MEMWB|plif_memwb.dmemload_l [28]),
	.datad(\MEMWB|plif_memwb.porto_l [28]),
	.cin(gnd),
	.combout(\wdat[28]~6_combout ),
	.cout());
// synopsys translate_off
defparam \wdat[28]~6 .lut_mask = 16'h5140;
defparam \wdat[28]~6 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y35_N6
cycloneive_lcell_comb \wdat[28]~7 (
// Equation(s):
// \wdat[28]~7_combout  = (\wdat[28]~6_combout ) # ((plif_memwbregsrc_l_1 & plif_memwbrtnaddr_l_28))

	.dataa(\MEMWB|plif_memwb.regsrc_l [1]),
	.datab(\MEMWB|plif_memwb.rtnaddr_l [28]),
	.datac(gnd),
	.datad(\wdat[28]~6_combout ),
	.cin(gnd),
	.combout(\wdat[28]~7_combout ),
	.cout());
// synopsys translate_off
defparam \wdat[28]~7 .lut_mask = 16'hFF88;
defparam \wdat[28]~7 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y35_N0
cycloneive_lcell_comb \portb~9 (
// Equation(s):
// \portb~9_combout  = (\portb~1_combout  & (((\portb~2_combout ) # (plif_idexextimm_l_28)))) # (!\portb~1_combout  & (plif_idexrdat2_l_28 & (!\portb~2_combout )))

	.dataa(\portb~1_combout ),
	.datab(\IDEX|plif_idex.rdat2_l [28]),
	.datac(\portb~2_combout ),
	.datad(\IDEX|plif_idex.extimm_l [28]),
	.cin(gnd),
	.combout(\portb~9_combout ),
	.cout());
// synopsys translate_off
defparam \portb~9 .lut_mask = 16'hAEA4;
defparam \portb~9 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y35_N14
cycloneive_lcell_comb \portb~10 (
// Equation(s):
// \portb~10_combout  = (\portb~2_combout  & ((\portb~9_combout  & ((plif_exmemporto_l_28))) # (!\portb~9_combout  & (\wdat[28]~7_combout )))) # (!\portb~2_combout  & (((\portb~9_combout ))))

	.dataa(\wdat[28]~7_combout ),
	.datab(plif_exmemporto_l_28),
	.datac(\portb~2_combout ),
	.datad(\portb~9_combout ),
	.cin(gnd),
	.combout(\portb~10_combout ),
	.cout());
// synopsys translate_off
defparam \portb~10 .lut_mask = 16'hCFA0;
defparam \portb~10 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y36_N20
cycloneive_lcell_comb \wdat[27]~8 (
// Equation(s):
// \wdat[27]~8_combout  = (!plif_memwbregsrc_l_1 & ((plif_memwbregsrc_l_0 & ((plif_memwbdmemload_l_27))) # (!plif_memwbregsrc_l_0 & (plif_memwbporto_l_27))))

	.dataa(\MEMWB|plif_memwb.regsrc_l [1]),
	.datab(\MEMWB|plif_memwb.porto_l [27]),
	.datac(\MEMWB|plif_memwb.dmemload_l [27]),
	.datad(\MEMWB|plif_memwb.regsrc_l [0]),
	.cin(gnd),
	.combout(\wdat[27]~8_combout ),
	.cout());
// synopsys translate_off
defparam \wdat[27]~8 .lut_mask = 16'h5044;
defparam \wdat[27]~8 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y36_N0
cycloneive_lcell_comb \wdat[27]~9 (
// Equation(s):
// \wdat[27]~9_combout  = (\wdat[27]~8_combout ) # ((plif_memwbregsrc_l_1 & plif_memwbrtnaddr_l_27))

	.dataa(gnd),
	.datab(\MEMWB|plif_memwb.regsrc_l [1]),
	.datac(\MEMWB|plif_memwb.rtnaddr_l [27]),
	.datad(\wdat[27]~8_combout ),
	.cin(gnd),
	.combout(\wdat[27]~9_combout ),
	.cout());
// synopsys translate_off
defparam \wdat[27]~9 .lut_mask = 16'hFFC0;
defparam \wdat[27]~9 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y36_N6
cycloneive_lcell_comb \portb~11 (
// Equation(s):
// \portb~11_combout  = (\portb~2_combout  & (((\wdat[27]~9_combout ) # (\portb~1_combout )))) # (!\portb~2_combout  & (plif_idexrdat2_l_27 & ((!\portb~1_combout ))))

	.dataa(\IDEX|plif_idex.rdat2_l [27]),
	.datab(\wdat[27]~9_combout ),
	.datac(\portb~2_combout ),
	.datad(\portb~1_combout ),
	.cin(gnd),
	.combout(\portb~11_combout ),
	.cout());
// synopsys translate_off
defparam \portb~11 .lut_mask = 16'hF0CA;
defparam \portb~11 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y36_N24
cycloneive_lcell_comb \portb~12 (
// Equation(s):
// \portb~12_combout  = (\portb~1_combout  & ((\portb~11_combout  & (plif_exmemporto_l_27)) # (!\portb~11_combout  & ((plif_idexextimm_l_27))))) # (!\portb~1_combout  & (((\portb~11_combout ))))

	.dataa(plif_exmemporto_l_27),
	.datab(\IDEX|plif_idex.extimm_l [27]),
	.datac(\portb~1_combout ),
	.datad(\portb~11_combout ),
	.cin(gnd),
	.combout(\portb~12_combout ),
	.cout());
// synopsys translate_off
defparam \portb~12 .lut_mask = 16'hAFC0;
defparam \portb~12 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y36_N4
cycloneive_lcell_comb \wdat[26]~10 (
// Equation(s):
// \wdat[26]~10_combout  = (!plif_memwbregsrc_l_1 & ((plif_memwbregsrc_l_0 & ((plif_memwbdmemload_l_26))) # (!plif_memwbregsrc_l_0 & (plif_memwbporto_l_26))))

	.dataa(\MEMWB|plif_memwb.regsrc_l [1]),
	.datab(\MEMWB|plif_memwb.porto_l [26]),
	.datac(\MEMWB|plif_memwb.dmemload_l [26]),
	.datad(\MEMWB|plif_memwb.regsrc_l [0]),
	.cin(gnd),
	.combout(\wdat[26]~10_combout ),
	.cout());
// synopsys translate_off
defparam \wdat[26]~10 .lut_mask = 16'h5044;
defparam \wdat[26]~10 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y36_N6
cycloneive_lcell_comb \wdat[26]~11 (
// Equation(s):
// \wdat[26]~11_combout  = (\wdat[26]~10_combout ) # ((plif_memwbrtnaddr_l_26 & plif_memwbregsrc_l_1))

	.dataa(\MEMWB|plif_memwb.rtnaddr_l [26]),
	.datab(\wdat[26]~10_combout ),
	.datac(gnd),
	.datad(\MEMWB|plif_memwb.regsrc_l [1]),
	.cin(gnd),
	.combout(\wdat[26]~11_combout ),
	.cout());
// synopsys translate_off
defparam \wdat[26]~11 .lut_mask = 16'hEECC;
defparam \wdat[26]~11 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y36_N12
cycloneive_lcell_comb \portb~13 (
// Equation(s):
// \portb~13_combout  = (\portb~1_combout  & (((\portb~2_combout ) # (plif_idexextimm_l_26)))) # (!\portb~1_combout  & (plif_idexrdat2_l_26 & (!\portb~2_combout )))

	.dataa(\portb~1_combout ),
	.datab(\IDEX|plif_idex.rdat2_l [26]),
	.datac(\portb~2_combout ),
	.datad(\IDEX|plif_idex.extimm_l [26]),
	.cin(gnd),
	.combout(\portb~13_combout ),
	.cout());
// synopsys translate_off
defparam \portb~13 .lut_mask = 16'hAEA4;
defparam \portb~13 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y36_N10
cycloneive_lcell_comb \portb~14 (
// Equation(s):
// \portb~14_combout  = (\portb~2_combout  & ((\portb~13_combout  & ((plif_exmemporto_l_26))) # (!\portb~13_combout  & (\wdat[26]~11_combout )))) # (!\portb~2_combout  & (((\portb~13_combout ))))

	.dataa(\wdat[26]~11_combout ),
	.datab(plif_exmemporto_l_26),
	.datac(\portb~2_combout ),
	.datad(\portb~13_combout ),
	.cin(gnd),
	.combout(\portb~14_combout ),
	.cout());
// synopsys translate_off
defparam \portb~14 .lut_mask = 16'hCFA0;
defparam \portb~14 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y36_N14
cycloneive_lcell_comb \wdat[25]~12 (
// Equation(s):
// \wdat[25]~12_combout  = (!plif_memwbregsrc_l_1 & ((plif_memwbregsrc_l_0 & ((plif_memwbdmemload_l_25))) # (!plif_memwbregsrc_l_0 & (plif_memwbporto_l_25))))

	.dataa(\MEMWB|plif_memwb.regsrc_l [1]),
	.datab(\MEMWB|plif_memwb.porto_l [25]),
	.datac(\MEMWB|plif_memwb.dmemload_l [25]),
	.datad(\MEMWB|plif_memwb.regsrc_l [0]),
	.cin(gnd),
	.combout(\wdat[25]~12_combout ),
	.cout());
// synopsys translate_off
defparam \wdat[25]~12 .lut_mask = 16'h5044;
defparam \wdat[25]~12 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y36_N30
cycloneive_lcell_comb \wdat[25]~13 (
// Equation(s):
// \wdat[25]~13_combout  = (\wdat[25]~12_combout ) # ((plif_memwbregsrc_l_1 & plif_memwbrtnaddr_l_25))

	.dataa(gnd),
	.datab(\MEMWB|plif_memwb.regsrc_l [1]),
	.datac(\MEMWB|plif_memwb.rtnaddr_l [25]),
	.datad(\wdat[25]~12_combout ),
	.cin(gnd),
	.combout(\wdat[25]~13_combout ),
	.cout());
// synopsys translate_off
defparam \wdat[25]~13 .lut_mask = 16'hFFC0;
defparam \wdat[25]~13 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y36_N12
cycloneive_lcell_comb \portb~15 (
// Equation(s):
// \portb~15_combout  = (\portb~2_combout  & ((\wdat[25]~13_combout ) # ((\portb~1_combout )))) # (!\portb~2_combout  & (((plif_idexrdat2_l_25 & !\portb~1_combout ))))

	.dataa(\wdat[25]~13_combout ),
	.datab(\IDEX|plif_idex.rdat2_l [25]),
	.datac(\portb~2_combout ),
	.datad(\portb~1_combout ),
	.cin(gnd),
	.combout(\portb~15_combout ),
	.cout());
// synopsys translate_off
defparam \portb~15 .lut_mask = 16'hF0AC;
defparam \portb~15 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y36_N22
cycloneive_lcell_comb \portb~16 (
// Equation(s):
// \portb~16_combout  = (\portb~1_combout  & ((\portb~15_combout  & ((plif_exmemporto_l_25))) # (!\portb~15_combout  & (plif_idexextimm_l_25)))) # (!\portb~1_combout  & (((\portb~15_combout ))))

	.dataa(\IDEX|plif_idex.extimm_l [25]),
	.datab(\portb~1_combout ),
	.datac(plif_exmemporto_l_25),
	.datad(\portb~15_combout ),
	.cin(gnd),
	.combout(\portb~16_combout ),
	.cout());
// synopsys translate_off
defparam \portb~16 .lut_mask = 16'hF388;
defparam \portb~16 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y35_N14
cycloneive_lcell_comb \wdat[24]~14 (
// Equation(s):
// \wdat[24]~14_combout  = (!plif_memwbregsrc_l_1 & ((plif_memwbregsrc_l_0 & ((plif_memwbdmemload_l_24))) # (!plif_memwbregsrc_l_0 & (plif_memwbporto_l_24))))

	.dataa(\MEMWB|plif_memwb.regsrc_l [0]),
	.datab(\MEMWB|plif_memwb.porto_l [24]),
	.datac(\MEMWB|plif_memwb.dmemload_l [24]),
	.datad(\MEMWB|plif_memwb.regsrc_l [1]),
	.cin(gnd),
	.combout(\wdat[24]~14_combout ),
	.cout());
// synopsys translate_off
defparam \wdat[24]~14 .lut_mask = 16'h00E4;
defparam \wdat[24]~14 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y35_N2
cycloneive_lcell_comb \wdat[24]~15 (
// Equation(s):
// \wdat[24]~15_combout  = (\wdat[24]~14_combout ) # ((plif_memwbrtnaddr_l_24 & plif_memwbregsrc_l_1))

	.dataa(gnd),
	.datab(\wdat[24]~14_combout ),
	.datac(\MEMWB|plif_memwb.rtnaddr_l [24]),
	.datad(\MEMWB|plif_memwb.regsrc_l [1]),
	.cin(gnd),
	.combout(\wdat[24]~15_combout ),
	.cout());
// synopsys translate_off
defparam \wdat[24]~15 .lut_mask = 16'hFCCC;
defparam \wdat[24]~15 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y35_N8
cycloneive_lcell_comb \portb~17 (
// Equation(s):
// \portb~17_combout  = (\portb~2_combout  & (((\portb~1_combout )))) # (!\portb~2_combout  & ((\portb~1_combout  & ((plif_idexextimm_l_24))) # (!\portb~1_combout  & (plif_idexrdat2_l_24))))

	.dataa(\IDEX|plif_idex.rdat2_l [24]),
	.datab(\IDEX|plif_idex.extimm_l [24]),
	.datac(\portb~2_combout ),
	.datad(\portb~1_combout ),
	.cin(gnd),
	.combout(\portb~17_combout ),
	.cout());
// synopsys translate_off
defparam \portb~17 .lut_mask = 16'hFC0A;
defparam \portb~17 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y35_N22
cycloneive_lcell_comb \portb~18 (
// Equation(s):
// \portb~18_combout  = (\portb~2_combout  & ((\portb~17_combout  & ((plif_exmemporto_l_24))) # (!\portb~17_combout  & (\wdat[24]~15_combout )))) # (!\portb~2_combout  & (((\portb~17_combout ))))

	.dataa(\portb~2_combout ),
	.datab(\wdat[24]~15_combout ),
	.datac(\portb~17_combout ),
	.datad(plif_exmemporto_l_24),
	.cin(gnd),
	.combout(\portb~18_combout ),
	.cout());
// synopsys translate_off
defparam \portb~18 .lut_mask = 16'hF858;
defparam \portb~18 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y35_N10
cycloneive_lcell_comb \wdat[23]~16 (
// Equation(s):
// \wdat[23]~16_combout  = (!plif_memwbregsrc_l_1 & ((plif_memwbregsrc_l_0 & (plif_memwbdmemload_l_23)) # (!plif_memwbregsrc_l_0 & ((plif_memwbporto_l_23)))))

	.dataa(\MEMWB|plif_memwb.regsrc_l [1]),
	.datab(\MEMWB|plif_memwb.regsrc_l [0]),
	.datac(\MEMWB|plif_memwb.dmemload_l [23]),
	.datad(\MEMWB|plif_memwb.porto_l [23]),
	.cin(gnd),
	.combout(\wdat[23]~16_combout ),
	.cout());
// synopsys translate_off
defparam \wdat[23]~16 .lut_mask = 16'h5140;
defparam \wdat[23]~16 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X52_Y39_N2
cycloneive_lcell_comb \wdat[23]~17 (
// Equation(s):
// \wdat[23]~17_combout  = (\wdat[23]~16_combout ) # ((plif_memwbrtnaddr_l_23 & plif_memwbregsrc_l_1))

	.dataa(\wdat[23]~16_combout ),
	.datab(gnd),
	.datac(\MEMWB|plif_memwb.rtnaddr_l [23]),
	.datad(\MEMWB|plif_memwb.regsrc_l [1]),
	.cin(gnd),
	.combout(\wdat[23]~17_combout ),
	.cout());
// synopsys translate_off
defparam \wdat[23]~17 .lut_mask = 16'hFAAA;
defparam \wdat[23]~17 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X52_Y39_N20
cycloneive_lcell_comb \portb~19 (
// Equation(s):
// \portb~19_combout  = (\portb~1_combout  & (((\portb~2_combout )))) # (!\portb~1_combout  & ((\portb~2_combout  & ((\wdat[23]~17_combout ))) # (!\portb~2_combout  & (plif_idexrdat2_l_23))))

	.dataa(\IDEX|plif_idex.rdat2_l [23]),
	.datab(\wdat[23]~17_combout ),
	.datac(\portb~1_combout ),
	.datad(\portb~2_combout ),
	.cin(gnd),
	.combout(\portb~19_combout ),
	.cout());
// synopsys translate_off
defparam \portb~19 .lut_mask = 16'hFC0A;
defparam \portb~19 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X52_Y39_N30
cycloneive_lcell_comb \portb~20 (
// Equation(s):
// \portb~20_combout  = (\portb~1_combout  & ((\portb~19_combout  & (plif_exmemporto_l_23)) # (!\portb~19_combout  & ((plif_idexextimm_l_23))))) # (!\portb~1_combout  & (((\portb~19_combout ))))

	.dataa(plif_exmemporto_l_23),
	.datab(\IDEX|plif_idex.extimm_l [23]),
	.datac(\portb~1_combout ),
	.datad(\portb~19_combout ),
	.cin(gnd),
	.combout(\portb~20_combout ),
	.cout());
// synopsys translate_off
defparam \portb~20 .lut_mask = 16'hAFC0;
defparam \portb~20 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y39_N4
cycloneive_lcell_comb \wdat[22]~18 (
// Equation(s):
// \wdat[22]~18_combout  = (!plif_memwbregsrc_l_1 & ((plif_memwbregsrc_l_0 & ((plif_memwbdmemload_l_22))) # (!plif_memwbregsrc_l_0 & (plif_memwbporto_l_22))))

	.dataa(\MEMWB|plif_memwb.porto_l [22]),
	.datab(\MEMWB|plif_memwb.regsrc_l [0]),
	.datac(\MEMWB|plif_memwb.dmemload_l [22]),
	.datad(\MEMWB|plif_memwb.regsrc_l [1]),
	.cin(gnd),
	.combout(\wdat[22]~18_combout ),
	.cout());
// synopsys translate_off
defparam \wdat[22]~18 .lut_mask = 16'h00E2;
defparam \wdat[22]~18 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y39_N14
cycloneive_lcell_comb \wdat[22]~19 (
// Equation(s):
// \wdat[22]~19_combout  = (\wdat[22]~18_combout ) # ((plif_memwbrtnaddr_l_22 & plif_memwbregsrc_l_1))

	.dataa(\MEMWB|plif_memwb.rtnaddr_l [22]),
	.datab(\MEMWB|plif_memwb.regsrc_l [1]),
	.datac(gnd),
	.datad(\wdat[22]~18_combout ),
	.cin(gnd),
	.combout(\wdat[22]~19_combout ),
	.cout());
// synopsys translate_off
defparam \wdat[22]~19 .lut_mask = 16'hFF88;
defparam \wdat[22]~19 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y39_N16
cycloneive_lcell_comb \portb~21 (
// Equation(s):
// \portb~21_combout  = (\portb~1_combout  & ((plif_idexextimm_l_22) # ((\portb~2_combout )))) # (!\portb~1_combout  & (((plif_idexrdat2_l_22 & !\portb~2_combout ))))

	.dataa(\IDEX|plif_idex.extimm_l [22]),
	.datab(\IDEX|plif_idex.rdat2_l [22]),
	.datac(\portb~1_combout ),
	.datad(\portb~2_combout ),
	.cin(gnd),
	.combout(\portb~21_combout ),
	.cout());
// synopsys translate_off
defparam \portb~21 .lut_mask = 16'hF0AC;
defparam \portb~21 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y39_N22
cycloneive_lcell_comb \portb~22 (
// Equation(s):
// \portb~22_combout  = (\portb~2_combout  & ((\portb~21_combout  & (plif_exmemporto_l_22)) # (!\portb~21_combout  & ((\wdat[22]~19_combout ))))) # (!\portb~2_combout  & (((\portb~21_combout ))))

	.dataa(\portb~2_combout ),
	.datab(plif_exmemporto_l_22),
	.datac(\wdat[22]~19_combout ),
	.datad(\portb~21_combout ),
	.cin(gnd),
	.combout(\portb~22_combout ),
	.cout());
// synopsys translate_off
defparam \portb~22 .lut_mask = 16'hDDA0;
defparam \portb~22 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y35_N20
cycloneive_lcell_comb \wdat[21]~20 (
// Equation(s):
// \wdat[21]~20_combout  = (!plif_memwbregsrc_l_1 & ((plif_memwbregsrc_l_0 & ((plif_memwbdmemload_l_21))) # (!plif_memwbregsrc_l_0 & (plif_memwbporto_l_21))))

	.dataa(\MEMWB|plif_memwb.porto_l [21]),
	.datab(\MEMWB|plif_memwb.regsrc_l [0]),
	.datac(\MEMWB|plif_memwb.dmemload_l [21]),
	.datad(\MEMWB|plif_memwb.regsrc_l [1]),
	.cin(gnd),
	.combout(\wdat[21]~20_combout ),
	.cout());
// synopsys translate_off
defparam \wdat[21]~20 .lut_mask = 16'h00E2;
defparam \wdat[21]~20 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y35_N0
cycloneive_lcell_comb \wdat[21]~21 (
// Equation(s):
// \wdat[21]~21_combout  = (\wdat[21]~20_combout ) # ((plif_memwbregsrc_l_1 & plif_memwbrtnaddr_l_21))

	.dataa(\MEMWB|plif_memwb.regsrc_l [1]),
	.datab(gnd),
	.datac(\MEMWB|plif_memwb.rtnaddr_l [21]),
	.datad(\wdat[21]~20_combout ),
	.cin(gnd),
	.combout(\wdat[21]~21_combout ),
	.cout());
// synopsys translate_off
defparam \wdat[21]~21 .lut_mask = 16'hFFA0;
defparam \wdat[21]~21 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y35_N2
cycloneive_lcell_comb \portb~23 (
// Equation(s):
// \portb~23_combout  = (\portb~1_combout  & (((\portb~2_combout )))) # (!\portb~1_combout  & ((\portb~2_combout  & (\wdat[21]~21_combout )) # (!\portb~2_combout  & ((plif_idexrdat2_l_21)))))

	.dataa(\portb~1_combout ),
	.datab(\wdat[21]~21_combout ),
	.datac(\IDEX|plif_idex.rdat2_l [21]),
	.datad(\portb~2_combout ),
	.cin(gnd),
	.combout(\portb~23_combout ),
	.cout());
// synopsys translate_off
defparam \portb~23 .lut_mask = 16'hEE50;
defparam \portb~23 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y35_N12
cycloneive_lcell_comb \portb~24 (
// Equation(s):
// \portb~24_combout  = (\portb~1_combout  & ((\portb~23_combout  & ((plif_exmemporto_l_21))) # (!\portb~23_combout  & (plif_idexextimm_l_21)))) # (!\portb~1_combout  & (((\portb~23_combout ))))

	.dataa(\IDEX|plif_idex.extimm_l [21]),
	.datab(\portb~1_combout ),
	.datac(plif_exmemporto_l_21),
	.datad(\portb~23_combout ),
	.cin(gnd),
	.combout(\portb~24_combout ),
	.cout());
// synopsys translate_off
defparam \portb~24 .lut_mask = 16'hF388;
defparam \portb~24 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y39_N8
cycloneive_lcell_comb \wdat[20]~22 (
// Equation(s):
// \wdat[20]~22_combout  = (!plif_memwbregsrc_l_1 & ((plif_memwbregsrc_l_0 & ((plif_memwbdmemload_l_20))) # (!plif_memwbregsrc_l_0 & (plif_memwbporto_l_20))))

	.dataa(\MEMWB|plif_memwb.porto_l [20]),
	.datab(\MEMWB|plif_memwb.regsrc_l [0]),
	.datac(\MEMWB|plif_memwb.dmemload_l [20]),
	.datad(\MEMWB|plif_memwb.regsrc_l [1]),
	.cin(gnd),
	.combout(\wdat[20]~22_combout ),
	.cout());
// synopsys translate_off
defparam \wdat[20]~22 .lut_mask = 16'h00E2;
defparam \wdat[20]~22 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y39_N16
cycloneive_lcell_comb \wdat[20]~23 (
// Equation(s):
// \wdat[20]~23_combout  = (\wdat[20]~22_combout ) # ((plif_memwbrtnaddr_l_20 & plif_memwbregsrc_l_1))

	.dataa(gnd),
	.datab(\wdat[20]~22_combout ),
	.datac(\MEMWB|plif_memwb.rtnaddr_l [20]),
	.datad(\MEMWB|plif_memwb.regsrc_l [1]),
	.cin(gnd),
	.combout(\wdat[20]~23_combout ),
	.cout());
// synopsys translate_off
defparam \wdat[20]~23 .lut_mask = 16'hFCCC;
defparam \wdat[20]~23 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y39_N2
cycloneive_lcell_comb \portb~25 (
// Equation(s):
// \portb~25_combout  = (\portb~2_combout  & (((\portb~1_combout )))) # (!\portb~2_combout  & ((\portb~1_combout  & ((plif_idexextimm_l_20))) # (!\portb~1_combout  & (plif_idexrdat2_l_20))))

	.dataa(\IDEX|plif_idex.rdat2_l [20]),
	.datab(\IDEX|plif_idex.extimm_l [20]),
	.datac(\portb~2_combout ),
	.datad(\portb~1_combout ),
	.cin(gnd),
	.combout(\portb~25_combout ),
	.cout());
// synopsys translate_off
defparam \portb~25 .lut_mask = 16'hFC0A;
defparam \portb~25 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y39_N30
cycloneive_lcell_comb \portb~26 (
// Equation(s):
// \portb~26_combout  = (\portb~2_combout  & ((\portb~25_combout  & (plif_exmemporto_l_20)) # (!\portb~25_combout  & ((\wdat[20]~23_combout ))))) # (!\portb~2_combout  & (((\portb~25_combout ))))

	.dataa(plif_exmemporto_l_20),
	.datab(\wdat[20]~23_combout ),
	.datac(\portb~2_combout ),
	.datad(\portb~25_combout ),
	.cin(gnd),
	.combout(\portb~26_combout ),
	.cout());
// synopsys translate_off
defparam \portb~26 .lut_mask = 16'hAFC0;
defparam \portb~26 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y34_N28
cycloneive_lcell_comb \wdat[19]~24 (
// Equation(s):
// \wdat[19]~24_combout  = (!plif_memwbregsrc_l_1 & ((plif_memwbregsrc_l_0 & ((plif_memwbdmemload_l_19))) # (!plif_memwbregsrc_l_0 & (plif_memwbporto_l_19))))

	.dataa(\MEMWB|plif_memwb.regsrc_l [0]),
	.datab(\MEMWB|plif_memwb.porto_l [19]),
	.datac(\MEMWB|plif_memwb.dmemload_l [19]),
	.datad(\MEMWB|plif_memwb.regsrc_l [1]),
	.cin(gnd),
	.combout(\wdat[19]~24_combout ),
	.cout());
// synopsys translate_off
defparam \wdat[19]~24 .lut_mask = 16'h00E4;
defparam \wdat[19]~24 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y34_N24
cycloneive_lcell_comb \wdat[19]~25 (
// Equation(s):
// \wdat[19]~25_combout  = (\wdat[19]~24_combout ) # ((plif_memwbregsrc_l_1 & plif_memwbrtnaddr_l_19))

	.dataa(\MEMWB|plif_memwb.regsrc_l [1]),
	.datab(gnd),
	.datac(\MEMWB|plif_memwb.rtnaddr_l [19]),
	.datad(\wdat[19]~24_combout ),
	.cin(gnd),
	.combout(\wdat[19]~25_combout ),
	.cout());
// synopsys translate_off
defparam \wdat[19]~25 .lut_mask = 16'hFFA0;
defparam \wdat[19]~25 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y34_N6
cycloneive_lcell_comb \portb~27 (
// Equation(s):
// \portb~27_combout  = (\portb~1_combout  & (((\portb~2_combout )))) # (!\portb~1_combout  & ((\portb~2_combout  & ((\wdat[19]~25_combout ))) # (!\portb~2_combout  & (plif_idexrdat2_l_19))))

	.dataa(\IDEX|plif_idex.rdat2_l [19]),
	.datab(\wdat[19]~25_combout ),
	.datac(\portb~1_combout ),
	.datad(\portb~2_combout ),
	.cin(gnd),
	.combout(\portb~27_combout ),
	.cout());
// synopsys translate_off
defparam \portb~27 .lut_mask = 16'hFC0A;
defparam \portb~27 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y34_N20
cycloneive_lcell_comb \portb~28 (
// Equation(s):
// \portb~28_combout  = (\portb~1_combout  & ((\portb~27_combout  & (plif_exmemporto_l_19)) # (!\portb~27_combout  & ((plif_idexextimm_l_19))))) # (!\portb~1_combout  & (((\portb~27_combout ))))

	.dataa(plif_exmemporto_l_19),
	.datab(\IDEX|plif_idex.extimm_l [19]),
	.datac(\portb~1_combout ),
	.datad(\portb~27_combout ),
	.cin(gnd),
	.combout(\portb~28_combout ),
	.cout());
// synopsys translate_off
defparam \portb~28 .lut_mask = 16'hAFC0;
defparam \portb~28 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y37_N12
cycloneive_lcell_comb \wdat[18]~26 (
// Equation(s):
// \wdat[18]~26_combout  = (!plif_memwbregsrc_l_1 & ((plif_memwbregsrc_l_0 & ((plif_memwbdmemload_l_18))) # (!plif_memwbregsrc_l_0 & (plif_memwbporto_l_18))))

	.dataa(\MEMWB|plif_memwb.regsrc_l [1]),
	.datab(\MEMWB|plif_memwb.porto_l [18]),
	.datac(\MEMWB|plif_memwb.dmemload_l [18]),
	.datad(\MEMWB|plif_memwb.regsrc_l [0]),
	.cin(gnd),
	.combout(\wdat[18]~26_combout ),
	.cout());
// synopsys translate_off
defparam \wdat[18]~26 .lut_mask = 16'h5044;
defparam \wdat[18]~26 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y37_N14
cycloneive_lcell_comb \wdat[18]~27 (
// Equation(s):
// \wdat[18]~27_combout  = (\wdat[18]~26_combout ) # ((plif_memwbregsrc_l_1 & plif_memwbrtnaddr_l_18))

	.dataa(\MEMWB|plif_memwb.regsrc_l [1]),
	.datab(gnd),
	.datac(\MEMWB|plif_memwb.rtnaddr_l [18]),
	.datad(\wdat[18]~26_combout ),
	.cin(gnd),
	.combout(\wdat[18]~27_combout ),
	.cout());
// synopsys translate_off
defparam \wdat[18]~27 .lut_mask = 16'hFFA0;
defparam \wdat[18]~27 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y37_N20
cycloneive_lcell_comb \portb~29 (
// Equation(s):
// \portb~29_combout  = (\portb~1_combout  & ((plif_idexextimm_l_18) # ((\portb~2_combout )))) # (!\portb~1_combout  & (((plif_idexrdat2_l_18 & !\portb~2_combout ))))

	.dataa(\IDEX|plif_idex.extimm_l [18]),
	.datab(\IDEX|plif_idex.rdat2_l [18]),
	.datac(\portb~1_combout ),
	.datad(\portb~2_combout ),
	.cin(gnd),
	.combout(\portb~29_combout ),
	.cout());
// synopsys translate_off
defparam \portb~29 .lut_mask = 16'hF0AC;
defparam \portb~29 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y37_N2
cycloneive_lcell_comb \portb~30 (
// Equation(s):
// \portb~30_combout  = (\portb~2_combout  & ((\portb~29_combout  & (plif_exmemporto_l_18)) # (!\portb~29_combout  & ((\wdat[18]~27_combout ))))) # (!\portb~2_combout  & (((\portb~29_combout ))))

	.dataa(plif_exmemporto_l_18),
	.datab(\portb~2_combout ),
	.datac(\wdat[18]~27_combout ),
	.datad(\portb~29_combout ),
	.cin(gnd),
	.combout(\portb~30_combout ),
	.cout());
// synopsys translate_off
defparam \portb~30 .lut_mask = 16'hBBC0;
defparam \portb~30 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y35_N6
cycloneive_lcell_comb \wdat[17]~28 (
// Equation(s):
// \wdat[17]~28_combout  = (!plif_memwbregsrc_l_1 & ((plif_memwbregsrc_l_0 & (plif_memwbdmemload_l_17)) # (!plif_memwbregsrc_l_0 & ((plif_memwbporto_l_17)))))

	.dataa(\MEMWB|plif_memwb.regsrc_l [1]),
	.datab(\MEMWB|plif_memwb.regsrc_l [0]),
	.datac(\MEMWB|plif_memwb.dmemload_l [17]),
	.datad(\MEMWB|plif_memwb.porto_l [17]),
	.cin(gnd),
	.combout(\wdat[17]~28_combout ),
	.cout());
// synopsys translate_off
defparam \wdat[17]~28 .lut_mask = 16'h5140;
defparam \wdat[17]~28 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y35_N14
cycloneive_lcell_comb \wdat[17]~29 (
// Equation(s):
// \wdat[17]~29_combout  = (\wdat[17]~28_combout ) # ((plif_memwbregsrc_l_1 & plif_memwbrtnaddr_l_17))

	.dataa(\MEMWB|plif_memwb.regsrc_l [1]),
	.datab(\MEMWB|plif_memwb.rtnaddr_l [17]),
	.datac(gnd),
	.datad(\wdat[17]~28_combout ),
	.cin(gnd),
	.combout(\wdat[17]~29_combout ),
	.cout());
// synopsys translate_off
defparam \wdat[17]~29 .lut_mask = 16'hFF88;
defparam \wdat[17]~29 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y35_N18
cycloneive_lcell_comb \portb~31 (
// Equation(s):
// \portb~31_combout  = (\portb~1_combout  & (((\portb~2_combout )))) # (!\portb~1_combout  & ((\portb~2_combout  & (\wdat[17]~29_combout )) # (!\portb~2_combout  & ((plif_idexrdat2_l_17)))))

	.dataa(\wdat[17]~29_combout ),
	.datab(\portb~1_combout ),
	.datac(\IDEX|plif_idex.rdat2_l [17]),
	.datad(\portb~2_combout ),
	.cin(gnd),
	.combout(\portb~31_combout ),
	.cout());
// synopsys translate_off
defparam \portb~31 .lut_mask = 16'hEE30;
defparam \portb~31 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y35_N8
cycloneive_lcell_comb \portb~32 (
// Equation(s):
// \portb~32_combout  = (\portb~1_combout  & ((\portb~31_combout  & ((plif_exmemporto_l_17))) # (!\portb~31_combout  & (plif_idexextimm_l_17)))) # (!\portb~1_combout  & (((\portb~31_combout ))))

	.dataa(\IDEX|plif_idex.extimm_l [17]),
	.datab(\portb~1_combout ),
	.datac(plif_exmemporto_l_17),
	.datad(\portb~31_combout ),
	.cin(gnd),
	.combout(\portb~32_combout ),
	.cout());
// synopsys translate_off
defparam \portb~32 .lut_mask = 16'hF388;
defparam \portb~32 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y35_N0
cycloneive_lcell_comb \wdat[16]~30 (
// Equation(s):
// \wdat[16]~30_combout  = (!plif_memwbregsrc_l_1 & ((plif_memwbregsrc_l_0 & ((plif_memwbdmemload_l_16))) # (!plif_memwbregsrc_l_0 & (plif_memwbporto_l_16))))

	.dataa(\MEMWB|plif_memwb.regsrc_l [0]),
	.datab(\MEMWB|plif_memwb.porto_l [16]),
	.datac(\MEMWB|plif_memwb.dmemload_l [16]),
	.datad(\MEMWB|plif_memwb.regsrc_l [1]),
	.cin(gnd),
	.combout(\wdat[16]~30_combout ),
	.cout());
// synopsys translate_off
defparam \wdat[16]~30 .lut_mask = 16'h00E4;
defparam \wdat[16]~30 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y35_N26
cycloneive_lcell_comb \wdat[16]~31 (
// Equation(s):
// \wdat[16]~31_combout  = (\wdat[16]~30_combout ) # ((plif_memwbregsrc_l_1 & plif_memwbrtnaddr_l_16))

	.dataa(gnd),
	.datab(\MEMWB|plif_memwb.regsrc_l [1]),
	.datac(\MEMWB|plif_memwb.rtnaddr_l [16]),
	.datad(\wdat[16]~30_combout ),
	.cin(gnd),
	.combout(\wdat[16]~31_combout ),
	.cout());
// synopsys translate_off
defparam \wdat[16]~31 .lut_mask = 16'hFFC0;
defparam \wdat[16]~31 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y35_N24
cycloneive_lcell_comb \portb~33 (
// Equation(s):
// \portb~33_combout  = (\portb~2_combout  & (((\portb~1_combout )))) # (!\portb~2_combout  & ((\portb~1_combout  & ((plif_idexextimm_l_16))) # (!\portb~1_combout  & (plif_idexrdat2_l_16))))

	.dataa(\IDEX|plif_idex.rdat2_l [16]),
	.datab(\IDEX|plif_idex.extimm_l [16]),
	.datac(\portb~2_combout ),
	.datad(\portb~1_combout ),
	.cin(gnd),
	.combout(\portb~33_combout ),
	.cout());
// synopsys translate_off
defparam \portb~33 .lut_mask = 16'hFC0A;
defparam \portb~33 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y35_N10
cycloneive_lcell_comb \portb~34 (
// Equation(s):
// \portb~34_combout  = (\portb~2_combout  & ((\portb~33_combout  & ((plif_exmemporto_l_16))) # (!\portb~33_combout  & (\wdat[16]~31_combout )))) # (!\portb~2_combout  & (((\portb~33_combout ))))

	.dataa(\wdat[16]~31_combout ),
	.datab(plif_exmemporto_l_16),
	.datac(\portb~2_combout ),
	.datad(\portb~33_combout ),
	.cin(gnd),
	.combout(\portb~34_combout ),
	.cout());
// synopsys translate_off
defparam \portb~34 .lut_mask = 16'hCFA0;
defparam \portb~34 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y38_N24
cycloneive_lcell_comb \wdat[15]~32 (
// Equation(s):
// \wdat[15]~32_combout  = (!plif_memwbregsrc_l_1 & ((plif_memwbregsrc_l_0 & (plif_memwbdmemload_l_15)) # (!plif_memwbregsrc_l_0 & ((plif_memwbporto_l_15)))))

	.dataa(\MEMWB|plif_memwb.regsrc_l [1]),
	.datab(\MEMWB|plif_memwb.regsrc_l [0]),
	.datac(\MEMWB|plif_memwb.dmemload_l [15]),
	.datad(\MEMWB|plif_memwb.porto_l [15]),
	.cin(gnd),
	.combout(\wdat[15]~32_combout ),
	.cout());
// synopsys translate_off
defparam \wdat[15]~32 .lut_mask = 16'h5140;
defparam \wdat[15]~32 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y38_N2
cycloneive_lcell_comb \wdat[15]~33 (
// Equation(s):
// \wdat[15]~33_combout  = (\wdat[15]~32_combout ) # ((plif_memwbregsrc_l_1 & plif_memwbrtnaddr_l_15))

	.dataa(\MEMWB|plif_memwb.regsrc_l [1]),
	.datab(gnd),
	.datac(\MEMWB|plif_memwb.rtnaddr_l [15]),
	.datad(\wdat[15]~32_combout ),
	.cin(gnd),
	.combout(\wdat[15]~33_combout ),
	.cout());
// synopsys translate_off
defparam \wdat[15]~33 .lut_mask = 16'hFFA0;
defparam \wdat[15]~33 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y38_N16
cycloneive_lcell_comb \portb~35 (
// Equation(s):
// \portb~35_combout  = (\portb~1_combout  & (((\portb~2_combout )))) # (!\portb~1_combout  & ((\portb~2_combout  & ((\wdat[15]~33_combout ))) # (!\portb~2_combout  & (plif_idexrdat2_l_15))))

	.dataa(\IDEX|plif_idex.rdat2_l [15]),
	.datab(\wdat[15]~33_combout ),
	.datac(\portb~1_combout ),
	.datad(\portb~2_combout ),
	.cin(gnd),
	.combout(\portb~35_combout ),
	.cout());
// synopsys translate_off
defparam \portb~35 .lut_mask = 16'hFC0A;
defparam \portb~35 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y38_N14
cycloneive_lcell_comb \portb~36 (
// Equation(s):
// \portb~36_combout  = (\portb~1_combout  & ((\portb~35_combout  & (plif_exmemporto_l_15)) # (!\portb~35_combout  & ((plif_idexextimm_l_15))))) # (!\portb~1_combout  & (((\portb~35_combout ))))

	.dataa(\portb~1_combout ),
	.datab(plif_exmemporto_l_15),
	.datac(\IDEX|plif_idex.extimm_l [15]),
	.datad(\portb~35_combout ),
	.cin(gnd),
	.combout(\portb~36_combout ),
	.cout());
// synopsys translate_off
defparam \portb~36 .lut_mask = 16'hDDA0;
defparam \portb~36 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y35_N2
cycloneive_lcell_comb \wdat[14]~34 (
// Equation(s):
// \wdat[14]~34_combout  = (!plif_memwbregsrc_l_1 & ((plif_memwbregsrc_l_0 & ((plif_memwbdmemload_l_14))) # (!plif_memwbregsrc_l_0 & (plif_memwbporto_l_14))))

	.dataa(\MEMWB|plif_memwb.regsrc_l [1]),
	.datab(\MEMWB|plif_memwb.porto_l [14]),
	.datac(\MEMWB|plif_memwb.dmemload_l [14]),
	.datad(\MEMWB|plif_memwb.regsrc_l [0]),
	.cin(gnd),
	.combout(\wdat[14]~34_combout ),
	.cout());
// synopsys translate_off
defparam \wdat[14]~34 .lut_mask = 16'h5044;
defparam \wdat[14]~34 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y35_N4
cycloneive_lcell_comb \wdat[14]~35 (
// Equation(s):
// \wdat[14]~35_combout  = (\wdat[14]~34_combout ) # ((plif_memwbrtnaddr_l_14 & plif_memwbregsrc_l_1))

	.dataa(\MEMWB|plif_memwb.rtnaddr_l [14]),
	.datab(\MEMWB|plif_memwb.regsrc_l [1]),
	.datac(gnd),
	.datad(\wdat[14]~34_combout ),
	.cin(gnd),
	.combout(\wdat[14]~35_combout ),
	.cout());
// synopsys translate_off
defparam \wdat[14]~35 .lut_mask = 16'hFF88;
defparam \wdat[14]~35 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y38_N4
cycloneive_lcell_comb \portb~37 (
// Equation(s):
// \portb~37_combout  = (\portb~1_combout  & ((\portb~2_combout  & (plif_exmemporto_l_14)) # (!\portb~2_combout  & ((plif_idexextimm_l_14))))) # (!\portb~1_combout  & (((\portb~2_combout ))))

	.dataa(plif_exmemporto_l_14),
	.datab(\IDEX|plif_idex.extimm_l [14]),
	.datac(\portb~1_combout ),
	.datad(\portb~2_combout ),
	.cin(gnd),
	.combout(\portb~37_combout ),
	.cout());
// synopsys translate_off
defparam \portb~37 .lut_mask = 16'hAFC0;
defparam \portb~37 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y38_N26
cycloneive_lcell_comb \portb~38 (
// Equation(s):
// \portb~38_combout  = (\portb~1_combout  & (\portb~37_combout )) # (!\portb~1_combout  & ((\portb~37_combout  & (\wdat[14]~35_combout )) # (!\portb~37_combout  & ((plif_idexrdat2_l_14)))))

	.dataa(\portb~1_combout ),
	.datab(\portb~37_combout ),
	.datac(\wdat[14]~35_combout ),
	.datad(\IDEX|plif_idex.rdat2_l [14]),
	.cin(gnd),
	.combout(\portb~38_combout ),
	.cout());
// synopsys translate_off
defparam \portb~38 .lut_mask = 16'hD9C8;
defparam \portb~38 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y38_N0
cycloneive_lcell_comb \wdat[13]~36 (
// Equation(s):
// \wdat[13]~36_combout  = (!plif_memwbregsrc_l_1 & ((plif_memwbregsrc_l_0 & ((plif_memwbdmemload_l_13))) # (!plif_memwbregsrc_l_0 & (plif_memwbporto_l_13))))

	.dataa(\MEMWB|plif_memwb.regsrc_l [1]),
	.datab(\MEMWB|plif_memwb.porto_l [13]),
	.datac(\MEMWB|plif_memwb.dmemload_l [13]),
	.datad(\MEMWB|plif_memwb.regsrc_l [0]),
	.cin(gnd),
	.combout(\wdat[13]~36_combout ),
	.cout());
// synopsys translate_off
defparam \wdat[13]~36 .lut_mask = 16'h5044;
defparam \wdat[13]~36 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y38_N8
cycloneive_lcell_comb \wdat[13]~37 (
// Equation(s):
// \wdat[13]~37_combout  = (\wdat[13]~36_combout ) # ((plif_memwbregsrc_l_1 & plif_memwbrtnaddr_l_13))

	.dataa(\MEMWB|plif_memwb.regsrc_l [1]),
	.datab(gnd),
	.datac(\MEMWB|plif_memwb.rtnaddr_l [13]),
	.datad(\wdat[13]~36_combout ),
	.cin(gnd),
	.combout(\wdat[13]~37_combout ),
	.cout());
// synopsys translate_off
defparam \wdat[13]~37 .lut_mask = 16'hFFA0;
defparam \wdat[13]~37 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y38_N20
cycloneive_lcell_comb \portb~39 (
// Equation(s):
// \portb~39_combout  = (\portb~1_combout  & (((\portb~2_combout )))) # (!\portb~1_combout  & ((\portb~2_combout  & ((\wdat[13]~37_combout ))) # (!\portb~2_combout  & (plif_idexrdat2_l_13))))

	.dataa(\IDEX|plif_idex.rdat2_l [13]),
	.datab(\wdat[13]~37_combout ),
	.datac(\portb~1_combout ),
	.datad(\portb~2_combout ),
	.cin(gnd),
	.combout(\portb~39_combout ),
	.cout());
// synopsys translate_off
defparam \portb~39 .lut_mask = 16'hFC0A;
defparam \portb~39 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y38_N6
cycloneive_lcell_comb \portb~40 (
// Equation(s):
// \portb~40_combout  = (\portb~1_combout  & ((\portb~39_combout  & ((plif_exmemporto_l_13))) # (!\portb~39_combout  & (plif_idexextimm_l_13)))) # (!\portb~1_combout  & (((\portb~39_combout ))))

	.dataa(\portb~1_combout ),
	.datab(\IDEX|plif_idex.extimm_l [13]),
	.datac(plif_exmemporto_l_13),
	.datad(\portb~39_combout ),
	.cin(gnd),
	.combout(\portb~40_combout ),
	.cout());
// synopsys translate_off
defparam \portb~40 .lut_mask = 16'hF588;
defparam \portb~40 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y34_N26
cycloneive_lcell_comb \wdat[12]~38 (
// Equation(s):
// \wdat[12]~38_combout  = (!plif_memwbregsrc_l_1 & ((plif_memwbregsrc_l_0 & ((plif_memwbdmemload_l_12))) # (!plif_memwbregsrc_l_0 & (plif_memwbporto_l_12))))

	.dataa(\MEMWB|plif_memwb.porto_l [12]),
	.datab(\MEMWB|plif_memwb.regsrc_l [1]),
	.datac(\MEMWB|plif_memwb.dmemload_l [12]),
	.datad(\MEMWB|plif_memwb.regsrc_l [0]),
	.cin(gnd),
	.combout(\wdat[12]~38_combout ),
	.cout());
// synopsys translate_off
defparam \wdat[12]~38 .lut_mask = 16'h3022;
defparam \wdat[12]~38 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y34_N2
cycloneive_lcell_comb \wdat[12]~39 (
// Equation(s):
// \wdat[12]~39_combout  = (\wdat[12]~38_combout ) # ((plif_memwbregsrc_l_1 & plif_memwbrtnaddr_l_12))

	.dataa(\wdat[12]~38_combout ),
	.datab(\MEMWB|plif_memwb.regsrc_l [1]),
	.datac(\MEMWB|plif_memwb.rtnaddr_l [12]),
	.datad(gnd),
	.cin(gnd),
	.combout(\wdat[12]~39_combout ),
	.cout());
// synopsys translate_off
defparam \wdat[12]~39 .lut_mask = 16'hEAEA;
defparam \wdat[12]~39 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y38_N30
cycloneive_lcell_comb \portb~41 (
// Equation(s):
// \portb~41_combout  = (\portb~1_combout  & ((\portb~2_combout  & ((plif_exmemporto_l_12))) # (!\portb~2_combout  & (plif_idexextimm_l_12)))) # (!\portb~1_combout  & (((\portb~2_combout ))))

	.dataa(\IDEX|plif_idex.extimm_l [12]),
	.datab(plif_exmemporto_l_12),
	.datac(\portb~1_combout ),
	.datad(\portb~2_combout ),
	.cin(gnd),
	.combout(\portb~41_combout ),
	.cout());
// synopsys translate_off
defparam \portb~41 .lut_mask = 16'hCFA0;
defparam \portb~41 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y38_N12
cycloneive_lcell_comb \portb~42 (
// Equation(s):
// \portb~42_combout  = (\portb~41_combout  & (((\portb~1_combout ) # (\wdat[12]~39_combout )))) # (!\portb~41_combout  & (plif_idexrdat2_l_12 & (!\portb~1_combout )))

	.dataa(\portb~41_combout ),
	.datab(\IDEX|plif_idex.rdat2_l [12]),
	.datac(\portb~1_combout ),
	.datad(\wdat[12]~39_combout ),
	.cin(gnd),
	.combout(\portb~42_combout ),
	.cout());
// synopsys translate_off
defparam \portb~42 .lut_mask = 16'hAEA4;
defparam \portb~42 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y38_N8
cycloneive_lcell_comb \wdat[11]~40 (
// Equation(s):
// \wdat[11]~40_combout  = (!plif_memwbregsrc_l_1 & ((plif_memwbregsrc_l_0 & ((plif_memwbdmemload_l_11))) # (!plif_memwbregsrc_l_0 & (plif_memwbporto_l_11))))

	.dataa(\MEMWB|plif_memwb.porto_l [11]),
	.datab(\MEMWB|plif_memwb.regsrc_l [0]),
	.datac(\MEMWB|plif_memwb.dmemload_l [11]),
	.datad(\MEMWB|plif_memwb.regsrc_l [1]),
	.cin(gnd),
	.combout(\wdat[11]~40_combout ),
	.cout());
// synopsys translate_off
defparam \wdat[11]~40 .lut_mask = 16'h00E2;
defparam \wdat[11]~40 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y38_N4
cycloneive_lcell_comb \wdat[11]~41 (
// Equation(s):
// \wdat[11]~41_combout  = (\wdat[11]~40_combout ) # ((plif_memwbrtnaddr_l_11 & plif_memwbregsrc_l_1))

	.dataa(gnd),
	.datab(\wdat[11]~40_combout ),
	.datac(\MEMWB|plif_memwb.rtnaddr_l [11]),
	.datad(\MEMWB|plif_memwb.regsrc_l [1]),
	.cin(gnd),
	.combout(\wdat[11]~41_combout ),
	.cout());
// synopsys translate_off
defparam \wdat[11]~41 .lut_mask = 16'hFCCC;
defparam \wdat[11]~41 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y38_N0
cycloneive_lcell_comb \portb~43 (
// Equation(s):
// \portb~43_combout  = (\portb~2_combout  & (((\wdat[11]~41_combout ) # (\portb~1_combout )))) # (!\portb~2_combout  & (plif_idexrdat2_l_11 & ((!\portb~1_combout ))))

	.dataa(\IDEX|plif_idex.rdat2_l [11]),
	.datab(\wdat[11]~41_combout ),
	.datac(\portb~2_combout ),
	.datad(\portb~1_combout ),
	.cin(gnd),
	.combout(\portb~43_combout ),
	.cout());
// synopsys translate_off
defparam \portb~43 .lut_mask = 16'hF0CA;
defparam \portb~43 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y38_N26
cycloneive_lcell_comb \portb~44 (
// Equation(s):
// \portb~44_combout  = (\portb~1_combout  & ((\portb~43_combout  & (plif_exmemporto_l_11)) # (!\portb~43_combout  & ((plif_idexextimm_l_11))))) # (!\portb~1_combout  & (\portb~43_combout ))

	.dataa(\portb~1_combout ),
	.datab(\portb~43_combout ),
	.datac(plif_exmemporto_l_11),
	.datad(\IDEX|plif_idex.extimm_l [11]),
	.cin(gnd),
	.combout(\portb~44_combout ),
	.cout());
// synopsys translate_off
defparam \portb~44 .lut_mask = 16'hE6C4;
defparam \portb~44 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y34_N30
cycloneive_lcell_comb \wdat[10]~42 (
// Equation(s):
// \wdat[10]~42_combout  = (!plif_memwbregsrc_l_1 & ((plif_memwbregsrc_l_0 & ((plif_memwbdmemload_l_10))) # (!plif_memwbregsrc_l_0 & (plif_memwbporto_l_10))))

	.dataa(\MEMWB|plif_memwb.regsrc_l [0]),
	.datab(\MEMWB|plif_memwb.porto_l [10]),
	.datac(\MEMWB|plif_memwb.dmemload_l [10]),
	.datad(\MEMWB|plif_memwb.regsrc_l [1]),
	.cin(gnd),
	.combout(\wdat[10]~42_combout ),
	.cout());
// synopsys translate_off
defparam \wdat[10]~42 .lut_mask = 16'h00E4;
defparam \wdat[10]~42 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y34_N18
cycloneive_lcell_comb \wdat[10]~43 (
// Equation(s):
// \wdat[10]~43_combout  = (\wdat[10]~42_combout ) # ((plif_memwbrtnaddr_l_10 & plif_memwbregsrc_l_1))

	.dataa(\wdat[10]~42_combout ),
	.datab(gnd),
	.datac(\MEMWB|plif_memwb.rtnaddr_l [10]),
	.datad(\MEMWB|plif_memwb.regsrc_l [1]),
	.cin(gnd),
	.combout(\wdat[10]~43_combout ),
	.cout());
// synopsys translate_off
defparam \wdat[10]~43 .lut_mask = 16'hFAAA;
defparam \wdat[10]~43 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y38_N20
cycloneive_lcell_comb \portb~45 (
// Equation(s):
// \portb~45_combout  = (\portb~2_combout  & ((plif_exmemporto_l_10) # ((!\portb~1_combout )))) # (!\portb~2_combout  & (((plif_idexextimm_l_10 & \portb~1_combout ))))

	.dataa(plif_exmemporto_l_10),
	.datab(\IDEX|plif_idex.extimm_l [10]),
	.datac(\portb~2_combout ),
	.datad(\portb~1_combout ),
	.cin(gnd),
	.combout(\portb~45_combout ),
	.cout());
// synopsys translate_off
defparam \portb~45 .lut_mask = 16'hACF0;
defparam \portb~45 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y38_N10
cycloneive_lcell_comb \portb~46 (
// Equation(s):
// \portb~46_combout  = (\portb~45_combout  & ((\wdat[10]~43_combout ) # ((\portb~1_combout )))) # (!\portb~45_combout  & (((plif_idexrdat2_l_10 & !\portb~1_combout ))))

	.dataa(\wdat[10]~43_combout ),
	.datab(\portb~45_combout ),
	.datac(\IDEX|plif_idex.rdat2_l [10]),
	.datad(\portb~1_combout ),
	.cin(gnd),
	.combout(\portb~46_combout ),
	.cout());
// synopsys translate_off
defparam \portb~46 .lut_mask = 16'hCCB8;
defparam \portb~46 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y35_N10
cycloneive_lcell_comb \wdat[9]~44 (
// Equation(s):
// \wdat[9]~44_combout  = (!plif_memwbregsrc_l_1 & ((plif_memwbregsrc_l_0 & ((plif_memwbdmemload_l_9))) # (!plif_memwbregsrc_l_0 & (plif_memwbporto_l_9))))

	.dataa(\MEMWB|plif_memwb.porto_l [9]),
	.datab(\MEMWB|plif_memwb.regsrc_l [1]),
	.datac(\MEMWB|plif_memwb.dmemload_l [9]),
	.datad(\MEMWB|plif_memwb.regsrc_l [0]),
	.cin(gnd),
	.combout(\wdat[9]~44_combout ),
	.cout());
// synopsys translate_off
defparam \wdat[9]~44 .lut_mask = 16'h3022;
defparam \wdat[9]~44 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y35_N8
cycloneive_lcell_comb \wdat[9]~45 (
// Equation(s):
// \wdat[9]~45_combout  = (\wdat[9]~44_combout ) # ((plif_memwbregsrc_l_1 & plif_memwbrtnaddr_l_9))

	.dataa(\MEMWB|plif_memwb.regsrc_l [1]),
	.datab(\MEMWB|plif_memwb.rtnaddr_l [9]),
	.datac(gnd),
	.datad(\wdat[9]~44_combout ),
	.cin(gnd),
	.combout(\wdat[9]~45_combout ),
	.cout());
// synopsys translate_off
defparam \wdat[9]~45 .lut_mask = 16'hFF88;
defparam \wdat[9]~45 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y38_N28
cycloneive_lcell_comb \portb~47 (
// Equation(s):
// \portb~47_combout  = (\portb~2_combout  & ((\wdat[9]~45_combout ) # ((\portb~1_combout )))) # (!\portb~2_combout  & (((plif_idexrdat2_l_9 & !\portb~1_combout ))))

	.dataa(\wdat[9]~45_combout ),
	.datab(\IDEX|plif_idex.rdat2_l [9]),
	.datac(\portb~2_combout ),
	.datad(\portb~1_combout ),
	.cin(gnd),
	.combout(\portb~47_combout ),
	.cout());
// synopsys translate_off
defparam \portb~47 .lut_mask = 16'hF0AC;
defparam \portb~47 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y38_N6
cycloneive_lcell_comb \portb~48 (
// Equation(s):
// \portb~48_combout  = (\portb~1_combout  & ((\portb~47_combout  & ((plif_exmemporto_l_9))) # (!\portb~47_combout  & (plif_idexextimm_l_9)))) # (!\portb~1_combout  & (((\portb~47_combout ))))

	.dataa(\portb~1_combout ),
	.datab(\IDEX|plif_idex.extimm_l [9]),
	.datac(plif_exmemporto_l_9),
	.datad(\portb~47_combout ),
	.cin(gnd),
	.combout(\portb~48_combout ),
	.cout());
// synopsys translate_off
defparam \portb~48 .lut_mask = 16'hF588;
defparam \portb~48 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y33_N2
cycloneive_lcell_comb \wdat[8]~46 (
// Equation(s):
// \wdat[8]~46_combout  = (!plif_memwbregsrc_l_1 & ((plif_memwbregsrc_l_0 & ((plif_memwbdmemload_l_8))) # (!plif_memwbregsrc_l_0 & (plif_memwbporto_l_8))))

	.dataa(\MEMWB|plif_memwb.regsrc_l [1]),
	.datab(\MEMWB|plif_memwb.porto_l [8]),
	.datac(\MEMWB|plif_memwb.dmemload_l [8]),
	.datad(\MEMWB|plif_memwb.regsrc_l [0]),
	.cin(gnd),
	.combout(\wdat[8]~46_combout ),
	.cout());
// synopsys translate_off
defparam \wdat[8]~46 .lut_mask = 16'h5044;
defparam \wdat[8]~46 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y33_N22
cycloneive_lcell_comb \wdat[8]~47 (
// Equation(s):
// \wdat[8]~47_combout  = (\wdat[8]~46_combout ) # ((plif_memwbregsrc_l_1 & plif_memwbrtnaddr_l_8))

	.dataa(\MEMWB|plif_memwb.regsrc_l [1]),
	.datab(gnd),
	.datac(\MEMWB|plif_memwb.rtnaddr_l [8]),
	.datad(\wdat[8]~46_combout ),
	.cin(gnd),
	.combout(\wdat[8]~47_combout ),
	.cout());
// synopsys translate_off
defparam \wdat[8]~47 .lut_mask = 16'hFFA0;
defparam \wdat[8]~47 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y38_N12
cycloneive_lcell_comb \portb~49 (
// Equation(s):
// \portb~49_combout  = (\portb~2_combout  & ((plif_exmemporto_l_8) # ((!\portb~1_combout )))) # (!\portb~2_combout  & (((plif_idexextimm_l_8 & \portb~1_combout ))))

	.dataa(plif_exmemporto_l_8),
	.datab(\IDEX|plif_idex.extimm_l [8]),
	.datac(\portb~2_combout ),
	.datad(\portb~1_combout ),
	.cin(gnd),
	.combout(\portb~49_combout ),
	.cout());
// synopsys translate_off
defparam \portb~49 .lut_mask = 16'hACF0;
defparam \portb~49 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y38_N14
cycloneive_lcell_comb \portb~50 (
// Equation(s):
// \portb~50_combout  = (\portb~1_combout  & (((\portb~49_combout )))) # (!\portb~1_combout  & ((\portb~49_combout  & ((\wdat[8]~47_combout ))) # (!\portb~49_combout  & (plif_idexrdat2_l_8))))

	.dataa(\portb~1_combout ),
	.datab(\IDEX|plif_idex.rdat2_l [8]),
	.datac(\wdat[8]~47_combout ),
	.datad(\portb~49_combout ),
	.cin(gnd),
	.combout(\portb~50_combout ),
	.cout());
// synopsys translate_off
defparam \portb~50 .lut_mask = 16'hFA44;
defparam \portb~50 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y38_N0
cycloneive_lcell_comb \wdat[7]~48 (
// Equation(s):
// \wdat[7]~48_combout  = (!plif_memwbregsrc_l_1 & ((plif_memwbregsrc_l_0 & ((plif_memwbdmemload_l_7))) # (!plif_memwbregsrc_l_0 & (plif_memwbporto_l_7))))

	.dataa(\MEMWB|plif_memwb.regsrc_l [1]),
	.datab(\MEMWB|plif_memwb.porto_l [7]),
	.datac(\MEMWB|plif_memwb.dmemload_l [7]),
	.datad(\MEMWB|plif_memwb.regsrc_l [0]),
	.cin(gnd),
	.combout(\wdat[7]~48_combout ),
	.cout());
// synopsys translate_off
defparam \wdat[7]~48 .lut_mask = 16'h5044;
defparam \wdat[7]~48 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y38_N16
cycloneive_lcell_comb \wdat[7]~49 (
// Equation(s):
// \wdat[7]~49_combout  = (\wdat[7]~48_combout ) # ((plif_memwbregsrc_l_1 & plif_memwbrtnaddr_l_7))

	.dataa(\MEMWB|plif_memwb.regsrc_l [1]),
	.datab(gnd),
	.datac(\MEMWB|plif_memwb.rtnaddr_l [7]),
	.datad(\wdat[7]~48_combout ),
	.cin(gnd),
	.combout(\wdat[7]~49_combout ),
	.cout());
// synopsys translate_off
defparam \wdat[7]~49 .lut_mask = 16'hFFA0;
defparam \wdat[7]~49 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y38_N24
cycloneive_lcell_comb \portb~51 (
// Equation(s):
// \portb~51_combout  = (\portb~1_combout  & (((\portb~2_combout )))) # (!\portb~1_combout  & ((\portb~2_combout  & ((\wdat[7]~49_combout ))) # (!\portb~2_combout  & (plif_idexrdat2_l_7))))

	.dataa(\IDEX|plif_idex.rdat2_l [7]),
	.datab(\portb~1_combout ),
	.datac(\portb~2_combout ),
	.datad(\wdat[7]~49_combout ),
	.cin(gnd),
	.combout(\portb~51_combout ),
	.cout());
// synopsys translate_off
defparam \portb~51 .lut_mask = 16'hF2C2;
defparam \portb~51 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y38_N6
cycloneive_lcell_comb \portb~52 (
// Equation(s):
// \portb~52_combout  = (\portb~1_combout  & ((\portb~51_combout  & ((plif_exmemporto_l_7))) # (!\portb~51_combout  & (plif_idexextimm_l_7)))) # (!\portb~1_combout  & (((\portb~51_combout ))))

	.dataa(\IDEX|plif_idex.extimm_l [7]),
	.datab(\portb~1_combout ),
	.datac(plif_exmemporto_l_7),
	.datad(\portb~51_combout ),
	.cin(gnd),
	.combout(\portb~52_combout ),
	.cout());
// synopsys translate_off
defparam \portb~52 .lut_mask = 16'hF388;
defparam \portb~52 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y39_N16
cycloneive_lcell_comb \wdat[6]~50 (
// Equation(s):
// \wdat[6]~50_combout  = (!plif_memwbregsrc_l_1 & ((plif_memwbregsrc_l_0 & ((plif_memwbdmemload_l_6))) # (!plif_memwbregsrc_l_0 & (plif_memwbporto_l_6))))

	.dataa(\MEMWB|plif_memwb.regsrc_l [1]),
	.datab(\MEMWB|plif_memwb.porto_l [6]),
	.datac(\MEMWB|plif_memwb.dmemload_l [6]),
	.datad(\MEMWB|plif_memwb.regsrc_l [0]),
	.cin(gnd),
	.combout(\wdat[6]~50_combout ),
	.cout());
// synopsys translate_off
defparam \wdat[6]~50 .lut_mask = 16'h5044;
defparam \wdat[6]~50 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y39_N30
cycloneive_lcell_comb \wdat[6]~51 (
// Equation(s):
// \wdat[6]~51_combout  = (\wdat[6]~50_combout ) # ((plif_memwbregsrc_l_1 & plif_memwbrtnaddr_l_6))

	.dataa(\MEMWB|plif_memwb.regsrc_l [1]),
	.datab(gnd),
	.datac(\MEMWB|plif_memwb.rtnaddr_l [6]),
	.datad(\wdat[6]~50_combout ),
	.cin(gnd),
	.combout(\wdat[6]~51_combout ),
	.cout());
// synopsys translate_off
defparam \wdat[6]~51 .lut_mask = 16'hFFA0;
defparam \wdat[6]~51 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y38_N20
cycloneive_lcell_comb \portb~53 (
// Equation(s):
// \portb~53_combout  = (\portb~2_combout  & (((plif_exmemporto_l_6) # (!\portb~1_combout )))) # (!\portb~2_combout  & (plif_idexextimm_l_6 & ((\portb~1_combout ))))

	.dataa(\IDEX|plif_idex.extimm_l [6]),
	.datab(plif_exmemporto_l_6),
	.datac(\portb~2_combout ),
	.datad(\portb~1_combout ),
	.cin(gnd),
	.combout(\portb~53_combout ),
	.cout());
// synopsys translate_off
defparam \portb~53 .lut_mask = 16'hCAF0;
defparam \portb~53 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y38_N26
cycloneive_lcell_comb \portb~54 (
// Equation(s):
// \portb~54_combout  = (\portb~1_combout  & (((\portb~53_combout )))) # (!\portb~1_combout  & ((\portb~53_combout  & ((\wdat[6]~51_combout ))) # (!\portb~53_combout  & (plif_idexrdat2_l_6))))

	.dataa(\IDEX|plif_idex.rdat2_l [6]),
	.datab(\portb~1_combout ),
	.datac(\wdat[6]~51_combout ),
	.datad(\portb~53_combout ),
	.cin(gnd),
	.combout(\portb~54_combout ),
	.cout());
// synopsys translate_off
defparam \portb~54 .lut_mask = 16'hFC22;
defparam \portb~54 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y38_N8
cycloneive_lcell_comb \wdat[5]~52 (
// Equation(s):
// \wdat[5]~52_combout  = (!plif_memwbregsrc_l_1 & ((plif_memwbregsrc_l_0 & (plif_memwbdmemload_l_5)) # (!plif_memwbregsrc_l_0 & ((plif_memwbporto_l_5)))))

	.dataa(\MEMWB|plif_memwb.regsrc_l [1]),
	.datab(\MEMWB|plif_memwb.regsrc_l [0]),
	.datac(\MEMWB|plif_memwb.dmemload_l [5]),
	.datad(\MEMWB|plif_memwb.porto_l [5]),
	.cin(gnd),
	.combout(\wdat[5]~52_combout ),
	.cout());
// synopsys translate_off
defparam \wdat[5]~52 .lut_mask = 16'h5140;
defparam \wdat[5]~52 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y38_N28
cycloneive_lcell_comb \wdat[5]~53 (
// Equation(s):
// \wdat[5]~53_combout  = (\wdat[5]~52_combout ) # ((plif_memwbregsrc_l_1 & plif_memwbrtnaddr_l_5))

	.dataa(\MEMWB|plif_memwb.regsrc_l [1]),
	.datab(\wdat[5]~52_combout ),
	.datac(\MEMWB|plif_memwb.rtnaddr_l [5]),
	.datad(gnd),
	.cin(gnd),
	.combout(\wdat[5]~53_combout ),
	.cout());
// synopsys translate_off
defparam \wdat[5]~53 .lut_mask = 16'hECEC;
defparam \wdat[5]~53 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y38_N18
cycloneive_lcell_comb \portb~55 (
// Equation(s):
// \portb~55_combout  = (\portb~1_combout  & (((\portb~2_combout )))) # (!\portb~1_combout  & ((\portb~2_combout  & (\wdat[5]~53_combout )) # (!\portb~2_combout  & ((plif_idexrdat2_l_5)))))

	.dataa(\wdat[5]~53_combout ),
	.datab(\portb~1_combout ),
	.datac(\portb~2_combout ),
	.datad(\IDEX|plif_idex.rdat2_l [5]),
	.cin(gnd),
	.combout(\portb~55_combout ),
	.cout());
// synopsys translate_off
defparam \portb~55 .lut_mask = 16'hE3E0;
defparam \portb~55 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y38_N4
cycloneive_lcell_comb \portb~56 (
// Equation(s):
// \portb~56_combout  = (\portb~1_combout  & ((\portb~55_combout  & ((plif_exmemporto_l_5))) # (!\portb~55_combout  & (plif_idexextimm_l_5)))) # (!\portb~1_combout  & (((\portb~55_combout ))))

	.dataa(\IDEX|plif_idex.extimm_l [5]),
	.datab(\portb~1_combout ),
	.datac(plif_exmemporto_l_5),
	.datad(\portb~55_combout ),
	.cin(gnd),
	.combout(\portb~56_combout ),
	.cout());
// synopsys translate_off
defparam \portb~56 .lut_mask = 16'hF388;
defparam \portb~56 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y35_N6
cycloneive_lcell_comb \wdat[2]~54 (
// Equation(s):
// \wdat[2]~54_combout  = (!plif_memwbregsrc_l_1 & ((plif_memwbregsrc_l_0 & ((plif_memwbdmemload_l_2))) # (!plif_memwbregsrc_l_0 & (plif_memwbporto_l_2))))

	.dataa(\MEMWB|plif_memwb.regsrc_l [1]),
	.datab(\MEMWB|plif_memwb.porto_l [2]),
	.datac(\MEMWB|plif_memwb.dmemload_l [2]),
	.datad(\MEMWB|plif_memwb.regsrc_l [0]),
	.cin(gnd),
	.combout(\wdat[2]~54_combout ),
	.cout());
// synopsys translate_off
defparam \wdat[2]~54 .lut_mask = 16'h5044;
defparam \wdat[2]~54 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y39_N8
cycloneive_lcell_comb \wdat[2]~55 (
// Equation(s):
// \wdat[2]~55_combout  = (\wdat[2]~54_combout ) # ((plif_memwbregsrc_l_1 & plif_memwbrtnaddr_l_2))

	.dataa(\MEMWB|plif_memwb.regsrc_l [1]),
	.datab(\MEMWB|plif_memwb.rtnaddr_l [2]),
	.datac(gnd),
	.datad(\wdat[2]~54_combout ),
	.cin(gnd),
	.combout(\wdat[2]~55_combout ),
	.cout());
// synopsys translate_off
defparam \wdat[2]~55 .lut_mask = 16'hFF88;
defparam \wdat[2]~55 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y39_N20
cycloneive_lcell_comb \porta~54 (
// Equation(s):
// \porta~54_combout  = (always03 & (((plif_exmemporto_l_2)))) # (!always03 & (fwda & ((\wdat[2]~55_combout ))))

	.dataa(\FU|fwda~3_combout ),
	.datab(plif_exmemporto_l_2),
	.datac(\wdat[2]~55_combout ),
	.datad(\FU|always0~8_combout ),
	.cin(gnd),
	.combout(\porta~54_combout ),
	.cout());
// synopsys translate_off
defparam \porta~54 .lut_mask = 16'hCCA0;
defparam \porta~54 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y39_N18
cycloneive_lcell_comb \porta~55 (
// Equation(s):
// \porta~55_combout  = (\porta~54_combout ) # ((!fwda & (!always03 & plif_idexrdat1_l_2)))

	.dataa(\FU|fwda~3_combout ),
	.datab(\FU|always0~8_combout ),
	.datac(\IDEX|plif_idex.rdat1_l [2]),
	.datad(\porta~54_combout ),
	.cin(gnd),
	.combout(\porta~55_combout ),
	.cout());
// synopsys translate_off
defparam \porta~55 .lut_mask = 16'hFF10;
defparam \porta~55 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y34_N0
cycloneive_lcell_comb \wdat[1]~56 (
// Equation(s):
// \wdat[1]~56_combout  = (!plif_memwbregsrc_l_1 & ((plif_memwbregsrc_l_0 & ((plif_memwbdmemload_l_1))) # (!plif_memwbregsrc_l_0 & (plif_memwbporto_l_1))))

	.dataa(\MEMWB|plif_memwb.porto_l [1]),
	.datab(\MEMWB|plif_memwb.regsrc_l [1]),
	.datac(\MEMWB|plif_memwb.dmemload_l [1]),
	.datad(\MEMWB|plif_memwb.regsrc_l [0]),
	.cin(gnd),
	.combout(\wdat[1]~56_combout ),
	.cout());
// synopsys translate_off
defparam \wdat[1]~56 .lut_mask = 16'h3022;
defparam \wdat[1]~56 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y34_N6
cycloneive_lcell_comb \wdat[1]~57 (
// Equation(s):
// \wdat[1]~57_combout  = (\wdat[1]~56_combout ) # ((plif_memwbregsrc_l_1 & plif_memwbrtnaddr_l_1))

	.dataa(gnd),
	.datab(\MEMWB|plif_memwb.regsrc_l [1]),
	.datac(\MEMWB|plif_memwb.rtnaddr_l [1]),
	.datad(\wdat[1]~56_combout ),
	.cin(gnd),
	.combout(\wdat[1]~57_combout ),
	.cout());
// synopsys translate_off
defparam \wdat[1]~57 .lut_mask = 16'hFFC0;
defparam \wdat[1]~57 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y34_N24
cycloneive_lcell_comb \porta~56 (
// Equation(s):
// \porta~56_combout  = (always03 & (plif_exmemporto_l_1)) # (!always03 & (((fwda & \wdat[1]~57_combout ))))

	.dataa(plif_exmemporto_l_1),
	.datab(\FU|fwda~3_combout ),
	.datac(\wdat[1]~57_combout ),
	.datad(\FU|always0~8_combout ),
	.cin(gnd),
	.combout(\porta~56_combout ),
	.cout());
// synopsys translate_off
defparam \porta~56 .lut_mask = 16'hAAC0;
defparam \porta~56 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y34_N10
cycloneive_lcell_comb \porta~57 (
// Equation(s):
// \porta~57_combout  = (\porta~56_combout ) # ((!always03 & (!fwda & plif_idexrdat1_l_1)))

	.dataa(\FU|always0~8_combout ),
	.datab(\FU|fwda~3_combout ),
	.datac(\IDEX|plif_idex.rdat1_l [1]),
	.datad(\porta~56_combout ),
	.cin(gnd),
	.combout(\porta~57_combout ),
	.cout());
// synopsys translate_off
defparam \porta~57 .lut_mask = 16'hFF10;
defparam \porta~57 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y33_N16
cycloneive_lcell_comb \wdat[0]~58 (
// Equation(s):
// \wdat[0]~58_combout  = (!plif_memwbregsrc_l_1 & ((plif_memwbregsrc_l_0 & ((plif_memwbdmemload_l_0))) # (!plif_memwbregsrc_l_0 & (plif_memwbporto_l_0))))

	.dataa(\MEMWB|plif_memwb.porto_l [0]),
	.datab(\MEMWB|plif_memwb.regsrc_l [1]),
	.datac(\MEMWB|plif_memwb.dmemload_l [0]),
	.datad(\MEMWB|plif_memwb.regsrc_l [0]),
	.cin(gnd),
	.combout(\wdat[0]~58_combout ),
	.cout());
// synopsys translate_off
defparam \wdat[0]~58 .lut_mask = 16'h3022;
defparam \wdat[0]~58 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y33_N10
cycloneive_lcell_comb \wdat[0]~59 (
// Equation(s):
// \wdat[0]~59_combout  = (\wdat[0]~58_combout ) # ((plif_memwbregsrc_l_1 & plif_memwbrtnaddr_l_0))

	.dataa(\MEMWB|plif_memwb.regsrc_l [1]),
	.datab(\MEMWB|plif_memwb.rtnaddr_l [0]),
	.datac(gnd),
	.datad(\wdat[0]~58_combout ),
	.cin(gnd),
	.combout(\wdat[0]~59_combout ),
	.cout());
// synopsys translate_off
defparam \wdat[0]~59 .lut_mask = 16'hFF88;
defparam \wdat[0]~59 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y37_N20
cycloneive_lcell_comb \portb~57 (
// Equation(s):
// \portb~57_combout  = (\portb~2_combout  & ((plif_exmemporto_l_0) # ((!\portb~1_combout )))) # (!\portb~2_combout  & (((plif_idexextimm_l_0 & \portb~1_combout ))))

	.dataa(plif_exmemporto_l_0),
	.datab(\portb~2_combout ),
	.datac(\IDEX|plif_idex.extimm_l [0]),
	.datad(\portb~1_combout ),
	.cin(gnd),
	.combout(\portb~57_combout ),
	.cout());
// synopsys translate_off
defparam \portb~57 .lut_mask = 16'hB8CC;
defparam \portb~57 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y37_N6
cycloneive_lcell_comb \portb~58 (
// Equation(s):
// \portb~58_combout  = (\portb~1_combout  & (((\portb~57_combout )))) # (!\portb~1_combout  & ((\portb~57_combout  & ((\wdat[0]~59_combout ))) # (!\portb~57_combout  & (plif_idexrdat2_l_0))))

	.dataa(\IDEX|plif_idex.rdat2_l [0]),
	.datab(\portb~1_combout ),
	.datac(\wdat[0]~59_combout ),
	.datad(\portb~57_combout ),
	.cin(gnd),
	.combout(\portb~58_combout ),
	.cout());
// synopsys translate_off
defparam \portb~58 .lut_mask = 16'hFC22;
defparam \portb~58 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y39_N28
cycloneive_lcell_comb \portb~59 (
// Equation(s):
// \portb~59_combout  = (\portb~1_combout  & (((\portb~2_combout )))) # (!\portb~1_combout  & ((\portb~2_combout  & ((\wdat[1]~57_combout ))) # (!\portb~2_combout  & (plif_idexrdat2_l_1))))

	.dataa(\portb~1_combout ),
	.datab(\IDEX|plif_idex.rdat2_l [1]),
	.datac(\wdat[1]~57_combout ),
	.datad(\portb~2_combout ),
	.cin(gnd),
	.combout(\portb~59_combout ),
	.cout());
// synopsys translate_off
defparam \portb~59 .lut_mask = 16'hFA44;
defparam \portb~59 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y39_N30
cycloneive_lcell_comb \portb~60 (
// Equation(s):
// \portb~60_combout  = (\portb~1_combout  & ((\portb~59_combout  & (plif_exmemporto_l_1)) # (!\portb~59_combout  & ((plif_idexextimm_l_1))))) # (!\portb~1_combout  & (((\portb~59_combout ))))

	.dataa(plif_exmemporto_l_1),
	.datab(\IDEX|plif_idex.extimm_l [1]),
	.datac(\portb~1_combout ),
	.datad(\portb~59_combout ),
	.cin(gnd),
	.combout(\portb~60_combout ),
	.cout());
// synopsys translate_off
defparam \portb~60 .lut_mask = 16'hAFC0;
defparam \portb~60 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y33_N20
cycloneive_lcell_comb \wdat[4]~60 (
// Equation(s):
// \wdat[4]~60_combout  = (!plif_memwbregsrc_l_1 & ((plif_memwbregsrc_l_0 & ((plif_memwbdmemload_l_4))) # (!plif_memwbregsrc_l_0 & (plif_memwbporto_l_4))))

	.dataa(\MEMWB|plif_memwb.porto_l [4]),
	.datab(\MEMWB|plif_memwb.regsrc_l [1]),
	.datac(\MEMWB|plif_memwb.dmemload_l [4]),
	.datad(\MEMWB|plif_memwb.regsrc_l [0]),
	.cin(gnd),
	.combout(\wdat[4]~60_combout ),
	.cout());
// synopsys translate_off
defparam \wdat[4]~60 .lut_mask = 16'h3022;
defparam \wdat[4]~60 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y33_N22
cycloneive_lcell_comb \wdat[4]~61 (
// Equation(s):
// \wdat[4]~61_combout  = (\wdat[4]~60_combout ) # ((plif_memwbregsrc_l_1 & plif_memwbrtnaddr_l_4))

	.dataa(\MEMWB|plif_memwb.regsrc_l [1]),
	.datab(\MEMWB|plif_memwb.rtnaddr_l [4]),
	.datac(gnd),
	.datad(\wdat[4]~60_combout ),
	.cin(gnd),
	.combout(\wdat[4]~61_combout ),
	.cout());
// synopsys translate_off
defparam \wdat[4]~61 .lut_mask = 16'hFF88;
defparam \wdat[4]~61 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y39_N6
cycloneive_lcell_comb \porta~58 (
// Equation(s):
// \porta~58_combout  = (fwda & ((\wdat[4]~61_combout ))) # (!fwda & (plif_idexrdat1_l_4))

	.dataa(gnd),
	.datab(\IDEX|plif_idex.rdat1_l [4]),
	.datac(\wdat[4]~61_combout ),
	.datad(\FU|fwda~3_combout ),
	.cin(gnd),
	.combout(\porta~58_combout ),
	.cout());
// synopsys translate_off
defparam \porta~58 .lut_mask = 16'hF0CC;
defparam \porta~58 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y39_N0
cycloneive_lcell_comb \porta~59 (
// Equation(s):
// \porta~59_combout  = (always03 & (plif_exmemporto_l_4)) # (!always03 & ((\porta~58_combout )))

	.dataa(gnd),
	.datab(\FU|always0~8_combout ),
	.datac(plif_exmemporto_l_4),
	.datad(\porta~58_combout ),
	.cin(gnd),
	.combout(\porta~59_combout ),
	.cout());
// synopsys translate_off
defparam \porta~59 .lut_mask = 16'hF3C0;
defparam \porta~59 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y35_N24
cycloneive_lcell_comb \wdat[3]~62 (
// Equation(s):
// \wdat[3]~62_combout  = (!plif_memwbregsrc_l_1 & ((plif_memwbregsrc_l_0 & (plif_memwbdmemload_l_3)) # (!plif_memwbregsrc_l_0 & ((plif_memwbporto_l_3)))))

	.dataa(\MEMWB|plif_memwb.regsrc_l [1]),
	.datab(\MEMWB|plif_memwb.regsrc_l [0]),
	.datac(\MEMWB|plif_memwb.dmemload_l [3]),
	.datad(\MEMWB|plif_memwb.porto_l [3]),
	.cin(gnd),
	.combout(\wdat[3]~62_combout ),
	.cout());
// synopsys translate_off
defparam \wdat[3]~62 .lut_mask = 16'h5140;
defparam \wdat[3]~62 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y35_N26
cycloneive_lcell_comb \wdat[3]~63 (
// Equation(s):
// \wdat[3]~63_combout  = (\wdat[3]~62_combout ) # ((plif_memwbrtnaddr_l_3 & plif_memwbregsrc_l_1))

	.dataa(\MEMWB|plif_memwb.rtnaddr_l [3]),
	.datab(\MEMWB|plif_memwb.regsrc_l [1]),
	.datac(gnd),
	.datad(\wdat[3]~62_combout ),
	.cin(gnd),
	.combout(\wdat[3]~63_combout ),
	.cout());
// synopsys translate_off
defparam \wdat[3]~63 .lut_mask = 16'hFF88;
defparam \wdat[3]~63 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y37_N22
cycloneive_lcell_comb \porta~60 (
// Equation(s):
// \porta~60_combout  = (fwda & ((\wdat[3]~63_combout ))) # (!fwda & (plif_idexrdat1_l_3))

	.dataa(gnd),
	.datab(\FU|fwda~3_combout ),
	.datac(\IDEX|plif_idex.rdat1_l [3]),
	.datad(\wdat[3]~63_combout ),
	.cin(gnd),
	.combout(\porta~60_combout ),
	.cout());
// synopsys translate_off
defparam \porta~60 .lut_mask = 16'hFC30;
defparam \porta~60 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y37_N16
cycloneive_lcell_comb \porta~61 (
// Equation(s):
// \porta~61_combout  = (always03 & ((plif_exmemporto_l_3))) # (!always03 & (\porta~60_combout ))

	.dataa(\porta~60_combout ),
	.datab(plif_exmemporto_l_3),
	.datac(gnd),
	.datad(\FU|always0~8_combout ),
	.cin(gnd),
	.combout(\porta~61_combout ),
	.cout());
// synopsys translate_off
defparam \porta~61 .lut_mask = 16'hCCAA;
defparam \porta~61 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y39_N2
cycloneive_lcell_comb \portb~61 (
// Equation(s):
// \portb~61_combout  = (\portb~1_combout  & ((\portb~2_combout  & ((plif_exmemporto_l_2))) # (!\portb~2_combout  & (plif_idexextimm_l_2)))) # (!\portb~1_combout  & (((\portb~2_combout ))))

	.dataa(\IDEX|plif_idex.extimm_l [2]),
	.datab(\portb~1_combout ),
	.datac(plif_exmemporto_l_2),
	.datad(\portb~2_combout ),
	.cin(gnd),
	.combout(\portb~61_combout ),
	.cout());
// synopsys translate_off
defparam \portb~61 .lut_mask = 16'hF388;
defparam \portb~61 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y39_N26
cycloneive_lcell_comb \portb~62 (
// Equation(s):
// \portb~62_combout  = (\portb~1_combout  & (((\portb~61_combout )))) # (!\portb~1_combout  & ((\portb~61_combout  & ((\wdat[2]~55_combout ))) # (!\portb~61_combout  & (plif_idexrdat2_l_2))))

	.dataa(\IDEX|plif_idex.rdat2_l [2]),
	.datab(\portb~1_combout ),
	.datac(\wdat[2]~55_combout ),
	.datad(\portb~61_combout ),
	.cin(gnd),
	.combout(\portb~62_combout ),
	.cout());
// synopsys translate_off
defparam \portb~62 .lut_mask = 16'hFC22;
defparam \portb~62 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y33_N24
cycloneive_lcell_comb \porta~62 (
// Equation(s):
// \porta~62_combout  = (always03 & (((plif_exmemporto_l_8)))) # (!always03 & (\wdat[8]~47_combout  & (fwda)))

	.dataa(\wdat[8]~47_combout ),
	.datab(\FU|fwda~3_combout ),
	.datac(plif_exmemporto_l_8),
	.datad(\FU|always0~8_combout ),
	.cin(gnd),
	.combout(\porta~62_combout ),
	.cout());
// synopsys translate_off
defparam \porta~62 .lut_mask = 16'hF088;
defparam \porta~62 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y36_N10
cycloneive_lcell_comb \porta~63 (
// Equation(s):
// \porta~63_combout  = (fwda) # (always03)

	.dataa(\FU|fwda~3_combout ),
	.datab(gnd),
	.datac(gnd),
	.datad(\FU|always0~8_combout ),
	.cin(gnd),
	.combout(\porta~63_combout ),
	.cout());
// synopsys translate_off
defparam \porta~63 .lut_mask = 16'hFFAA;
defparam \porta~63 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y38_N30
cycloneive_lcell_comb \porta~64 (
// Equation(s):
// \porta~64_combout  = (always03 & (((plif_exmemporto_l_7)))) # (!always03 & ((fwda & (\wdat[7]~49_combout )) # (!fwda & ((plif_exmemporto_l_7)))))

	.dataa(\wdat[7]~49_combout ),
	.datab(\FU|always0~8_combout ),
	.datac(plif_exmemporto_l_7),
	.datad(\FU|fwda~3_combout ),
	.cin(gnd),
	.combout(\porta~64_combout ),
	.cout());
// synopsys translate_off
defparam \porta~64 .lut_mask = 16'hE2F0;
defparam \porta~64 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y39_N28
cycloneive_lcell_comb \porta~65 (
// Equation(s):
// \porta~65_combout  = (always03 & (((plif_exmemporto_l_6)))) # (!always03 & (fwda & ((\wdat[6]~51_combout ))))

	.dataa(\FU|fwda~3_combout ),
	.datab(plif_exmemporto_l_6),
	.datac(\wdat[6]~51_combout ),
	.datad(\FU|always0~8_combout ),
	.cin(gnd),
	.combout(\porta~65_combout ),
	.cout());
// synopsys translate_off
defparam \porta~65 .lut_mask = 16'hCCA0;
defparam \porta~65 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y38_N14
cycloneive_lcell_comb \porta~66 (
// Equation(s):
// \porta~66_combout  = (always03 & (((plif_exmemporto_l_5)))) # (!always03 & (\wdat[5]~53_combout  & ((fwda))))

	.dataa(\wdat[5]~53_combout ),
	.datab(\FU|always0~8_combout ),
	.datac(plif_exmemporto_l_5),
	.datad(\FU|fwda~3_combout ),
	.cin(gnd),
	.combout(\porta~66_combout ),
	.cout());
// synopsys translate_off
defparam \porta~66 .lut_mask = 16'hE2C0;
defparam \porta~66 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y36_N0
cycloneive_lcell_comb \portb~63 (
// Equation(s):
// \portb~63_combout  = (\portb~2_combout  & ((\wdat[3]~63_combout ) # ((\portb~1_combout )))) # (!\portb~2_combout  & (((plif_idexrdat2_l_3 & !\portb~1_combout ))))

	.dataa(\wdat[3]~63_combout ),
	.datab(\IDEX|plif_idex.rdat2_l [3]),
	.datac(\portb~2_combout ),
	.datad(\portb~1_combout ),
	.cin(gnd),
	.combout(\portb~63_combout ),
	.cout());
// synopsys translate_off
defparam \portb~63 .lut_mask = 16'hF0AC;
defparam \portb~63 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y36_N6
cycloneive_lcell_comb \portb~64 (
// Equation(s):
// \portb~64_combout  = (\portb~1_combout  & ((\portb~63_combout  & (plif_exmemporto_l_3)) # (!\portb~63_combout  & ((plif_idexextimm_l_3))))) # (!\portb~1_combout  & (((\portb~63_combout ))))

	.dataa(plif_exmemporto_l_3),
	.datab(\IDEX|plif_idex.extimm_l [3]),
	.datac(\portb~1_combout ),
	.datad(\portb~63_combout ),
	.cin(gnd),
	.combout(\portb~64_combout ),
	.cout());
// synopsys translate_off
defparam \portb~64 .lut_mask = 16'hAFC0;
defparam \portb~64 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y35_N16
cycloneive_lcell_comb \porta~67 (
// Equation(s):
// \porta~67_combout  = (always03 & (((plif_exmemporto_l_16)))) # (!always03 & (\wdat[16]~31_combout  & ((fwda))))

	.dataa(\wdat[16]~31_combout ),
	.datab(plif_exmemporto_l_16),
	.datac(\FU|fwda~3_combout ),
	.datad(\FU|always0~8_combout ),
	.cin(gnd),
	.combout(\porta~67_combout ),
	.cout());
// synopsys translate_off
defparam \porta~67 .lut_mask = 16'hCCA0;
defparam \porta~67 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y40_N0
cycloneive_lcell_comb \porta~68 (
// Equation(s):
// \porta~68_combout  = (always03 & (((plif_exmemporto_l_15)))) # (!always03 & (\wdat[15]~33_combout  & ((fwda))))

	.dataa(\wdat[15]~33_combout ),
	.datab(plif_exmemporto_l_15),
	.datac(\FU|fwda~3_combout ),
	.datad(\FU|always0~8_combout ),
	.cin(gnd),
	.combout(\porta~68_combout ),
	.cout());
// synopsys translate_off
defparam \porta~68 .lut_mask = 16'hCCA0;
defparam \porta~68 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y41_N20
cycloneive_lcell_comb \porta~69 (
// Equation(s):
// \porta~69_combout  = (always03 & (((plif_exmemporto_l_14)))) # (!always03 & (fwda & ((\wdat[14]~35_combout ))))

	.dataa(\FU|always0~8_combout ),
	.datab(\FU|fwda~3_combout ),
	.datac(plif_exmemporto_l_14),
	.datad(\wdat[14]~35_combout ),
	.cin(gnd),
	.combout(\porta~69_combout ),
	.cout());
// synopsys translate_off
defparam \porta~69 .lut_mask = 16'hE4A0;
defparam \porta~69 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y38_N28
cycloneive_lcell_comb \porta~70 (
// Equation(s):
// \porta~70_combout  = (always03 & (plif_exmemporto_l_13)) # (!always03 & (((\wdat[13]~37_combout  & fwda))))

	.dataa(plif_exmemporto_l_13),
	.datab(\wdat[13]~37_combout ),
	.datac(\FU|fwda~3_combout ),
	.datad(\FU|always0~8_combout ),
	.cin(gnd),
	.combout(\porta~70_combout ),
	.cout());
// synopsys translate_off
defparam \porta~70 .lut_mask = 16'hAAC0;
defparam \porta~70 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y34_N20
cycloneive_lcell_comb \porta~71 (
// Equation(s):
// \porta~71_combout  = (always03 & (((plif_exmemporto_l_12)))) # (!always03 & (\wdat[12]~39_combout  & ((fwda))))

	.dataa(\FU|always0~8_combout ),
	.datab(\wdat[12]~39_combout ),
	.datac(plif_exmemporto_l_12),
	.datad(\FU|fwda~3_combout ),
	.cin(gnd),
	.combout(\porta~71_combout ),
	.cout());
// synopsys translate_off
defparam \porta~71 .lut_mask = 16'hE4A0;
defparam \porta~71 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y38_N18
cycloneive_lcell_comb \porta~72 (
// Equation(s):
// \porta~72_combout  = (always03 & (plif_exmemporto_l_11)) # (!always03 & (((\wdat[11]~41_combout  & fwda))))

	.dataa(plif_exmemporto_l_11),
	.datab(\wdat[11]~41_combout ),
	.datac(\FU|fwda~3_combout ),
	.datad(\FU|always0~8_combout ),
	.cin(gnd),
	.combout(\porta~72_combout ),
	.cout());
// synopsys translate_off
defparam \porta~72 .lut_mask = 16'hAAC0;
defparam \porta~72 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y34_N16
cycloneive_lcell_comb \porta~73 (
// Equation(s):
// \porta~73_combout  = (always03 & (plif_exmemporto_l_10)) # (!always03 & (((\wdat[10]~43_combout  & fwda))))

	.dataa(plif_exmemporto_l_10),
	.datab(\wdat[10]~43_combout ),
	.datac(\FU|always0~8_combout ),
	.datad(\FU|fwda~3_combout ),
	.cin(gnd),
	.combout(\porta~73_combout ),
	.cout());
// synopsys translate_off
defparam \porta~73 .lut_mask = 16'hACA0;
defparam \porta~73 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y41_N2
cycloneive_lcell_comb \porta~74 (
// Equation(s):
// \porta~74_combout  = (always03 & (plif_exmemporto_l_9)) # (!always03 & (((fwda & \wdat[9]~45_combout ))))

	.dataa(plif_exmemporto_l_9),
	.datab(\FU|fwda~3_combout ),
	.datac(\wdat[9]~45_combout ),
	.datad(\FU|always0~8_combout ),
	.cin(gnd),
	.combout(\porta~74_combout ),
	.cout());
// synopsys translate_off
defparam \porta~74 .lut_mask = 16'hAAC0;
defparam \porta~74 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y41_N2
cycloneive_lcell_comb \portb~65 (
// Equation(s):
// \portb~65_combout  = (\portb~2_combout  & ((plif_exmemporto_l_4) # ((!\portb~1_combout )))) # (!\portb~2_combout  & (((plif_idexextimm_l_4 & \portb~1_combout ))))

	.dataa(plif_exmemporto_l_4),
	.datab(\IDEX|plif_idex.extimm_l [4]),
	.datac(\portb~2_combout ),
	.datad(\portb~1_combout ),
	.cin(gnd),
	.combout(\portb~65_combout ),
	.cout());
// synopsys translate_off
defparam \portb~65 .lut_mask = 16'hACF0;
defparam \portb~65 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y41_N8
cycloneive_lcell_comb \portb~66 (
// Equation(s):
// \portb~66_combout  = (\portb~1_combout  & (((\portb~65_combout )))) # (!\portb~1_combout  & ((\portb~65_combout  & ((\wdat[4]~61_combout ))) # (!\portb~65_combout  & (plif_idexrdat2_l_4))))

	.dataa(\portb~1_combout ),
	.datab(\IDEX|plif_idex.rdat2_l [4]),
	.datac(\wdat[4]~61_combout ),
	.datad(\portb~65_combout ),
	.cin(gnd),
	.combout(\portb~66_combout ),
	.cout());
// synopsys translate_off
defparam \portb~66 .lut_mask = 16'hFA44;
defparam \portb~66 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y41_N28
cycloneive_lcell_comb \porta~75 (
// Equation(s):
// \porta~75_combout  = (always03 & (((plif_exmemporto_l_31)))) # (!always03 & (\wdat[31]~1_combout  & ((fwda))))

	.dataa(\wdat[31]~1_combout ),
	.datab(\FU|always0~8_combout ),
	.datac(plif_exmemporto_l_31),
	.datad(\FU|fwda~3_combout ),
	.cin(gnd),
	.combout(\porta~75_combout ),
	.cout());
// synopsys translate_off
defparam \porta~75 .lut_mask = 16'hE2C0;
defparam \porta~75 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y33_N18
cycloneive_lcell_comb \porta~76 (
// Equation(s):
// \porta~76_combout  = (always03 & (plif_exmemporto_l_29)) # (!always03 & (((fwda & \wdat[29]~5_combout ))))

	.dataa(plif_exmemporto_l_29),
	.datab(\FU|fwda~3_combout ),
	.datac(\wdat[29]~5_combout ),
	.datad(\FU|always0~8_combout ),
	.cin(gnd),
	.combout(\porta~76_combout ),
	.cout());
// synopsys translate_off
defparam \porta~76 .lut_mask = 16'hAAC0;
defparam \porta~76 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y42_N28
cycloneive_lcell_comb \porta~77 (
// Equation(s):
// \porta~77_combout  = (always03 & (((plif_exmemporto_l_30)))) # (!always03 & (\wdat[30]~3_combout  & ((fwda))))

	.dataa(\wdat[30]~3_combout ),
	.datab(plif_exmemporto_l_30),
	.datac(\FU|fwda~3_combout ),
	.datad(\FU|always0~8_combout ),
	.cin(gnd),
	.combout(\porta~77_combout ),
	.cout());
// synopsys translate_off
defparam \porta~77 .lut_mask = 16'hCCA0;
defparam \porta~77 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y35_N4
cycloneive_lcell_comb \porta~78 (
// Equation(s):
// \porta~78_combout  = (always03 & (((plif_exmemporto_l_28)))) # (!always03 & (fwda & ((\wdat[28]~7_combout ))))

	.dataa(\FU|always0~8_combout ),
	.datab(\FU|fwda~3_combout ),
	.datac(plif_exmemporto_l_28),
	.datad(\wdat[28]~7_combout ),
	.cin(gnd),
	.combout(\porta~78_combout ),
	.cout());
// synopsys translate_off
defparam \porta~78 .lut_mask = 16'hE4A0;
defparam \porta~78 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y36_N16
cycloneive_lcell_comb \porta~79 (
// Equation(s):
// \porta~79_combout  = (always03 & (plif_exmemporto_l_27)) # (!always03 & (((fwda & \wdat[27]~9_combout ))))

	.dataa(\FU|always0~8_combout ),
	.datab(plif_exmemporto_l_27),
	.datac(\FU|fwda~3_combout ),
	.datad(\wdat[27]~9_combout ),
	.cin(gnd),
	.combout(\porta~79_combout ),
	.cout());
// synopsys translate_off
defparam \porta~79 .lut_mask = 16'hD888;
defparam \porta~79 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y36_N24
cycloneive_lcell_comb \porta~80 (
// Equation(s):
// \porta~80_combout  = (always03 & (((plif_exmemporto_l_26)))) # (!always03 & (\wdat[26]~11_combout  & ((fwda))))

	.dataa(\wdat[26]~11_combout ),
	.datab(plif_exmemporto_l_26),
	.datac(\FU|fwda~3_combout ),
	.datad(\FU|always0~8_combout ),
	.cin(gnd),
	.combout(\porta~80_combout ),
	.cout());
// synopsys translate_off
defparam \porta~80 .lut_mask = 16'hCCA0;
defparam \porta~80 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y36_N18
cycloneive_lcell_comb \porta~81 (
// Equation(s):
// \porta~81_combout  = (always03 & (((plif_exmemporto_l_25)))) # (!always03 & (\wdat[25]~13_combout  & (fwda)))

	.dataa(\wdat[25]~13_combout ),
	.datab(\FU|fwda~3_combout ),
	.datac(\FU|always0~8_combout ),
	.datad(plif_exmemporto_l_25),
	.cin(gnd),
	.combout(\porta~81_combout ),
	.cout());
// synopsys translate_off
defparam \porta~81 .lut_mask = 16'hF808;
defparam \porta~81 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y35_N20
cycloneive_lcell_comb \porta~82 (
// Equation(s):
// \porta~82_combout  = (always03 & (plif_exmemporto_l_24)) # (!always03 & (((\wdat[24]~15_combout  & fwda))))

	.dataa(plif_exmemporto_l_24),
	.datab(\wdat[24]~15_combout ),
	.datac(\FU|fwda~3_combout ),
	.datad(\FU|always0~8_combout ),
	.cin(gnd),
	.combout(\porta~82_combout ),
	.cout());
// synopsys translate_off
defparam \porta~82 .lut_mask = 16'hAAC0;
defparam \porta~82 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X52_Y39_N0
cycloneive_lcell_comb \porta~83 (
// Equation(s):
// \porta~83_combout  = (always03 & (plif_exmemporto_l_23)) # (!always03 & (((\wdat[23]~17_combout  & fwda))))

	.dataa(plif_exmemporto_l_23),
	.datab(\wdat[23]~17_combout ),
	.datac(\FU|always0~8_combout ),
	.datad(\FU|fwda~3_combout ),
	.cin(gnd),
	.combout(\porta~83_combout ),
	.cout());
// synopsys translate_off
defparam \porta~83 .lut_mask = 16'hACA0;
defparam \porta~83 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y39_N20
cycloneive_lcell_comb \porta~84 (
// Equation(s):
// \porta~84_combout  = (always03 & (plif_exmemporto_l_22)) # (!always03 & (((\wdat[22]~19_combout  & fwda))))

	.dataa(plif_exmemporto_l_22),
	.datab(\wdat[22]~19_combout ),
	.datac(\FU|fwda~3_combout ),
	.datad(\FU|always0~8_combout ),
	.cin(gnd),
	.combout(\porta~84_combout ),
	.cout());
// synopsys translate_off
defparam \porta~84 .lut_mask = 16'hAAC0;
defparam \porta~84 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y38_N12
cycloneive_lcell_comb \porta~85 (
// Equation(s):
// \porta~85_combout  = (always03 & (((plif_exmemporto_l_21)))) # (!always03 & (\wdat[21]~21_combout  & (fwda)))

	.dataa(\FU|always0~8_combout ),
	.datab(\wdat[21]~21_combout ),
	.datac(\FU|fwda~3_combout ),
	.datad(plif_exmemporto_l_21),
	.cin(gnd),
	.combout(\porta~85_combout ),
	.cout());
// synopsys translate_off
defparam \porta~85 .lut_mask = 16'hEA40;
defparam \porta~85 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y39_N28
cycloneive_lcell_comb \porta~86 (
// Equation(s):
// \porta~86_combout  = (always03 & (plif_exmemporto_l_20)) # (!always03 & (((\wdat[20]~23_combout  & fwda))))

	.dataa(plif_exmemporto_l_20),
	.datab(\wdat[20]~23_combout ),
	.datac(\FU|always0~8_combout ),
	.datad(\FU|fwda~3_combout ),
	.cin(gnd),
	.combout(\porta~86_combout ),
	.cout());
// synopsys translate_off
defparam \porta~86 .lut_mask = 16'hACA0;
defparam \porta~86 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y36_N28
cycloneive_lcell_comb \porta~87 (
// Equation(s):
// \porta~87_combout  = (always03 & (((plif_exmemporto_l_19)))) # (!always03 & (\wdat[19]~25_combout  & ((fwda))))

	.dataa(\wdat[19]~25_combout ),
	.datab(plif_exmemporto_l_19),
	.datac(\FU|always0~8_combout ),
	.datad(\FU|fwda~3_combout ),
	.cin(gnd),
	.combout(\porta~87_combout ),
	.cout());
// synopsys translate_off
defparam \porta~87 .lut_mask = 16'hCAC0;
defparam \porta~87 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y37_N28
cycloneive_lcell_comb \porta~88 (
// Equation(s):
// \porta~88_combout  = (always03 & (plif_exmemporto_l_18)) # (!always03 & (((\wdat[18]~27_combout  & fwda))))

	.dataa(plif_exmemporto_l_18),
	.datab(\wdat[18]~27_combout ),
	.datac(\FU|always0~8_combout ),
	.datad(\FU|fwda~3_combout ),
	.cin(gnd),
	.combout(\porta~88_combout ),
	.cout());
// synopsys translate_off
defparam \porta~88 .lut_mask = 16'hACA0;
defparam \porta~88 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y40_N6
cycloneive_lcell_comb \porta~89 (
// Equation(s):
// \porta~89_combout  = (always03 & (((plif_exmemporto_l_17)))) # (!always03 & (\wdat[17]~29_combout  & ((fwda))))

	.dataa(\wdat[17]~29_combout ),
	.datab(plif_exmemporto_l_17),
	.datac(\FU|fwda~3_combout ),
	.datad(\FU|always0~8_combout ),
	.cin(gnd),
	.combout(\porta~89_combout ),
	.cout());
// synopsys translate_off
defparam \porta~89 .lut_mask = 16'hCCA0;
defparam \porta~89 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y40_N18
cycloneive_lcell_comb \porta~90 (
// Equation(s):
// \porta~90_combout  = (fwda & ((\wdat[0]~59_combout ))) # (!fwda & (plif_idexrdat1_l_0))

	.dataa(gnd),
	.datab(\IDEX|plif_idex.rdat1_l [0]),
	.datac(\wdat[0]~59_combout ),
	.datad(\FU|fwda~3_combout ),
	.cin(gnd),
	.combout(\porta~90_combout ),
	.cout());
// synopsys translate_off
defparam \porta~90 .lut_mask = 16'hF0CC;
defparam \porta~90 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y40_N20
cycloneive_lcell_comb \porta~91 (
// Equation(s):
// \porta~91_combout  = (always03 & (plif_exmemporto_l_0)) # (!always03 & ((\porta~90_combout )))

	.dataa(\FU|always0~8_combout ),
	.datab(plif_exmemporto_l_0),
	.datac(gnd),
	.datad(\porta~90_combout ),
	.cin(gnd),
	.combout(\porta~91_combout ),
	.cout());
// synopsys translate_off
defparam \porta~91 .lut_mask = 16'hDD88;
defparam \porta~91 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y32_N16
cycloneive_lcell_comb \pcsrc~0 (
// Equation(s):
// \pcsrc~0_combout  = (plif_memwbpcsrc_l_0 & ((plif_memwbpcsrc_l_1) # (plif_memwbbtype_l $ (plif_memwbzero_l))))

	.dataa(\MEMWB|plif_memwb.btype_l~q ),
	.datab(\MEMWB|plif_memwb.pcsrc_l [1]),
	.datac(\MEMWB|plif_memwb.zero_l~q ),
	.datad(\MEMWB|plif_memwb.pcsrc_l [0]),
	.cin(gnd),
	.combout(\pcsrc~0_combout ),
	.cout());
// synopsys translate_off
defparam \pcsrc~0 .lut_mask = 16'hDE00;
defparam \pcsrc~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y39_N4
cycloneive_lcell_comb \rdat2~64 (
// Equation(s):
// \rdat2~64_combout  = (always02 & (((plif_exmemporto_l_0)))) # (!always02 & (fwdc & ((\wdat[0]~59_combout ))))

	.dataa(\FU|fwdc~2_combout ),
	.datab(plif_exmemporto_l_0),
	.datac(\FU|always0~4_combout ),
	.datad(\wdat[0]~59_combout ),
	.cin(gnd),
	.combout(\rdat2~64_combout ),
	.cout());
// synopsys translate_off
defparam \rdat2~64 .lut_mask = 16'hCAC0;
defparam \rdat2~64 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y33_N2
cycloneive_lcell_comb \extimm[30]~0 (
// Equation(s):
// \extimm[30]~0_combout  = (!WideOr151 & (plif_ifidinstr_l_15 & WideOr142))

	.dataa(gnd),
	.datab(\CU|WideOr15~combout ),
	.datac(\IFID|plif_ifid.instr_l [15]),
	.datad(\CU|WideOr14~combout ),
	.cin(gnd),
	.combout(\extimm[30]~0_combout ),
	.cout());
// synopsys translate_off
defparam \extimm[30]~0 .lut_mask = 16'h3000;
defparam \extimm[30]~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y33_N24
cycloneive_lcell_comb \Equal0~0 (
// Equation(s):
// \Equal0~0_combout  = (Equal20 & (!Equal22 & (Selector22 & WideOr141)))

	.dataa(\CU|Equal20~0_combout ),
	.datab(\CU|Equal22~0_combout ),
	.datac(\CU|Selector22~6_combout ),
	.datad(\CU|WideOr14~0_combout ),
	.cin(gnd),
	.combout(\Equal0~0_combout ),
	.cout());
// synopsys translate_off
defparam \Equal0~0 .lut_mask = 16'h2000;
defparam \Equal0~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y34_N18
cycloneive_lcell_comb \rdat2~65 (
// Equation(s):
// \rdat2~65_combout  = (always02 & (((plif_exmemporto_l_1)))) # (!always02 & (fwdc & ((\wdat[1]~57_combout ))))

	.dataa(\FU|always0~4_combout ),
	.datab(\FU|fwdc~2_combout ),
	.datac(plif_exmemporto_l_1),
	.datad(\wdat[1]~57_combout ),
	.cin(gnd),
	.combout(\rdat2~65_combout ),
	.cout());
// synopsys translate_off
defparam \rdat2~65 .lut_mask = 16'hE4A0;
defparam \rdat2~65 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y35_N2
cycloneive_lcell_comb \rdat2~66 (
// Equation(s):
// \rdat2~66_combout  = (always02 & (plif_exmemporto_l_2)) # (!always02 & (((\wdat[2]~55_combout  & fwdc))))

	.dataa(plif_exmemporto_l_2),
	.datab(\wdat[2]~55_combout ),
	.datac(\FU|always0~4_combout ),
	.datad(\FU|fwdc~2_combout ),
	.cin(gnd),
	.combout(\rdat2~66_combout ),
	.cout());
// synopsys translate_off
defparam \rdat2~66 .lut_mask = 16'hACA0;
defparam \rdat2~66 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y34_N18
cycloneive_lcell_comb \rdat2~67 (
// Equation(s):
// \rdat2~67_combout  = (always02 & (((plif_exmemporto_l_3)))) # (!always02 & (fwdc & ((\wdat[3]~63_combout ))))

	.dataa(\FU|fwdc~2_combout ),
	.datab(\FU|always0~4_combout ),
	.datac(plif_exmemporto_l_3),
	.datad(\wdat[3]~63_combout ),
	.cin(gnd),
	.combout(\rdat2~67_combout ),
	.cout());
// synopsys translate_off
defparam \rdat2~67 .lut_mask = 16'hE2C0;
defparam \rdat2~67 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y41_N12
cycloneive_lcell_comb \rdat2~68 (
// Equation(s):
// \rdat2~68_combout  = (always02 & (((plif_exmemporto_l_4)))) # (!always02 & (\wdat[4]~61_combout  & (fwdc)))

	.dataa(\wdat[4]~61_combout ),
	.datab(\FU|fwdc~2_combout ),
	.datac(plif_exmemporto_l_4),
	.datad(\FU|always0~4_combout ),
	.cin(gnd),
	.combout(\rdat2~68_combout ),
	.cout());
// synopsys translate_off
defparam \rdat2~68 .lut_mask = 16'hF088;
defparam \rdat2~68 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y39_N22
cycloneive_lcell_comb \rdat2~69 (
// Equation(s):
// \rdat2~69_combout  = (always02 & (((plif_exmemporto_l_5)))) # (!always02 & (\wdat[5]~53_combout  & ((fwdc))))

	.dataa(\FU|always0~4_combout ),
	.datab(\wdat[5]~53_combout ),
	.datac(plif_exmemporto_l_5),
	.datad(\FU|fwdc~2_combout ),
	.cin(gnd),
	.combout(\rdat2~69_combout ),
	.cout());
// synopsys translate_off
defparam \rdat2~69 .lut_mask = 16'hE4A0;
defparam \rdat2~69 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y39_N12
cycloneive_lcell_comb \rdat2~70 (
// Equation(s):
// \rdat2~70_combout  = (always02 & (((plif_exmemporto_l_6)))) # (!always02 & (fwdc & ((\wdat[6]~51_combout ))))

	.dataa(\FU|fwdc~2_combout ),
	.datab(plif_exmemporto_l_6),
	.datac(\wdat[6]~51_combout ),
	.datad(\FU|always0~4_combout ),
	.cin(gnd),
	.combout(\rdat2~70_combout ),
	.cout());
// synopsys translate_off
defparam \rdat2~70 .lut_mask = 16'hCCA0;
defparam \rdat2~70 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y34_N26
cycloneive_lcell_comb \rdat2~71 (
// Equation(s):
// \rdat2~71_combout  = (always02 & (((plif_exmemporto_l_7)))) # (!always02 & (fwdc & (\wdat[7]~49_combout )))

	.dataa(\FU|always0~4_combout ),
	.datab(\FU|fwdc~2_combout ),
	.datac(\wdat[7]~49_combout ),
	.datad(plif_exmemporto_l_7),
	.cin(gnd),
	.combout(\rdat2~71_combout ),
	.cout());
// synopsys translate_off
defparam \rdat2~71 .lut_mask = 16'hEA40;
defparam \rdat2~71 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y34_N24
cycloneive_lcell_comb \rdat2~72 (
// Equation(s):
// \rdat2~72_combout  = (always02 & (plif_exmemporto_l_8)) # (!always02 & (((\wdat[8]~47_combout  & fwdc))))

	.dataa(plif_exmemporto_l_8),
	.datab(\FU|always0~4_combout ),
	.datac(\wdat[8]~47_combout ),
	.datad(\FU|fwdc~2_combout ),
	.cin(gnd),
	.combout(\rdat2~72_combout ),
	.cout());
// synopsys translate_off
defparam \rdat2~72 .lut_mask = 16'hB888;
defparam \rdat2~72 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y35_N0
cycloneive_lcell_comb \rdat2~73 (
// Equation(s):
// \rdat2~73_combout  = (always02 & (plif_exmemporto_l_9)) # (!always02 & (((\wdat[9]~45_combout  & fwdc))))

	.dataa(\FU|always0~4_combout ),
	.datab(plif_exmemporto_l_9),
	.datac(\wdat[9]~45_combout ),
	.datad(\FU|fwdc~2_combout ),
	.cin(gnd),
	.combout(\rdat2~73_combout ),
	.cout());
// synopsys translate_off
defparam \rdat2~73 .lut_mask = 16'hD888;
defparam \rdat2~73 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y34_N10
cycloneive_lcell_comb \rdat2~74 (
// Equation(s):
// \rdat2~74_combout  = (always02 & (plif_exmemporto_l_10)) # (!always02 & (((fwdc & \wdat[10]~43_combout ))))

	.dataa(plif_exmemporto_l_10),
	.datab(\FU|fwdc~2_combout ),
	.datac(\FU|always0~4_combout ),
	.datad(\wdat[10]~43_combout ),
	.cin(gnd),
	.combout(\rdat2~74_combout ),
	.cout());
// synopsys translate_off
defparam \rdat2~74 .lut_mask = 16'hACA0;
defparam \rdat2~74 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y39_N20
cycloneive_lcell_comb \rdat2~75 (
// Equation(s):
// \rdat2~75_combout  = (always02 & (plif_exmemporto_l_11)) # (!always02 & (((\wdat[11]~41_combout  & fwdc))))

	.dataa(\FU|always0~4_combout ),
	.datab(plif_exmemporto_l_11),
	.datac(\wdat[11]~41_combout ),
	.datad(\FU|fwdc~2_combout ),
	.cin(gnd),
	.combout(\rdat2~75_combout ),
	.cout());
// synopsys translate_off
defparam \rdat2~75 .lut_mask = 16'hD888;
defparam \rdat2~75 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y34_N12
cycloneive_lcell_comb \rdat2~76 (
// Equation(s):
// \rdat2~76_combout  = (always02 & (((plif_exmemporto_l_12)))) # (!always02 & (fwdc & ((\wdat[12]~39_combout ))))

	.dataa(\FU|always0~4_combout ),
	.datab(\FU|fwdc~2_combout ),
	.datac(plif_exmemporto_l_12),
	.datad(\wdat[12]~39_combout ),
	.cin(gnd),
	.combout(\rdat2~76_combout ),
	.cout());
// synopsys translate_off
defparam \rdat2~76 .lut_mask = 16'hE4A0;
defparam \rdat2~76 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y39_N14
cycloneive_lcell_comb \rdat2~77 (
// Equation(s):
// \rdat2~77_combout  = (always02 & (((plif_exmemporto_l_13)))) # (!always02 & (\wdat[13]~37_combout  & ((fwdc))))

	.dataa(\FU|always0~4_combout ),
	.datab(\wdat[13]~37_combout ),
	.datac(plif_exmemporto_l_13),
	.datad(\FU|fwdc~2_combout ),
	.cin(gnd),
	.combout(\rdat2~77_combout ),
	.cout());
// synopsys translate_off
defparam \rdat2~77 .lut_mask = 16'hE4A0;
defparam \rdat2~77 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y35_N22
cycloneive_lcell_comb \rdat2~78 (
// Equation(s):
// \rdat2~78_combout  = (always02 & (plif_exmemporto_l_14)) # (!always02 & (((fwdc & \wdat[14]~35_combout ))))

	.dataa(plif_exmemporto_l_14),
	.datab(\FU|fwdc~2_combout ),
	.datac(\wdat[14]~35_combout ),
	.datad(\FU|always0~4_combout ),
	.cin(gnd),
	.combout(\rdat2~78_combout ),
	.cout());
// synopsys translate_off
defparam \rdat2~78 .lut_mask = 16'hAAC0;
defparam \rdat2~78 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y40_N28
cycloneive_lcell_comb \rdat2~79 (
// Equation(s):
// \rdat2~79_combout  = (always02 & (((plif_exmemporto_l_15)))) # (!always02 & (\wdat[15]~33_combout  & ((fwdc))))

	.dataa(\wdat[15]~33_combout ),
	.datab(plif_exmemporto_l_15),
	.datac(\FU|always0~4_combout ),
	.datad(\FU|fwdc~2_combout ),
	.cin(gnd),
	.combout(\rdat2~79_combout ),
	.cout());
// synopsys translate_off
defparam \rdat2~79 .lut_mask = 16'hCAC0;
defparam \rdat2~79 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y35_N20
cycloneive_lcell_comb \rdat2~80 (
// Equation(s):
// \rdat2~80_combout  = (always02 & (((plif_exmemporto_l_16)))) # (!always02 & (\wdat[16]~31_combout  & ((fwdc))))

	.dataa(\wdat[16]~31_combout ),
	.datab(plif_exmemporto_l_16),
	.datac(\FU|always0~4_combout ),
	.datad(\FU|fwdc~2_combout ),
	.cin(gnd),
	.combout(\rdat2~80_combout ),
	.cout());
// synopsys translate_off
defparam \rdat2~80 .lut_mask = 16'hCAC0;
defparam \rdat2~80 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y39_N28
cycloneive_lcell_comb \rdat2~81 (
// Equation(s):
// \rdat2~81_combout  = (always02 & (((plif_exmemporto_l_17)))) # (!always02 & (fwdc & (\wdat[17]~29_combout )))

	.dataa(\FU|fwdc~2_combout ),
	.datab(\wdat[17]~29_combout ),
	.datac(\FU|always0~4_combout ),
	.datad(plif_exmemporto_l_17),
	.cin(gnd),
	.combout(\rdat2~81_combout ),
	.cout());
// synopsys translate_off
defparam \rdat2~81 .lut_mask = 16'hF808;
defparam \rdat2~81 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y37_N6
cycloneive_lcell_comb \rdat2~82 (
// Equation(s):
// \rdat2~82_combout  = (always02 & (((plif_exmemporto_l_18)))) # (!always02 & (fwdc & (\wdat[18]~27_combout )))

	.dataa(\FU|fwdc~2_combout ),
	.datab(\wdat[18]~27_combout ),
	.datac(plif_exmemporto_l_18),
	.datad(\FU|always0~4_combout ),
	.cin(gnd),
	.combout(\rdat2~82_combout ),
	.cout());
// synopsys translate_off
defparam \rdat2~82 .lut_mask = 16'hF088;
defparam \rdat2~82 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y34_N0
cycloneive_lcell_comb \rdat2~83 (
// Equation(s):
// \rdat2~83_combout  = (always02 & (((plif_exmemporto_l_19)))) # (!always02 & (\wdat[19]~25_combout  & (fwdc)))

	.dataa(\FU|always0~4_combout ),
	.datab(\wdat[19]~25_combout ),
	.datac(\FU|fwdc~2_combout ),
	.datad(plif_exmemporto_l_19),
	.cin(gnd),
	.combout(\rdat2~83_combout ),
	.cout());
// synopsys translate_off
defparam \rdat2~83 .lut_mask = 16'hEA40;
defparam \rdat2~83 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y39_N12
cycloneive_lcell_comb \rdat2~84 (
// Equation(s):
// \rdat2~84_combout  = (always02 & (((plif_exmemporto_l_20)))) # (!always02 & (fwdc & ((\wdat[20]~23_combout ))))

	.dataa(\FU|fwdc~2_combout ),
	.datab(\FU|always0~4_combout ),
	.datac(plif_exmemporto_l_20),
	.datad(\wdat[20]~23_combout ),
	.cin(gnd),
	.combout(\rdat2~84_combout ),
	.cout());
// synopsys translate_off
defparam \rdat2~84 .lut_mask = 16'hE2C0;
defparam \rdat2~84 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y38_N28
cycloneive_lcell_comb \rdat2~85 (
// Equation(s):
// \rdat2~85_combout  = (always02 & (((plif_exmemporto_l_21)))) # (!always02 & (fwdc & (\wdat[21]~21_combout )))

	.dataa(\FU|fwdc~2_combout ),
	.datab(\FU|always0~4_combout ),
	.datac(\wdat[21]~21_combout ),
	.datad(plif_exmemporto_l_21),
	.cin(gnd),
	.combout(\rdat2~85_combout ),
	.cout());
// synopsys translate_off
defparam \rdat2~85 .lut_mask = 16'hEC20;
defparam \rdat2~85 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y39_N2
cycloneive_lcell_comb \rdat2~86 (
// Equation(s):
// \rdat2~86_combout  = (always02 & (((plif_exmemporto_l_22)))) # (!always02 & (fwdc & (\wdat[22]~19_combout )))

	.dataa(\FU|fwdc~2_combout ),
	.datab(\wdat[22]~19_combout ),
	.datac(plif_exmemporto_l_22),
	.datad(\FU|always0~4_combout ),
	.cin(gnd),
	.combout(\rdat2~86_combout ),
	.cout());
// synopsys translate_off
defparam \rdat2~86 .lut_mask = 16'hF088;
defparam \rdat2~86 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X52_Y39_N4
cycloneive_lcell_comb \rdat2~87 (
// Equation(s):
// \rdat2~87_combout  = (always02 & (((plif_exmemporto_l_23)))) # (!always02 & (fwdc & ((\wdat[23]~17_combout ))))

	.dataa(\FU|always0~4_combout ),
	.datab(\FU|fwdc~2_combout ),
	.datac(plif_exmemporto_l_23),
	.datad(\wdat[23]~17_combout ),
	.cin(gnd),
	.combout(\rdat2~87_combout ),
	.cout());
// synopsys translate_off
defparam \rdat2~87 .lut_mask = 16'hE4A0;
defparam \rdat2~87 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y35_N4
cycloneive_lcell_comb \rdat2~88 (
// Equation(s):
// \rdat2~88_combout  = (always02 & (((plif_exmemporto_l_24)))) # (!always02 & (\wdat[24]~15_combout  & (fwdc)))

	.dataa(\FU|always0~4_combout ),
	.datab(\wdat[24]~15_combout ),
	.datac(\FU|fwdc~2_combout ),
	.datad(plif_exmemporto_l_24),
	.cin(gnd),
	.combout(\rdat2~88_combout ),
	.cout());
// synopsys translate_off
defparam \rdat2~88 .lut_mask = 16'hEA40;
defparam \rdat2~88 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y36_N28
cycloneive_lcell_comb \rdat2~89 (
// Equation(s):
// \rdat2~89_combout  = (always02 & (((plif_exmemporto_l_25)))) # (!always02 & (fwdc & ((\wdat[25]~13_combout ))))

	.dataa(\FU|always0~4_combout ),
	.datab(\FU|fwdc~2_combout ),
	.datac(plif_exmemporto_l_25),
	.datad(\wdat[25]~13_combout ),
	.cin(gnd),
	.combout(\rdat2~89_combout ),
	.cout());
// synopsys translate_off
defparam \rdat2~89 .lut_mask = 16'hE4A0;
defparam \rdat2~89 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y36_N8
cycloneive_lcell_comb \rdat2~90 (
// Equation(s):
// \rdat2~90_combout  = (always02 & (((plif_exmemporto_l_26)))) # (!always02 & (fwdc & ((\wdat[26]~11_combout ))))

	.dataa(\FU|always0~4_combout ),
	.datab(\FU|fwdc~2_combout ),
	.datac(plif_exmemporto_l_26),
	.datad(\wdat[26]~11_combout ),
	.cin(gnd),
	.combout(\rdat2~90_combout ),
	.cout());
// synopsys translate_off
defparam \rdat2~90 .lut_mask = 16'hE4A0;
defparam \rdat2~90 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y36_N22
cycloneive_lcell_comb \rdat2~91 (
// Equation(s):
// \rdat2~91_combout  = (always02 & (((plif_exmemporto_l_27)))) # (!always02 & (\wdat[27]~9_combout  & ((fwdc))))

	.dataa(\FU|always0~4_combout ),
	.datab(\wdat[27]~9_combout ),
	.datac(plif_exmemporto_l_27),
	.datad(\FU|fwdc~2_combout ),
	.cin(gnd),
	.combout(\rdat2~91_combout ),
	.cout());
// synopsys translate_off
defparam \rdat2~91 .lut_mask = 16'hE4A0;
defparam \rdat2~91 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y35_N8
cycloneive_lcell_comb \rdat2~92 (
// Equation(s):
// \rdat2~92_combout  = (always02 & (((plif_exmemporto_l_28)))) # (!always02 & (\wdat[28]~7_combout  & (fwdc)))

	.dataa(\wdat[28]~7_combout ),
	.datab(\FU|fwdc~2_combout ),
	.datac(plif_exmemporto_l_28),
	.datad(\FU|always0~4_combout ),
	.cin(gnd),
	.combout(\rdat2~92_combout ),
	.cout());
// synopsys translate_off
defparam \rdat2~92 .lut_mask = 16'hF088;
defparam \rdat2~92 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y34_N28
cycloneive_lcell_comb \rdat2~93 (
// Equation(s):
// \rdat2~93_combout  = (always02 & (((plif_exmemporto_l_29)))) # (!always02 & (\wdat[29]~5_combout  & (fwdc)))

	.dataa(\wdat[29]~5_combout ),
	.datab(\FU|fwdc~2_combout ),
	.datac(\FU|always0~4_combout ),
	.datad(plif_exmemporto_l_29),
	.cin(gnd),
	.combout(\rdat2~93_combout ),
	.cout());
// synopsys translate_off
defparam \rdat2~93 .lut_mask = 16'hF808;
defparam \rdat2~93 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y42_N6
cycloneive_lcell_comb \rdat2~94 (
// Equation(s):
// \rdat2~94_combout  = (always02 & (((plif_exmemporto_l_30)))) # (!always02 & (\wdat[30]~3_combout  & ((fwdc))))

	.dataa(\wdat[30]~3_combout ),
	.datab(plif_exmemporto_l_30),
	.datac(\FU|always0~4_combout ),
	.datad(\FU|fwdc~2_combout ),
	.cin(gnd),
	.combout(\rdat2~94_combout ),
	.cout());
// synopsys translate_off
defparam \rdat2~94 .lut_mask = 16'hCAC0;
defparam \rdat2~94 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y41_N2
cycloneive_lcell_comb \rdat2~95 (
// Equation(s):
// \rdat2~95_combout  = (always02 & (((plif_exmemporto_l_31)))) # (!always02 & (fwdc & ((\wdat[31]~1_combout ))))

	.dataa(\FU|always0~4_combout ),
	.datab(\FU|fwdc~2_combout ),
	.datac(plif_exmemporto_l_31),
	.datad(\wdat[31]~1_combout ),
	.cin(gnd),
	.combout(\rdat2~95_combout ),
	.cout());
// synopsys translate_off
defparam \rdat2~95 .lut_mask = 16'hE4A0;
defparam \rdat2~95 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y33_N16
cycloneive_lcell_comb \porta~92 (
// Equation(s):
// \porta~92_combout  = (\porta~62_combout ) # ((!always03 & (!fwda & plif_idexrdat1_l_8)))

	.dataa(\FU|always0~8_combout ),
	.datab(\FU|fwda~3_combout ),
	.datac(\IDEX|plif_idex.rdat1_l [8]),
	.datad(\porta~62_combout ),
	.cin(gnd),
	.combout(\porta~92_combout ),
	.cout());
// synopsys translate_off
defparam \porta~92 .lut_mask = 16'hFF10;
defparam \porta~92 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y38_N12
cycloneive_lcell_comb \porta~93 (
// Equation(s):
// \porta~93_combout  = (fwda & (((\porta~64_combout )))) # (!fwda & ((always03 & ((\porta~64_combout ))) # (!always03 & (plif_idexrdat1_l_7))))

	.dataa(\FU|fwda~3_combout ),
	.datab(\IDEX|plif_idex.rdat1_l [7]),
	.datac(\porta~64_combout ),
	.datad(\FU|always0~8_combout ),
	.cin(gnd),
	.combout(\porta~93_combout ),
	.cout());
// synopsys translate_off
defparam \porta~93 .lut_mask = 16'hF0E4;
defparam \porta~93 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y39_N24
cycloneive_lcell_comb \porta~94 (
// Equation(s):
// \porta~94_combout  = (\porta~65_combout ) # ((!fwda & (!always03 & plif_idexrdat1_l_6)))

	.dataa(\FU|fwda~3_combout ),
	.datab(\FU|always0~8_combout ),
	.datac(\IDEX|plif_idex.rdat1_l [6]),
	.datad(\porta~65_combout ),
	.cin(gnd),
	.combout(\porta~94_combout ),
	.cout());
// synopsys translate_off
defparam \porta~94 .lut_mask = 16'hFF10;
defparam \porta~94 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y38_N2
cycloneive_lcell_comb \porta~95 (
// Equation(s):
// \porta~95_combout  = (\porta~66_combout ) # ((!fwda & (plif_idexrdat1_l_5 & !always03)))

	.dataa(\FU|fwda~3_combout ),
	.datab(\IDEX|plif_idex.rdat1_l [5]),
	.datac(\porta~66_combout ),
	.datad(\FU|always0~8_combout ),
	.cin(gnd),
	.combout(\porta~95_combout ),
	.cout());
// synopsys translate_off
defparam \porta~95 .lut_mask = 16'hF0F4;
defparam \porta~95 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y35_N30
cycloneive_lcell_comb \porta~96 (
// Equation(s):
// \porta~96_combout  = (\porta~67_combout ) # ((plif_idexrdat1_l_16 & (!always03 & !fwda)))

	.dataa(\IDEX|plif_idex.rdat1_l [16]),
	.datab(\FU|always0~8_combout ),
	.datac(\FU|fwda~3_combout ),
	.datad(\porta~67_combout ),
	.cin(gnd),
	.combout(\porta~96_combout ),
	.cout());
// synopsys translate_off
defparam \porta~96 .lut_mask = 16'hFF02;
defparam \porta~96 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y40_N10
cycloneive_lcell_comb \porta~97 (
// Equation(s):
// \porta~97_combout  = (\porta~68_combout ) # ((!always03 & (plif_idexrdat1_l_15 & !fwda)))

	.dataa(\FU|always0~8_combout ),
	.datab(\IDEX|plif_idex.rdat1_l [15]),
	.datac(\FU|fwda~3_combout ),
	.datad(\porta~68_combout ),
	.cin(gnd),
	.combout(\porta~97_combout ),
	.cout());
// synopsys translate_off
defparam \porta~97 .lut_mask = 16'hFF04;
defparam \porta~97 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y41_N28
cycloneive_lcell_comb \porta~98 (
// Equation(s):
// \porta~98_combout  = (\porta~69_combout ) # ((!always03 & (!fwda & plif_idexrdat1_l_14)))

	.dataa(\FU|always0~8_combout ),
	.datab(\FU|fwda~3_combout ),
	.datac(\IDEX|plif_idex.rdat1_l [14]),
	.datad(\porta~69_combout ),
	.cin(gnd),
	.combout(\porta~98_combout ),
	.cout());
// synopsys translate_off
defparam \porta~98 .lut_mask = 16'hFF10;
defparam \porta~98 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y38_N22
cycloneive_lcell_comb \porta~99 (
// Equation(s):
// \porta~99_combout  = (\porta~70_combout ) # ((!always03 & (plif_idexrdat1_l_13 & !fwda)))

	.dataa(\FU|always0~8_combout ),
	.datab(\IDEX|plif_idex.rdat1_l [13]),
	.datac(\FU|fwda~3_combout ),
	.datad(\porta~70_combout ),
	.cin(gnd),
	.combout(\porta~99_combout ),
	.cout());
// synopsys translate_off
defparam \porta~99 .lut_mask = 16'hFF04;
defparam \porta~99 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y34_N30
cycloneive_lcell_comb \porta~100 (
// Equation(s):
// \porta~100_combout  = (\porta~71_combout ) # ((!always03 & (!fwda & plif_idexrdat1_l_12)))

	.dataa(\FU|always0~8_combout ),
	.datab(\FU|fwda~3_combout ),
	.datac(\IDEX|plif_idex.rdat1_l [12]),
	.datad(\porta~71_combout ),
	.cin(gnd),
	.combout(\porta~100_combout ),
	.cout());
// synopsys translate_off
defparam \porta~100 .lut_mask = 16'hFF10;
defparam \porta~100 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y38_N30
cycloneive_lcell_comb \porta~101 (
// Equation(s):
// \porta~101_combout  = (\porta~72_combout ) # ((plif_idexrdat1_l_11 & (!always03 & !fwda)))

	.dataa(\IDEX|plif_idex.rdat1_l [11]),
	.datab(\FU|always0~8_combout ),
	.datac(\FU|fwda~3_combout ),
	.datad(\porta~72_combout ),
	.cin(gnd),
	.combout(\porta~101_combout ),
	.cout());
// synopsys translate_off
defparam \porta~101 .lut_mask = 16'hFF02;
defparam \porta~101 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y34_N2
cycloneive_lcell_comb \porta~102 (
// Equation(s):
// \porta~102_combout  = (\porta~73_combout ) # ((plif_idexrdat1_l_10 & (!fwda & !always03)))

	.dataa(\IDEX|plif_idex.rdat1_l [10]),
	.datab(\FU|fwda~3_combout ),
	.datac(\FU|always0~8_combout ),
	.datad(\porta~73_combout ),
	.cin(gnd),
	.combout(\porta~102_combout ),
	.cout());
// synopsys translate_off
defparam \porta~102 .lut_mask = 16'hFF02;
defparam \porta~102 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y41_N22
cycloneive_lcell_comb \porta~103 (
// Equation(s):
// \porta~103_combout  = (\porta~74_combout ) # ((!always03 & (!fwda & plif_idexrdat1_l_9)))

	.dataa(\FU|always0~8_combout ),
	.datab(\FU|fwda~3_combout ),
	.datac(\IDEX|plif_idex.rdat1_l [9]),
	.datad(\porta~74_combout ),
	.cin(gnd),
	.combout(\porta~103_combout ),
	.cout());
// synopsys translate_off
defparam \porta~103 .lut_mask = 16'hFF10;
defparam \porta~103 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y41_N6
cycloneive_lcell_comb \porta~104 (
// Equation(s):
// \porta~104_combout  = (\porta~75_combout ) # ((plif_idexrdat1_l_31 & (!fwda & !always03)))

	.dataa(\IDEX|plif_idex.rdat1_l [31]),
	.datab(\FU|fwda~3_combout ),
	.datac(\FU|always0~8_combout ),
	.datad(\porta~75_combout ),
	.cin(gnd),
	.combout(\porta~104_combout ),
	.cout());
// synopsys translate_off
defparam \porta~104 .lut_mask = 16'hFF02;
defparam \porta~104 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y33_N10
cycloneive_lcell_comb \porta~105 (
// Equation(s):
// \porta~105_combout  = (\porta~76_combout ) # ((!always03 & (!fwda & plif_idexrdat1_l_29)))

	.dataa(\FU|always0~8_combout ),
	.datab(\FU|fwda~3_combout ),
	.datac(\IDEX|plif_idex.rdat1_l [29]),
	.datad(\porta~76_combout ),
	.cin(gnd),
	.combout(\porta~105_combout ),
	.cout());
// synopsys translate_off
defparam \porta~105 .lut_mask = 16'hFF10;
defparam \porta~105 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y42_N30
cycloneive_lcell_comb \porta~106 (
// Equation(s):
// \porta~106_combout  = (\porta~77_combout ) # ((plif_idexrdat1_l_30 & (!always03 & !fwda)))

	.dataa(\IDEX|plif_idex.rdat1_l [30]),
	.datab(\FU|always0~8_combout ),
	.datac(\FU|fwda~3_combout ),
	.datad(\porta~77_combout ),
	.cin(gnd),
	.combout(\porta~106_combout ),
	.cout());
// synopsys translate_off
defparam \porta~106 .lut_mask = 16'hFF02;
defparam \porta~106 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y35_N22
cycloneive_lcell_comb \porta~107 (
// Equation(s):
// \porta~107_combout  = (\porta~78_combout ) # ((!always03 & (plif_idexrdat1_l_28 & !fwda)))

	.dataa(\FU|always0~8_combout ),
	.datab(\IDEX|plif_idex.rdat1_l [28]),
	.datac(\porta~78_combout ),
	.datad(\FU|fwda~3_combout ),
	.cin(gnd),
	.combout(\porta~107_combout ),
	.cout());
// synopsys translate_off
defparam \porta~107 .lut_mask = 16'hF0F4;
defparam \porta~107 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y36_N4
cycloneive_lcell_comb \porta~108 (
// Equation(s):
// \porta~108_combout  = (\porta~79_combout ) # ((!always03 & (plif_idexrdat1_l_27 & !fwda)))

	.dataa(\FU|always0~8_combout ),
	.datab(\IDEX|plif_idex.rdat1_l [27]),
	.datac(\FU|fwda~3_combout ),
	.datad(\porta~79_combout ),
	.cin(gnd),
	.combout(\porta~108_combout ),
	.cout());
// synopsys translate_off
defparam \porta~108 .lut_mask = 16'hFF04;
defparam \porta~108 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y36_N2
cycloneive_lcell_comb \porta~109 (
// Equation(s):
// \porta~109_combout  = (\porta~80_combout ) # ((plif_idexrdat1_l_26 & (!always03 & !fwda)))

	.dataa(\IDEX|plif_idex.rdat1_l [26]),
	.datab(\FU|always0~8_combout ),
	.datac(\FU|fwda~3_combout ),
	.datad(\porta~80_combout ),
	.cin(gnd),
	.combout(\porta~109_combout ),
	.cout());
// synopsys translate_off
defparam \porta~109 .lut_mask = 16'hFF02;
defparam \porta~109 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y36_N10
cycloneive_lcell_comb \porta~110 (
// Equation(s):
// \porta~110_combout  = (\porta~81_combout ) # ((!always03 & (plif_idexrdat1_l_25 & !fwda)))

	.dataa(\FU|always0~8_combout ),
	.datab(\IDEX|plif_idex.rdat1_l [25]),
	.datac(\FU|fwda~3_combout ),
	.datad(\porta~81_combout ),
	.cin(gnd),
	.combout(\porta~110_combout ),
	.cout());
// synopsys translate_off
defparam \porta~110 .lut_mask = 16'hFF04;
defparam \porta~110 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y35_N6
cycloneive_lcell_comb \porta~111 (
// Equation(s):
// \porta~111_combout  = (\porta~82_combout ) # ((plif_idexrdat1_l_24 & (!always03 & !fwda)))

	.dataa(\IDEX|plif_idex.rdat1_l [24]),
	.datab(\FU|always0~8_combout ),
	.datac(\FU|fwda~3_combout ),
	.datad(\porta~82_combout ),
	.cin(gnd),
	.combout(\porta~111_combout ),
	.cout());
// synopsys translate_off
defparam \porta~111 .lut_mask = 16'hFF02;
defparam \porta~111 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X52_Y39_N18
cycloneive_lcell_comb \porta~112 (
// Equation(s):
// \porta~112_combout  = (\porta~83_combout ) # ((plif_idexrdat1_l_23 & (!fwda & !always03)))

	.dataa(\IDEX|plif_idex.rdat1_l [23]),
	.datab(\FU|fwda~3_combout ),
	.datac(\FU|always0~8_combout ),
	.datad(\porta~83_combout ),
	.cin(gnd),
	.combout(\porta~112_combout ),
	.cout());
// synopsys translate_off
defparam \porta~112 .lut_mask = 16'hFF02;
defparam \porta~112 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y39_N18
cycloneive_lcell_comb \porta~113 (
// Equation(s):
// \porta~113_combout  = (\porta~84_combout ) # ((plif_idexrdat1_l_22 & (!always03 & !fwda)))

	.dataa(\IDEX|plif_idex.rdat1_l [22]),
	.datab(\FU|always0~8_combout ),
	.datac(\FU|fwda~3_combout ),
	.datad(\porta~84_combout ),
	.cin(gnd),
	.combout(\porta~113_combout ),
	.cout());
// synopsys translate_off
defparam \porta~113 .lut_mask = 16'hFF02;
defparam \porta~113 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y38_N6
cycloneive_lcell_comb \porta~114 (
// Equation(s):
// \porta~114_combout  = (\porta~85_combout ) # ((!always03 & (plif_idexrdat1_l_21 & !fwda)))

	.dataa(\FU|always0~8_combout ),
	.datab(\IDEX|plif_idex.rdat1_l [21]),
	.datac(\FU|fwda~3_combout ),
	.datad(\porta~85_combout ),
	.cin(gnd),
	.combout(\porta~114_combout ),
	.cout());
// synopsys translate_off
defparam \porta~114 .lut_mask = 16'hFF04;
defparam \porta~114 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y39_N10
cycloneive_lcell_comb \porta~115 (
// Equation(s):
// \porta~115_combout  = (\porta~86_combout ) # ((!fwda & (plif_idexrdat1_l_20 & !always03)))

	.dataa(\FU|fwda~3_combout ),
	.datab(\IDEX|plif_idex.rdat1_l [20]),
	.datac(\FU|always0~8_combout ),
	.datad(\porta~86_combout ),
	.cin(gnd),
	.combout(\porta~115_combout ),
	.cout());
// synopsys translate_off
defparam \porta~115 .lut_mask = 16'hFF04;
defparam \porta~115 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y36_N22
cycloneive_lcell_comb \porta~116 (
// Equation(s):
// \porta~116_combout  = (\porta~87_combout ) # ((!fwda & (plif_idexrdat1_l_19 & !always03)))

	.dataa(\FU|fwda~3_combout ),
	.datab(\IDEX|plif_idex.rdat1_l [19]),
	.datac(\FU|always0~8_combout ),
	.datad(\porta~87_combout ),
	.cin(gnd),
	.combout(\porta~116_combout ),
	.cout());
// synopsys translate_off
defparam \porta~116 .lut_mask = 16'hFF04;
defparam \porta~116 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y37_N18
cycloneive_lcell_comb \porta~117 (
// Equation(s):
// \porta~117_combout  = (\porta~88_combout ) # ((!fwda & (plif_idexrdat1_l_18 & !always03)))

	.dataa(\FU|fwda~3_combout ),
	.datab(\IDEX|plif_idex.rdat1_l [18]),
	.datac(\FU|always0~8_combout ),
	.datad(\porta~88_combout ),
	.cin(gnd),
	.combout(\porta~117_combout ),
	.cout());
// synopsys translate_off
defparam \porta~117 .lut_mask = 16'hFF04;
defparam \porta~117 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y40_N26
cycloneive_lcell_comb \porta~118 (
// Equation(s):
// \porta~118_combout  = (\porta~89_combout ) # ((!always03 & (plif_idexrdat1_l_17 & !fwda)))

	.dataa(\FU|always0~8_combout ),
	.datab(\IDEX|plif_idex.rdat1_l [17]),
	.datac(\FU|fwda~3_combout ),
	.datad(\porta~89_combout ),
	.cin(gnd),
	.combout(\porta~118_combout ),
	.cout());
// synopsys translate_off
defparam \porta~118 .lut_mask = 16'hFF04;
defparam \porta~118 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y39_N0
cycloneive_lcell_comb \rdat2~96 (
// Equation(s):
// \rdat2~96_combout  = (\rdat2~64_combout ) # ((!fwdc & (!always02 & plif_idexrdat2_l_0)))

	.dataa(\FU|fwdc~2_combout ),
	.datab(\rdat2~64_combout ),
	.datac(\FU|always0~4_combout ),
	.datad(\IDEX|plif_idex.rdat2_l [0]),
	.cin(gnd),
	.combout(\rdat2~96_combout ),
	.cout());
// synopsys translate_off
defparam \rdat2~96 .lut_mask = 16'hCDCC;
defparam \rdat2~96 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y35_N2
cycloneive_lcell_comb \rdat2~97 (
// Equation(s):
// \rdat2~97_combout  = (\rdat2~65_combout ) # ((plif_idexrdat2_l_1 & (!fwdc & !always02)))

	.dataa(\IDEX|plif_idex.rdat2_l [1]),
	.datab(\FU|fwdc~2_combout ),
	.datac(\FU|always0~4_combout ),
	.datad(\rdat2~65_combout ),
	.cin(gnd),
	.combout(\rdat2~97_combout ),
	.cout());
// synopsys translate_off
defparam \rdat2~97 .lut_mask = 16'hFF02;
defparam \rdat2~97 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y39_N22
cycloneive_lcell_comb \rdat2~98 (
// Equation(s):
// \rdat2~98_combout  = (\rdat2~66_combout ) # ((!fwdc & (!always02 & plif_idexrdat2_l_2)))

	.dataa(\rdat2~66_combout ),
	.datab(\FU|fwdc~2_combout ),
	.datac(\FU|always0~4_combout ),
	.datad(\IDEX|plif_idex.rdat2_l [2]),
	.cin(gnd),
	.combout(\rdat2~98_combout ),
	.cout());
// synopsys translate_off
defparam \rdat2~98 .lut_mask = 16'hABAA;
defparam \rdat2~98 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y34_N28
cycloneive_lcell_comb \rdat2~99 (
// Equation(s):
// \rdat2~99_combout  = (\rdat2~67_combout ) # ((!fwdc & (!always02 & plif_idexrdat2_l_3)))

	.dataa(\FU|fwdc~2_combout ),
	.datab(\FU|always0~4_combout ),
	.datac(\IDEX|plif_idex.rdat2_l [3]),
	.datad(\rdat2~67_combout ),
	.cin(gnd),
	.combout(\rdat2~99_combout ),
	.cout());
// synopsys translate_off
defparam \rdat2~99 .lut_mask = 16'hFF10;
defparam \rdat2~99 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y41_N18
cycloneive_lcell_comb \rdat2~100 (
// Equation(s):
// \rdat2~100_combout  = (\rdat2~68_combout ) # ((!always02 & (plif_idexrdat2_l_4 & !fwdc)))

	.dataa(\FU|always0~4_combout ),
	.datab(\rdat2~68_combout ),
	.datac(\IDEX|plif_idex.rdat2_l [4]),
	.datad(\FU|fwdc~2_combout ),
	.cin(gnd),
	.combout(\rdat2~100_combout ),
	.cout());
// synopsys translate_off
defparam \rdat2~100 .lut_mask = 16'hCCDC;
defparam \rdat2~100 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y39_N2
cycloneive_lcell_comb \rdat2~101 (
// Equation(s):
// \rdat2~101_combout  = (\rdat2~69_combout ) # ((!always02 & (plif_idexrdat2_l_5 & !fwdc)))

	.dataa(\rdat2~69_combout ),
	.datab(\FU|always0~4_combout ),
	.datac(\IDEX|plif_idex.rdat2_l [5]),
	.datad(\FU|fwdc~2_combout ),
	.cin(gnd),
	.combout(\rdat2~101_combout ),
	.cout());
// synopsys translate_off
defparam \rdat2~101 .lut_mask = 16'hAABA;
defparam \rdat2~101 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y35_N6
cycloneive_lcell_comb \rdat2~102 (
// Equation(s):
// \rdat2~102_combout  = (\rdat2~70_combout ) # ((plif_idexrdat2_l_6 & (!always02 & !fwdc)))

	.dataa(\IDEX|plif_idex.rdat2_l [6]),
	.datab(\rdat2~70_combout ),
	.datac(\FU|always0~4_combout ),
	.datad(\FU|fwdc~2_combout ),
	.cin(gnd),
	.combout(\rdat2~102_combout ),
	.cout());
// synopsys translate_off
defparam \rdat2~102 .lut_mask = 16'hCCCE;
defparam \rdat2~102 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y34_N12
cycloneive_lcell_comb \rdat2~103 (
// Equation(s):
// \rdat2~103_combout  = (\rdat2~71_combout ) # ((!fwdc & (!always02 & plif_idexrdat2_l_7)))

	.dataa(\FU|fwdc~2_combout ),
	.datab(\FU|always0~4_combout ),
	.datac(\IDEX|plif_idex.rdat2_l [7]),
	.datad(\rdat2~71_combout ),
	.cin(gnd),
	.combout(\rdat2~103_combout ),
	.cout());
// synopsys translate_off
defparam \rdat2~103 .lut_mask = 16'hFF10;
defparam \rdat2~103 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y34_N20
cycloneive_lcell_comb \rdat2~104 (
// Equation(s):
// \rdat2~104_combout  = (\rdat2~72_combout ) # ((plif_idexrdat2_l_8 & (!fwdc & !always02)))

	.dataa(\IDEX|plif_idex.rdat2_l [8]),
	.datab(\rdat2~72_combout ),
	.datac(\FU|fwdc~2_combout ),
	.datad(\FU|always0~4_combout ),
	.cin(gnd),
	.combout(\rdat2~104_combout ),
	.cout());
// synopsys translate_off
defparam \rdat2~104 .lut_mask = 16'hCCCE;
defparam \rdat2~104 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y35_N18
cycloneive_lcell_comb \rdat2~105 (
// Equation(s):
// \rdat2~105_combout  = (\rdat2~73_combout ) # ((!always02 & (!fwdc & plif_idexrdat2_l_9)))

	.dataa(\FU|always0~4_combout ),
	.datab(\rdat2~73_combout ),
	.datac(\FU|fwdc~2_combout ),
	.datad(\IDEX|plif_idex.rdat2_l [9]),
	.cin(gnd),
	.combout(\rdat2~105_combout ),
	.cout());
// synopsys translate_off
defparam \rdat2~105 .lut_mask = 16'hCDCC;
defparam \rdat2~105 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y34_N14
cycloneive_lcell_comb \rdat2~106 (
// Equation(s):
// \rdat2~106_combout  = (\rdat2~74_combout ) # ((!always02 & (plif_idexrdat2_l_10 & !fwdc)))

	.dataa(\FU|always0~4_combout ),
	.datab(\IDEX|plif_idex.rdat2_l [10]),
	.datac(\FU|fwdc~2_combout ),
	.datad(\rdat2~74_combout ),
	.cin(gnd),
	.combout(\rdat2~106_combout ),
	.cout());
// synopsys translate_off
defparam \rdat2~106 .lut_mask = 16'hFF04;
defparam \rdat2~106 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y35_N24
cycloneive_lcell_comb \rdat2~107 (
// Equation(s):
// \rdat2~107_combout  = (\rdat2~75_combout ) # ((!fwdc & (plif_idexrdat2_l_11 & !always02)))

	.dataa(\rdat2~75_combout ),
	.datab(\FU|fwdc~2_combout ),
	.datac(\IDEX|plif_idex.rdat2_l [11]),
	.datad(\FU|always0~4_combout ),
	.cin(gnd),
	.combout(\rdat2~107_combout ),
	.cout());
// synopsys translate_off
defparam \rdat2~107 .lut_mask = 16'hAABA;
defparam \rdat2~107 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y34_N2
cycloneive_lcell_comb \rdat2~108 (
// Equation(s):
// \rdat2~108_combout  = (\rdat2~76_combout ) # ((!fwdc & (plif_idexrdat2_l_12 & !always02)))

	.dataa(\FU|fwdc~2_combout ),
	.datab(\rdat2~76_combout ),
	.datac(\IDEX|plif_idex.rdat2_l [12]),
	.datad(\FU|always0~4_combout ),
	.cin(gnd),
	.combout(\rdat2~108_combout ),
	.cout());
// synopsys translate_off
defparam \rdat2~108 .lut_mask = 16'hCCDC;
defparam \rdat2~108 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y39_N26
cycloneive_lcell_comb \rdat2~109 (
// Equation(s):
// \rdat2~109_combout  = (\rdat2~77_combout ) # ((!fwdc & (!always02 & plif_idexrdat2_l_13)))

	.dataa(\FU|fwdc~2_combout ),
	.datab(\rdat2~77_combout ),
	.datac(\FU|always0~4_combout ),
	.datad(\IDEX|plif_idex.rdat2_l [13]),
	.cin(gnd),
	.combout(\rdat2~109_combout ),
	.cout());
// synopsys translate_off
defparam \rdat2~109 .lut_mask = 16'hCDCC;
defparam \rdat2~109 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y35_N14
cycloneive_lcell_comb \rdat2~110 (
// Equation(s):
// \rdat2~110_combout  = (\rdat2~78_combout ) # ((!always02 & (plif_idexrdat2_l_14 & !fwdc)))

	.dataa(\FU|always0~4_combout ),
	.datab(\IDEX|plif_idex.rdat2_l [14]),
	.datac(\FU|fwdc~2_combout ),
	.datad(\rdat2~78_combout ),
	.cin(gnd),
	.combout(\rdat2~110_combout ),
	.cout());
// synopsys translate_off
defparam \rdat2~110 .lut_mask = 16'hFF04;
defparam \rdat2~110 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y35_N28
cycloneive_lcell_comb \rdat2~111 (
// Equation(s):
// \rdat2~111_combout  = (\rdat2~79_combout ) # ((!always02 & (!fwdc & plif_idexrdat2_l_15)))

	.dataa(\FU|always0~4_combout ),
	.datab(\FU|fwdc~2_combout ),
	.datac(\IDEX|plif_idex.rdat2_l [15]),
	.datad(\rdat2~79_combout ),
	.cin(gnd),
	.combout(\rdat2~111_combout ),
	.cout());
// synopsys translate_off
defparam \rdat2~111 .lut_mask = 16'hFF10;
defparam \rdat2~111 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y35_N12
cycloneive_lcell_comb \rdat2~112 (
// Equation(s):
// \rdat2~112_combout  = (\rdat2~80_combout ) # ((plif_idexrdat2_l_16 & (!always02 & !fwdc)))

	.dataa(\IDEX|plif_idex.rdat2_l [16]),
	.datab(\rdat2~80_combout ),
	.datac(\FU|always0~4_combout ),
	.datad(\FU|fwdc~2_combout ),
	.cin(gnd),
	.combout(\rdat2~112_combout ),
	.cout());
// synopsys translate_off
defparam \rdat2~112 .lut_mask = 16'hCCCE;
defparam \rdat2~112 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y39_N6
cycloneive_lcell_comb \rdat2~113 (
// Equation(s):
// \rdat2~113_combout  = (\rdat2~81_combout ) # ((!fwdc & (!always02 & plif_idexrdat2_l_17)))

	.dataa(\FU|fwdc~2_combout ),
	.datab(\FU|always0~4_combout ),
	.datac(\IDEX|plif_idex.rdat2_l [17]),
	.datad(\rdat2~81_combout ),
	.cin(gnd),
	.combout(\rdat2~113_combout ),
	.cout());
// synopsys translate_off
defparam \rdat2~113 .lut_mask = 16'hFF10;
defparam \rdat2~113 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y37_N22
cycloneive_lcell_comb \rdat2~114 (
// Equation(s):
// \rdat2~114_combout  = (\rdat2~82_combout ) # ((!fwdc & (plif_idexrdat2_l_18 & !always02)))

	.dataa(\FU|fwdc~2_combout ),
	.datab(\IDEX|plif_idex.rdat2_l [18]),
	.datac(\FU|always0~4_combout ),
	.datad(\rdat2~82_combout ),
	.cin(gnd),
	.combout(\rdat2~114_combout ),
	.cout());
// synopsys translate_off
defparam \rdat2~114 .lut_mask = 16'hFF04;
defparam \rdat2~114 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y34_N8
cycloneive_lcell_comb \rdat2~115 (
// Equation(s):
// \rdat2~115_combout  = (\rdat2~83_combout ) # ((!fwdc & (!always02 & plif_idexrdat2_l_19)))

	.dataa(\rdat2~83_combout ),
	.datab(\FU|fwdc~2_combout ),
	.datac(\FU|always0~4_combout ),
	.datad(\IDEX|plif_idex.rdat2_l [19]),
	.cin(gnd),
	.combout(\rdat2~115_combout ),
	.cout());
// synopsys translate_off
defparam \rdat2~115 .lut_mask = 16'hABAA;
defparam \rdat2~115 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y39_N14
cycloneive_lcell_comb \rdat2~116 (
// Equation(s):
// \rdat2~116_combout  = (\rdat2~84_combout ) # ((!always02 & (!fwdc & plif_idexrdat2_l_20)))

	.dataa(\rdat2~84_combout ),
	.datab(\FU|always0~4_combout ),
	.datac(\FU|fwdc~2_combout ),
	.datad(\IDEX|plif_idex.rdat2_l [20]),
	.cin(gnd),
	.combout(\rdat2~116_combout ),
	.cout());
// synopsys translate_off
defparam \rdat2~116 .lut_mask = 16'hABAA;
defparam \rdat2~116 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y34_N0
cycloneive_lcell_comb \rdat2~117 (
// Equation(s):
// \rdat2~117_combout  = (\rdat2~85_combout ) # ((!fwdc & (plif_idexrdat2_l_21 & !always02)))

	.dataa(\FU|fwdc~2_combout ),
	.datab(\rdat2~85_combout ),
	.datac(\IDEX|plif_idex.rdat2_l [21]),
	.datad(\FU|always0~4_combout ),
	.cin(gnd),
	.combout(\rdat2~117_combout ),
	.cout());
// synopsys translate_off
defparam \rdat2~117 .lut_mask = 16'hCCDC;
defparam \rdat2~117 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y39_N12
cycloneive_lcell_comb \rdat2~118 (
// Equation(s):
// \rdat2~118_combout  = (\rdat2~86_combout ) # ((!fwdc & (!always02 & plif_idexrdat2_l_22)))

	.dataa(\FU|fwdc~2_combout ),
	.datab(\rdat2~86_combout ),
	.datac(\FU|always0~4_combout ),
	.datad(\IDEX|plif_idex.rdat2_l [22]),
	.cin(gnd),
	.combout(\rdat2~118_combout ),
	.cout());
// synopsys translate_off
defparam \rdat2~118 .lut_mask = 16'hCDCC;
defparam \rdat2~118 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X52_Y39_N26
cycloneive_lcell_comb \rdat2~119 (
// Equation(s):
// \rdat2~119_combout  = (\rdat2~87_combout ) # ((plif_idexrdat2_l_23 & (!always02 & !fwdc)))

	.dataa(\IDEX|plif_idex.rdat2_l [23]),
	.datab(\rdat2~87_combout ),
	.datac(\FU|always0~4_combout ),
	.datad(\FU|fwdc~2_combout ),
	.cin(gnd),
	.combout(\rdat2~119_combout ),
	.cout());
// synopsys translate_off
defparam \rdat2~119 .lut_mask = 16'hCCCE;
defparam \rdat2~119 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y35_N18
cycloneive_lcell_comb \rdat2~120 (
// Equation(s):
// \rdat2~120_combout  = (\rdat2~88_combout ) # ((plif_idexrdat2_l_24 & (!fwdc & !always02)))

	.dataa(\IDEX|plif_idex.rdat2_l [24]),
	.datab(\FU|fwdc~2_combout ),
	.datac(\FU|always0~4_combout ),
	.datad(\rdat2~88_combout ),
	.cin(gnd),
	.combout(\rdat2~120_combout ),
	.cout());
// synopsys translate_off
defparam \rdat2~120 .lut_mask = 16'hFF02;
defparam \rdat2~120 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y36_N20
cycloneive_lcell_comb \rdat2~121 (
// Equation(s):
// \rdat2~121_combout  = (\rdat2~89_combout ) # ((!always02 & (!fwdc & plif_idexrdat2_l_25)))

	.dataa(\FU|always0~4_combout ),
	.datab(\FU|fwdc~2_combout ),
	.datac(\IDEX|plif_idex.rdat2_l [25]),
	.datad(\rdat2~89_combout ),
	.cin(gnd),
	.combout(\rdat2~121_combout ),
	.cout());
// synopsys translate_off
defparam \rdat2~121 .lut_mask = 16'hFF10;
defparam \rdat2~121 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y36_N2
cycloneive_lcell_comb \rdat2~122 (
// Equation(s):
// \rdat2~122_combout  = (\rdat2~90_combout ) # ((!always02 & (!fwdc & plif_idexrdat2_l_26)))

	.dataa(\FU|always0~4_combout ),
	.datab(\FU|fwdc~2_combout ),
	.datac(\IDEX|plif_idex.rdat2_l [26]),
	.datad(\rdat2~90_combout ),
	.cin(gnd),
	.combout(\rdat2~122_combout ),
	.cout());
// synopsys translate_off
defparam \rdat2~122 .lut_mask = 16'hFF10;
defparam \rdat2~122 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y36_N4
cycloneive_lcell_comb \rdat2~123 (
// Equation(s):
// \rdat2~123_combout  = (\rdat2~91_combout ) # ((!always02 & (plif_idexrdat2_l_27 & !fwdc)))

	.dataa(\FU|always0~4_combout ),
	.datab(\IDEX|plif_idex.rdat2_l [27]),
	.datac(\rdat2~91_combout ),
	.datad(\FU|fwdc~2_combout ),
	.cin(gnd),
	.combout(\rdat2~123_combout ),
	.cout());
// synopsys translate_off
defparam \rdat2~123 .lut_mask = 16'hF0F4;
defparam \rdat2~123 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y35_N30
cycloneive_lcell_comb \rdat2~124 (
// Equation(s):
// \rdat2~124_combout  = (\rdat2~92_combout ) # ((plif_idexrdat2_l_28 & (!fwdc & !always02)))

	.dataa(\IDEX|plif_idex.rdat2_l [28]),
	.datab(\FU|fwdc~2_combout ),
	.datac(\FU|always0~4_combout ),
	.datad(\rdat2~92_combout ),
	.cin(gnd),
	.combout(\rdat2~124_combout ),
	.cout());
// synopsys translate_off
defparam \rdat2~124 .lut_mask = 16'hFF02;
defparam \rdat2~124 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y34_N10
cycloneive_lcell_comb \rdat2~125 (
// Equation(s):
// \rdat2~125_combout  = (\rdat2~93_combout ) # ((!fwdc & (plif_idexrdat2_l_29 & !always02)))

	.dataa(\FU|fwdc~2_combout ),
	.datab(\rdat2~93_combout ),
	.datac(\IDEX|plif_idex.rdat2_l [29]),
	.datad(\FU|always0~4_combout ),
	.cin(gnd),
	.combout(\rdat2~125_combout ),
	.cout());
// synopsys translate_off
defparam \rdat2~125 .lut_mask = 16'hCCDC;
defparam \rdat2~125 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y42_N26
cycloneive_lcell_comb \rdat2~126 (
// Equation(s):
// \rdat2~126_combout  = (\rdat2~94_combout ) # ((!fwdc & (!always02 & plif_idexrdat2_l_30)))

	.dataa(\rdat2~94_combout ),
	.datab(\FU|fwdc~2_combout ),
	.datac(\FU|always0~4_combout ),
	.datad(\IDEX|plif_idex.rdat2_l [30]),
	.cin(gnd),
	.combout(\rdat2~126_combout ),
	.cout());
// synopsys translate_off
defparam \rdat2~126 .lut_mask = 16'hABAA;
defparam \rdat2~126 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y41_N24
cycloneive_lcell_comb \rdat2~127 (
// Equation(s):
// \rdat2~127_combout  = (\rdat2~95_combout ) # ((!always02 & (!fwdc & plif_idexrdat2_l_31)))

	.dataa(\FU|always0~4_combout ),
	.datab(\FU|fwdc~2_combout ),
	.datac(\rdat2~95_combout ),
	.datad(\IDEX|plif_idex.rdat2_l [31]),
	.cin(gnd),
	.combout(\rdat2~127_combout ),
	.cout());
// synopsys translate_off
defparam \rdat2~127 .lut_mask = 16'hF1F0;
defparam \rdat2~127 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X53_Y33_N25
dffeas \dpif.imemREN (
	.clk(CLK),
	.d(\dpif.imemREN~0_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(dpifimemREN),
	.prn(vcc));
// synopsys translate_off
defparam \dpif.imemREN .is_wysiwyg = "true";
defparam \dpif.imemREN .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X53_Y33_N24
cycloneive_lcell_comb \dpif.imemREN~0 (
// Equation(s):
// \dpif.imemREN~0_combout  = (dpifimemREN) # (plif_idexhlt_l)

	.dataa(gnd),
	.datab(gnd),
	.datac(dpifimemREN),
	.datad(\IDEX|plif_idex.hlt_l~q ),
	.cin(gnd),
	.combout(\dpif.imemREN~0_combout ),
	.cout());
// synopsys translate_off
defparam \dpif.imemREN~0 .lut_mask = 16'hFFF0;
defparam \dpif.imemREN~0 .sum_lutc_input = "datac";
// synopsys translate_on

endmodule

module alu (
	plif_idexaluop_l_3,
	plif_idexaluop_l_2,
	plif_idexaluop_l_1,
	plif_idexaluop_l_0,
	portb,
	portb1,
	portb2,
	portb3,
	portb4,
	portb5,
	portb6,
	portb7,
	portb8,
	portb9,
	portb10,
	portb11,
	portb12,
	portb13,
	portb14,
	portb15,
	portb16,
	portb17,
	portb18,
	portb19,
	portb20,
	portb21,
	portb22,
	portb23,
	portb24,
	portb25,
	portb26,
	porta,
	porta1,
	portb27,
	portb28,
	porta2,
	porta3,
	portb29,
	porta4,
	portb30,
	portb31,
	porta5,
	plif_idexrdat1_l_29,
	porta6,
	plif_idexrdat1_l_25,
	porta7,
	Selector30,
	Selector31,
	Selector28,
	Selector29,
	Selector26,
	Selector27,
	Selector24,
	Selector25,
	Selector22,
	Selector23,
	Selector20,
	Selector21,
	Selector18,
	Selector19,
	Selector16,
	Selector17,
	Selector14,
	Selector15,
	Selector12,
	Selector13,
	Selector10,
	Selector11,
	Selector8,
	Selector9,
	Selector6,
	Selector7,
	Selector4,
	Selector5,
	Selector2,
	Selector3,
	Selector0,
	Selector1,
	WideOr11,
	porta8,
	porta9,
	porta10,
	porta11,
	porta12,
	porta13,
	porta14,
	porta15,
	porta16,
	porta17,
	porta18,
	porta19,
	porta20,
	porta21,
	porta22,
	porta23,
	porta24,
	porta25,
	porta26,
	porta27,
	porta28,
	porta29,
	porta30,
	porta31,
	porta32,
	porta33,
	porta34,
	devpor,
	devclrn,
	devoe);
input 	plif_idexaluop_l_3;
input 	plif_idexaluop_l_2;
input 	plif_idexaluop_l_1;
input 	plif_idexaluop_l_0;
input 	portb;
input 	portb1;
input 	portb2;
input 	portb3;
input 	portb4;
input 	portb5;
input 	portb6;
input 	portb7;
input 	portb8;
input 	portb9;
input 	portb10;
input 	portb11;
input 	portb12;
input 	portb13;
input 	portb14;
input 	portb15;
input 	portb16;
input 	portb17;
input 	portb18;
input 	portb19;
input 	portb20;
input 	portb21;
input 	portb22;
input 	portb23;
input 	portb24;
input 	portb25;
input 	portb26;
input 	porta;
input 	porta1;
input 	portb27;
input 	portb28;
input 	porta2;
input 	porta3;
input 	portb29;
input 	porta4;
input 	portb30;
input 	portb31;
input 	porta5;
input 	plif_idexrdat1_l_29;
input 	porta6;
input 	plif_idexrdat1_l_25;
input 	porta7;
output 	Selector30;
output 	Selector31;
output 	Selector28;
output 	Selector29;
output 	Selector26;
output 	Selector27;
output 	Selector24;
output 	Selector25;
output 	Selector22;
output 	Selector23;
output 	Selector20;
output 	Selector21;
output 	Selector18;
output 	Selector19;
output 	Selector16;
output 	Selector17;
output 	Selector14;
output 	Selector15;
output 	Selector12;
output 	Selector13;
output 	Selector10;
output 	Selector11;
output 	Selector8;
output 	Selector9;
output 	Selector6;
output 	Selector7;
output 	Selector4;
output 	Selector5;
output 	Selector2;
output 	Selector3;
output 	Selector0;
output 	Selector1;
output 	WideOr11;
input 	porta8;
input 	porta9;
input 	porta10;
input 	porta11;
input 	porta12;
input 	porta13;
input 	porta14;
input 	porta15;
input 	porta16;
input 	porta17;
input 	porta18;
input 	porta19;
input 	porta20;
input 	porta21;
input 	porta22;
input 	porta23;
input 	porta24;
input 	porta25;
input 	porta26;
input 	porta27;
input 	porta28;
input 	porta29;
input 	porta30;
input 	porta31;
input 	porta32;
input 	porta33;
input 	porta34;

// Design Ports Information

input 	devpor;
input 	devclrn;
input 	devoe;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
assign unknown = 1'bx;

wire \Add1~0_combout ;
wire \Add1~2_combout ;
wire \Add0~14_combout ;
wire \ShiftRight0~7_combout ;
wire \ShiftRight0~12_combout ;
wire \ShiftRight0~14_combout ;
wire \ShiftRight0~16_combout ;
wire \ShiftRight0~18_combout ;
wire \ShiftRight0~37_combout ;
wire \ShiftRight0~42_combout ;
wire \ShiftRight0~43_combout ;
wire \ShiftRight0~44_combout ;
wire \ShiftRight0~48_combout ;
wire \Selector0~14_combout ;
wire \Selector29~5_combout ;
wire \ShiftRight0~100_combout ;
wire \Selector20~2_combout ;
wire \Selector21~3_combout ;
wire \Selector18~3_combout ;
wire \Selector19~2_combout ;
wire \Selector14~1_combout ;
wire \Selector13~4_combout ;
wire \Selector11~2_combout ;
wire \Selector8~6_combout ;
wire \Selector9~3_combout ;
wire \Selector9~4_combout ;
wire \ShiftLeft0~72_combout ;
wire \ShiftLeft0~79_combout ;
wire \WideOr1~5_combout ;
wire \ShiftRight0~22_combout ;
wire \ShiftRight0~24_combout ;
wire \ShiftRight0~25_combout ;
wire \ShiftRight0~26_combout ;
wire \ShiftRight0~10_combout ;
wire \ShiftRight0~11_combout ;
wire \ShiftRight0~9_combout ;
wire \Selector0~0_combout ;
wire \Selector24~0_combout ;
wire \ShiftRight0~27_combout ;
wire \ShiftRight0~28_combout ;
wire \ShiftRight0~30_combout ;
wire \ShiftRight0~29_combout ;
wire \ShiftRight0~31_combout ;
wire \ShiftRight0~32_combout ;
wire \ShiftRight0~36_combout ;
wire \ShiftRight0~38_combout ;
wire \ShiftRight0~34_combout ;
wire \ShiftRight0~33_combout ;
wire \ShiftRight0~35_combout ;
wire \Selector22~0_combout ;
wire \ShiftRight0~39_combout ;
wire \Selector30~0_combout ;
wire \Selector0~3_combout ;
wire \Selector0~7_combout ;
wire \Selector30~6_combout ;
wire \Selector0~4_combout ;
wire \Selector30~4_combout ;
wire \Selector0~2_combout ;
wire \ShiftLeft0~2_combout ;
wire \Selector1~0_combout ;
wire \Selector0~1_combout ;
wire \ShiftRight0~40_combout ;
wire \ShiftRight0~41_combout ;
wire \Selector30~1_combout ;
wire \Selector30~2_combout ;
wire \Selector30~3_combout ;
wire \Selector0~5_combout ;
wire \Selector0~6_combout ;
wire \Add0~1 ;
wire \Add0~2_combout ;
wire \Selector30~5_combout ;
wire \Selector30~7_combout ;
wire \Add0~0_combout ;
wire \Selector31~3_combout ;
wire \Selector31~4_combout ;
wire \ShiftRight0~71_combout ;
wire \Selector31~5_combout ;
wire \Selector31~6_combout ;
wire \Selector31~7_combout ;
wire \Selector31~1_combout ;
wire \LessThan0~1_cout ;
wire \LessThan0~3_cout ;
wire \LessThan0~5_cout ;
wire \LessThan0~7_cout ;
wire \LessThan0~9_cout ;
wire \LessThan0~11_cout ;
wire \LessThan0~13_cout ;
wire \LessThan0~15_cout ;
wire \LessThan0~17_cout ;
wire \LessThan0~19_cout ;
wire \LessThan0~21_cout ;
wire \LessThan0~23_cout ;
wire \LessThan0~25_cout ;
wire \LessThan0~27_cout ;
wire \LessThan0~29_cout ;
wire \LessThan0~31_cout ;
wire \LessThan0~33_cout ;
wire \LessThan0~35_cout ;
wire \LessThan0~37_cout ;
wire \LessThan0~39_cout ;
wire \LessThan0~41_cout ;
wire \LessThan0~43_cout ;
wire \LessThan0~45_cout ;
wire \LessThan0~47_cout ;
wire \LessThan0~49_cout ;
wire \LessThan0~51_cout ;
wire \LessThan0~53_cout ;
wire \LessThan0~55_cout ;
wire \LessThan0~57_cout ;
wire \LessThan0~59_cout ;
wire \LessThan0~61_cout ;
wire \LessThan0~62_combout ;
wire \LessThan1~1_cout ;
wire \LessThan1~3_cout ;
wire \LessThan1~5_cout ;
wire \LessThan1~7_cout ;
wire \LessThan1~9_cout ;
wire \LessThan1~11_cout ;
wire \LessThan1~13_cout ;
wire \LessThan1~15_cout ;
wire \LessThan1~17_cout ;
wire \LessThan1~19_cout ;
wire \LessThan1~21_cout ;
wire \LessThan1~23_cout ;
wire \LessThan1~25_cout ;
wire \LessThan1~27_cout ;
wire \LessThan1~29_cout ;
wire \LessThan1~31_cout ;
wire \LessThan1~33_cout ;
wire \LessThan1~35_cout ;
wire \LessThan1~37_cout ;
wire \LessThan1~39_cout ;
wire \LessThan1~41_cout ;
wire \LessThan1~43_cout ;
wire \LessThan1~45_cout ;
wire \LessThan1~47_cout ;
wire \LessThan1~49_cout ;
wire \LessThan1~51_cout ;
wire \LessThan1~53_cout ;
wire \LessThan1~55_cout ;
wire \LessThan1~57_cout ;
wire \LessThan1~59_cout ;
wire \LessThan1~61_cout ;
wire \LessThan1~62_combout ;
wire \Selector31~2_combout ;
wire \ShiftRight0~60_combout ;
wire \ShiftRight0~61_combout ;
wire \ShiftRight0~62_combout ;
wire \ShiftRight0~58_combout ;
wire \ShiftRight0~57_combout ;
wire \ShiftRight0~59_combout ;
wire \ShiftRight0~63_combout ;
wire \ShiftRight0~68_combout ;
wire \ShiftRight0~67_combout ;
wire \ShiftRight0~69_combout ;
wire \ShiftRight0~65_combout ;
wire \ShiftRight0~64_combout ;
wire \ShiftRight0~66_combout ;
wire \Selector23~0_combout ;
wire \ShiftRight0~70_combout ;
wire \ShiftRight0~50_combout ;
wire \ShiftRight0~49_combout ;
wire \ShiftRight0~51_combout ;
wire \ShiftRight0~52_combout ;
wire \ShiftRight0~53_combout ;
wire \ShiftRight0~54_combout ;
wire \ShiftRight0~55_combout ;
wire \ShiftRight0~56_combout ;
wire \Selector31~0_combout ;
wire \ShiftRight0~5_combout ;
wire \ShiftRight0~4_combout ;
wire \ShiftRight0~6_combout ;
wire \ShiftRight0~8_combout ;
wire \Selector0~15_combout ;
wire \Selector23~1_combout ;
wire \ShiftRight0~72_combout ;
wire \Selector3~0_combout ;
wire \Selector28~1_combout ;
wire \Selector3~1_combout ;
wire \ShiftRight0~13_combout ;
wire \ShiftRight0~15_combout ;
wire \ShiftRight0~23_combout ;
wire \ShiftRight0~73_combout ;
wire \Selector28~2_combout ;
wire \ShiftRight0~19_combout ;
wire \ShiftRight0~75_combout ;
wire \ShiftRight0~20_combout ;
wire \ShiftRight0~76_combout ;
wire \ShiftRight0~77_combout ;
wire \Selector28~3_combout ;
wire \Selector0~9_combout ;
wire \Add1~1 ;
wire \Add1~3 ;
wire \Add1~5 ;
wire \Add1~6_combout ;
wire \Add0~3 ;
wire \Add0~5 ;
wire \Add0~6_combout ;
wire \Selector28~0_combout ;
wire \Selector28~4_combout ;
wire \ShiftRight0~78_combout ;
wire \ShiftRight0~79_combout ;
wire \ShiftRight0~80_combout ;
wire \ShiftRight0~81_combout ;
wire \ShiftRight0~83_combout ;
wire \ShiftRight0~82_combout ;
wire \Selector20~0_combout ;
wire \ShiftRight0~84_combout ;
wire \ShiftLeft0~3_combout ;
wire \ShiftLeft0~4_combout ;
wire \Selector0~12_combout ;
wire \Selector28~6_combout ;
wire \Selector28~7_combout ;
wire \ShiftRight0~74_combout ;
wire \Selector28~8_combout ;
wire \Selector0~10_combout ;
wire \Selector0~11_combout ;
wire \Selector28~5_combout ;
wire \Selector28~9_combout ;
wire \Selector16~0_combout ;
wire \ShiftLeft0~5_combout ;
wire \ShiftLeft0~6_combout ;
wire \Selector29~0_combout ;
wire \ShiftRight0~92_combout ;
wire \ShiftRight0~91_combout ;
wire \Selector21~0_combout ;
wire \ShiftRight0~89_combout ;
wire \ShiftRight0~90_combout ;
wire \ShiftRight0~93_combout ;
wire \Selector0~13_combout ;
wire \Selector29~2_combout ;
wire \Selector29~3_combout ;
wire \Selector29~4_combout ;
wire \ShiftRight0~46_combout ;
wire \ShiftRight0~87_combout ;
wire \ShiftRight0~86_combout ;
wire \ShiftRight0~88_combout ;
wire \Selector29~6_combout ;
wire \Add1~4_combout ;
wire \Add0~4_combout ;
wire \Selector29~1_combout ;
wire \Selector29~7_combout ;
wire \Selector26~5_combout ;
wire \Selector26~6_combout ;
wire \Selector26~7_combout ;
wire \Selector1~1_combout ;
wire \ShiftLeft0~7_combout ;
wire \ShiftLeft0~8_combout ;
wire \ShiftLeft0~9_combout ;
wire \Selector26~0_combout ;
wire \Add1~7 ;
wire \Add1~9 ;
wire \Add1~10_combout ;
wire \Add0~7 ;
wire \Add0~9 ;
wire \Add0~10_combout ;
wire \Selector26~1_combout ;
wire \ShiftRight0~17_combout ;
wire \Selector7~0_combout ;
wire \Selector26~2_combout ;
wire \ShiftRight0~95_combout ;
wire \ShiftRight0~96_combout ;
wire \ShiftRight0~21_combout ;
wire \ShiftRight0~94_combout ;
wire \Selector26~3_combout ;
wire \Selector26~4_combout ;
wire \ShiftLeft0~10_combout ;
wire \ShiftLeft0~12_combout ;
wire \ShiftLeft0~11_combout ;
wire \ShiftLeft0~13_combout ;
wire \ShiftLeft0~14_combout ;
wire \Selector27~0_combout ;
wire \Selector27~5_combout ;
wire \Selector27~6_combout ;
wire \Selector27~7_combout ;
wire \Add0~8_combout ;
wire \Add1~8_combout ;
wire \Selector27~1_combout ;
wire \Selector7~1_combout ;
wire \ShiftRight0~98_combout ;
wire \ShiftRight0~99_combout ;
wire \ShiftRight0~45_combout ;
wire \ShiftRight0~47_combout ;
wire \ShiftRight0~97_combout ;
wire \Selector27~2_combout ;
wire \Selector27~3_combout ;
wire \Selector27~4_combout ;
wire \Selector24~6_combout ;
wire \Selector24~7_combout ;
wire \Selector24~8_combout ;
wire \Add1~11 ;
wire \Add1~13 ;
wire \Add1~14_combout ;
wire \Selector24~2_combout ;
wire \ShiftRight0~101_combout ;
wire \ShiftRight0~105_combout ;
wire \Selector24~3_combout ;
wire \Selector24~4_combout ;
wire \Selector24~5_combout ;
wire \ShiftLeft0~16_combout ;
wire \ShiftLeft0~17_combout ;
wire \Selector24~1_combout ;
wire \Selector24~10_combout ;
wire \ShiftLeft0~18_combout ;
wire \ShiftLeft0~19_combout ;
wire \ShiftLeft0~20_combout ;
wire \Selector25~5_combout ;
wire \Selector25~4_combout ;
wire \Selector25~6_combout ;
wire \Add0~11 ;
wire \Add0~12_combout ;
wire \Add1~12_combout ;
wire \Selector25~0_combout ;
wire \ShiftRight0~103_combout ;
wire \ShiftRight0~104_combout ;
wire \ShiftRight0~106_combout ;
wire \ShiftRight0~85_combout ;
wire \ShiftRight0~102_combout ;
wire \Selector25~1_combout ;
wire \Selector25~2_combout ;
wire \Selector25~3_combout ;
wire \Add0~13 ;
wire \Add0~15 ;
wire \Add0~17 ;
wire \Add0~18_combout ;
wire \Selector1~2_combout ;
wire \Selector16~1_combout ;
wire \Selector1~3_combout ;
wire \Selector20~1_combout ;
wire \Selector22~1_combout ;
wire \Add1~15 ;
wire \Add1~17 ;
wire \Add1~18_combout ;
wire \Selector0~8_combout ;
wire \ShiftLeft0~22_combout ;
wire \ShiftLeft0~21_combout ;
wire \ShiftLeft0~25_combout ;
wire \Selector22~2_combout ;
wire \Selector22~4_combout ;
wire \Selector22~5_combout ;
wire \Selector22~3_combout ;
wire \Selector22~6_combout ;
wire \Selector22~7_combout ;
wire \ShiftLeft0~27_combout ;
wire \ShiftLeft0~28_combout ;
wire \ShiftLeft0~26_combout ;
wire \ShiftLeft0~80_combout ;
wire \Add1~16_combout ;
wire \Selector23~6_combout ;
wire \Add0~16_combout ;
wire \Selector23~2_combout ;
wire \Selector23~3_combout ;
wire \Selector23~4_combout ;
wire \Selector23~5_combout ;
wire \Selector23~7_combout ;
wire \Selector0~16_combout ;
wire \Selector0~17_combout ;
wire \Selector23~8_combout ;
wire \ShiftLeft0~23_combout ;
wire \ShiftLeft0~29_combout ;
wire \ShiftLeft0~30_combout ;
wire \ShiftLeft0~31_combout ;
wire \ShiftLeft0~32_combout ;
wire \Selector20~8_combout ;
wire \Add1~19 ;
wire \Add1~21 ;
wire \Add1~22_combout ;
wire \Add0~19 ;
wire \Add0~21 ;
wire \Add0~22_combout ;
wire \Selector20~6_combout ;
wire \Selector20~3_combout ;
wire \Selector0~18_combout ;
wire \Selector20~4_combout ;
wire \Selector20~5_combout ;
wire \Selector20~7_combout ;
wire \ShiftLeft0~33_combout ;
wire \ShiftLeft0~34_combout ;
wire \ShiftLeft0~35_combout ;
wire \ShiftLeft0~36_combout ;
wire \Selector21~7_combout ;
wire \Selector21~4_combout ;
wire \Selector21~2_combout ;
wire \Add0~20_combout ;
wire \Add1~20_combout ;
wire \Selector21~1_combout ;
wire \Selector21~5_combout ;
wire \Selector21~6_combout ;
wire \Selector18~7_combout ;
wire \Selector18~6_combout ;
wire \Add1~23 ;
wire \Add1~25 ;
wire \Add1~26_combout ;
wire \Selector18~8_combout ;
wire \Add0~23 ;
wire \Add0~25 ;
wire \Add0~26_combout ;
wire \Selector18~0_combout ;
wire \Selector18~1_combout ;
wire \ShiftLeft0~37_combout ;
wire \ShiftLeft0~38_combout ;
wire \ShiftLeft0~15_combout ;
wire \ShiftLeft0~24_combout ;
wire \Selector10~0_combout ;
wire \ShiftLeft0~39_combout ;
wire \Selector18~4_combout ;
wire \Selector18~2_combout ;
wire \Selector18~5_combout ;
wire \Selector19~6_combout ;
wire \ShiftLeft0~40_combout ;
wire \ShiftLeft0~41_combout ;
wire \Selector11~0_combout ;
wire \Selector19~0_combout ;
wire \Selector19~3_combout ;
wire \Selector19~4_combout ;
wire \Selector19~1_combout ;
wire \Selector19~5_combout ;
wire \Add1~24_combout ;
wire \Add0~24_combout ;
wire \Selector19~7_combout ;
wire \Add1~27 ;
wire \Add1~29 ;
wire \Add1~30_combout ;
wire \Selector16~3_combout ;
wire \Selector16~2_combout ;
wire \Add0~27 ;
wire \Add0~29 ;
wire \Add0~30_combout ;
wire \Selector16~4_combout ;
wire \Selector16~5_combout ;
wire \Selector16~7_combout ;
wire \Selector16~8_combout ;
wire \ShiftLeft0~42_combout ;
wire \ShiftLeft0~43_combout ;
wire \Selector8~0_combout ;
wire \ShiftLeft0~44_combout ;
wire \Selector16~6_combout ;
wire \Selector16~9_combout ;
wire \Add0~28_combout ;
wire \Selector17~4_combout ;
wire \Selector17~5_combout ;
wire \Add1~28_combout ;
wire \Selector17~6_combout ;
wire \Selector17~2_combout ;
wire \ShiftLeft0~46_combout ;
wire \Selector9~0_combout ;
wire \ShiftLeft0~47_combout ;
wire \Selector17~0_combout ;
wire \Selector17~1_combout ;
wire \Selector17~3_combout ;
wire \Add1~31 ;
wire \Add1~33 ;
wire \Add1~34_combout ;
wire \Selector1~4_combout ;
wire \Selector14~6_combout ;
wire \Selector14~7_combout ;
wire \Add0~31 ;
wire \Add0~33 ;
wire \Add0~34_combout ;
wire \Selector14~2_combout ;
wire \Selector14~0_combout ;
wire \Selector0~19_combout ;
wire \Selector14~3_combout ;
wire \Selector0~21_combout ;
wire \ShiftLeft0~48_combout ;
wire \ShiftLeft0~49_combout ;
wire \ShiftLeft0~50_combout ;
wire \Selector14~4_combout ;
wire \Selector14~5_combout ;
wire \Selector0~20_combout ;
wire \Selector8~1_combout ;
wire \Selector15~0_combout ;
wire \Add1~32_combout ;
wire \Selector15~3_combout ;
wire \ShiftLeft0~45_combout ;
wire \ShiftLeft0~51_combout ;
wire \ShiftLeft0~52_combout ;
wire \ShiftLeft0~53_combout ;
wire \Selector15~1_combout ;
wire \Selector15~2_combout ;
wire \Selector15~4_combout ;
wire \Add0~32_combout ;
wire \Selector15~5_combout ;
wire \Selector15~6_combout ;
wire \Selector15~7_combout ;
wire \Add0~35 ;
wire \Add0~37 ;
wire \Add0~38_combout ;
wire \Add1~35 ;
wire \Add1~37 ;
wire \Add1~38_combout ;
wire \Selector12~9_combout ;
wire \Selector12~2_combout ;
wire \Selector12~5_combout ;
wire \Selector12~6_combout ;
wire \Selector12~4_combout ;
wire \Selector12~12_combout ;
wire \ShiftLeft0~54_combout ;
wire \ShiftLeft0~55_combout ;
wire \ShiftLeft0~56_combout ;
wire \Selector12~3_combout ;
wire \Selector12~7_combout ;
wire \Selector12~8_combout ;
wire \Add1~36_combout ;
wire \Add0~36_combout ;
wire \Selector13~1_combout ;
wire \Selector13~2_combout ;
wire \Selector13~3_combout ;
wire \Selector12~11_combout ;
wire \Selector13~5_combout ;
wire \Selector13~6_combout ;
wire \Selector13~7_combout ;
wire \Selector13~0_combout ;
wire \Selector10~1_combout ;
wire \Add0~39 ;
wire \Add0~41 ;
wire \Add0~42_combout ;
wire \Selector10~5_combout ;
wire \Selector10~6_combout ;
wire \Add1~39 ;
wire \Add1~41 ;
wire \Add1~42_combout ;
wire \Selector8~2_combout ;
wire \Selector10~3_combout ;
wire \ShiftLeft0~62_combout ;
wire \Selector10~2_combout ;
wire \Selector10~4_combout ;
wire \Selector10~7_combout ;
wire \Add0~40_combout ;
wire \Add1~40_combout ;
wire \Selector11~4_combout ;
wire \Selector11~1_combout ;
wire \Selector11~3_combout ;
wire \Selector11~5_combout ;
wire \Selector11~7_combout ;
wire \Selector11~6_combout ;
wire \Selector11~8_combout ;
wire \Selector8~7_combout ;
wire \Selector8~8_combout ;
wire \Add0~43 ;
wire \Add0~45 ;
wire \Add0~46_combout ;
wire \Selector8~9_combout ;
wire \Add1~43 ;
wire \Add1~45 ;
wire \Add1~46_combout ;
wire \ShiftLeft0~60_combout ;
wire \ShiftLeft0~66_combout ;
wire \ShiftLeft0~67_combout ;
wire \Selector8~3_combout ;
wire \Selector8~4_combout ;
wire \Selector8~5_combout ;
wire \Selector9~1_combout ;
wire \Add1~44_combout ;
wire \Selector9~2_combout ;
wire \Add0~44_combout ;
wire \ShiftLeft0~57_combout ;
wire \ShiftLeft0~58_combout ;
wire \ShiftLeft0~68_combout ;
wire \ShiftLeft0~69_combout ;
wire \Selector1~5_combout ;
wire \Selector9~5_combout ;
wire \Selector9~6_combout ;
wire \Selector9~7_combout ;
wire \Add1~47 ;
wire \Add1~49 ;
wire \Add1~50_combout ;
wire \Add0~47 ;
wire \Add0~49 ;
wire \Add0~50_combout ;
wire \Selector6~7_combout ;
wire \Selector4~0_combout ;
wire \Selector6~0_combout ;
wire \porto~0_combout ;
wire \Selector6~1_combout ;
wire \Selector6~2_combout ;
wire \ShiftLeft0~70_combout ;
wire \ShiftLeft0~71_combout ;
wire \ShiftLeft0~61_combout ;
wire \Selector6~3_combout ;
wire \Selector6~4_combout ;
wire \Selector6~5_combout ;
wire \Selector6~6_combout ;
wire \Selector7~9_combout ;
wire \Selector7~8_combout ;
wire \Selector7~10_combout ;
wire \Add0~48_combout ;
wire \Add1~48_combout ;
wire \Selector7~2_combout ;
wire \Selector7~3_combout ;
wire \ShiftLeft0~73_combout ;
wire \Selector7~4_combout ;
wire \ShiftLeft0~63_combout ;
wire \ShiftLeft0~64_combout ;
wire \Selector7~5_combout ;
wire \Selector7~6_combout ;
wire \Selector7~7_combout ;
wire \Selector4~8_combout ;
wire \Selector4~7_combout ;
wire \Selector4~9_combout ;
wire \Add1~51 ;
wire \Add1~53 ;
wire \Add1~54_combout ;
wire \Selector4~4_combout ;
wire \Selector4~5_combout ;
wire \Add0~51 ;
wire \Add0~53 ;
wire \Add0~54_combout ;
wire \ShiftLeft0~74_combout ;
wire \ShiftLeft0~75_combout ;
wire \Selector4~1_combout ;
wire \Selector4~2_combout ;
wire \Selector4~3_combout ;
wire \Selector4~6_combout ;
wire \Add0~52_combout ;
wire \Selector5~0_combout ;
wire \Selector5~1_combout ;
wire \Selector5~2_combout ;
wire \ShiftLeft0~76_combout ;
wire \ShiftLeft0~77_combout ;
wire \ShiftLeft0~59_combout ;
wire \Selector5~3_combout ;
wire \Selector5~4_combout ;
wire \Selector5~5_combout ;
wire \Selector5~6_combout ;
wire \Add1~52_combout ;
wire \Selector5~7_combout ;
wire \Add1~55 ;
wire \Add1~57 ;
wire \Add1~58_combout ;
wire \Add0~55 ;
wire \Add0~57 ;
wire \Add0~58_combout ;
wire \Selector2~10_combout ;
wire \Selector2~0_combout ;
wire \Selector2~1_combout ;
wire \porto~1_combout ;
wire \Selector2~2_combout ;
wire \Selector2~3_combout ;
wire \Selector2~4_combout ;
wire \ShiftLeft0~78_combout ;
wire \Selector2~6_combout ;
wire \Selector2~7_combout ;
wire \Selector2~5_combout ;
wire \Selector2~8_combout ;
wire \Selector2~9_combout ;
wire \Add0~56_combout ;
wire \Selector3~10_combout ;
wire \Add1~56_combout ;
wire \Selector3~3_combout ;
wire \Selector3~4_combout ;
wire \Selector3~2_combout ;
wire \Selector3~5_combout ;
wire \Selector3~6_combout ;
wire \ShiftLeft0~65_combout ;
wire \Selector3~7_combout ;
wire \Selector3~8_combout ;
wire \Selector3~9_combout ;
wire \Selector0~23_combout ;
wire \Selector0~24_combout ;
wire \Add0~59 ;
wire \Add0~61 ;
wire \Add0~62_combout ;
wire \Selector0~25_combout ;
wire \Selector0~26_combout ;
wire \Selector0~27_combout ;
wire \Selector0~28_combout ;
wire \Selector0~29_combout ;
wire \Add1~59 ;
wire \Add1~61 ;
wire \Add1~62_combout ;
wire \Selector1~6_combout ;
wire \Selector0~30_combout ;
wire \Selector0~31_combout ;
wire \Selector0~32_combout ;
wire \Selector0~33_combout ;
wire \Selector0~22_combout ;
wire \Selector1~7_combout ;
wire \Selector1~8_combout ;
wire \Add0~60_combout ;
wire \Selector1~18_combout ;
wire \Add1~60_combout ;
wire \Selector1~9_combout ;
wire \Selector1~10_combout ;
wire \Selector1~14_combout ;
wire \Selector1~15_combout ;
wire \Selector1~16_combout ;
wire \Selector1~11_combout ;
wire \Selector1~12_combout ;
wire \Selector1~13_combout ;
wire \Selector1~17_combout ;
wire \Selector1~19_combout ;
wire \WideOr1~0_combout ;
wire \WideOr1~6_combout ;
wire \WideOr1~7_combout ;
wire \WideOr1~8_combout ;
wire \WideOr1~9_combout ;
wire \WideOr1~10_combout ;
wire \WideOr1~1_combout ;
wire \WideOr1~2_combout ;
wire \WideOr1~3_combout ;
wire \WideOr1~4_combout ;
wire \WideOr1~11_combout ;


// Location: LCCOMB_X57_Y40_N0
cycloneive_lcell_comb \Add1~0 (
// Equation(s):
// \Add1~0_combout  = (\portb~58_combout  & (\porta~91_combout  $ (VCC))) # (!\portb~58_combout  & ((\porta~91_combout ) # (GND)))
// \Add1~1  = CARRY((\porta~91_combout ) # (!\portb~58_combout ))

	.dataa(portb27),
	.datab(porta7),
	.datac(gnd),
	.datad(vcc),
	.cin(gnd),
	.combout(\Add1~0_combout ),
	.cout(\Add1~1 ));
// synopsys translate_off
defparam \Add1~0 .lut_mask = 16'h66DD;
defparam \Add1~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y40_N2
cycloneive_lcell_comb \Add1~2 (
// Equation(s):
// \Add1~2_combout  = (\portb~60_combout  & ((\porta~57_combout  & (!\Add1~1 )) # (!\porta~57_combout  & ((\Add1~1 ) # (GND))))) # (!\portb~60_combout  & ((\porta~57_combout  & (\Add1~1  & VCC)) # (!\porta~57_combout  & (!\Add1~1 ))))
// \Add1~3  = CARRY((\portb~60_combout  & ((!\Add1~1 ) # (!\porta~57_combout ))) # (!\portb~60_combout  & (!\porta~57_combout  & !\Add1~1 )))

	.dataa(portb28),
	.datab(porta1),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add1~1 ),
	.combout(\Add1~2_combout ),
	.cout(\Add1~3 ));
// synopsys translate_off
defparam \Add1~2 .lut_mask = 16'h692B;
defparam \Add1~2 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X52_Y38_N14
cycloneive_lcell_comb \Add0~14 (
// Equation(s):
// \Add0~14_combout  = (\portb~52_combout  & ((\porta~93_combout  & (\Add0~13  & VCC)) # (!\porta~93_combout  & (!\Add0~13 )))) # (!\portb~52_combout  & ((\porta~93_combout  & (!\Add0~13 )) # (!\porta~93_combout  & ((\Add0~13 ) # (GND)))))
// \Add0~15  = CARRY((\portb~52_combout  & (!\porta~93_combout  & !\Add0~13 )) # (!\portb~52_combout  & ((!\Add0~13 ) # (!\porta~93_combout ))))

	.dataa(portb24),
	.datab(porta9),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add0~13 ),
	.combout(\Add0~14_combout ),
	.cout(\Add0~15 ));
// synopsys translate_off
defparam \Add0~14 .lut_mask = 16'h9617;
defparam \Add0~14 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X54_Y38_N6
cycloneive_lcell_comb \ShiftRight0~7 (
// Equation(s):
// \ShiftRight0~7_combout  = (\portb~30_combout ) # ((\portb~32_combout ) # ((\portb~34_combout ) # (\portb~28_combout )))

	.dataa(portb13),
	.datab(portb14),
	.datac(portb15),
	.datad(portb12),
	.cin(gnd),
	.combout(\ShiftRight0~7_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftRight0~7 .lut_mask = 16'hFFFE;
defparam \ShiftRight0~7 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y41_N16
cycloneive_lcell_comb \ShiftRight0~12 (
// Equation(s):
// \ShiftRight0~12_combout  = (!\portb~60_combout  & ((\portb~58_combout  & (\porta~55_combout )) # (!\portb~58_combout  & ((\porta~57_combout )))))

	.dataa(porta),
	.datab(portb27),
	.datac(porta1),
	.datad(portb28),
	.cin(gnd),
	.combout(\ShiftRight0~12_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftRight0~12 .lut_mask = 16'h00B8;
defparam \ShiftRight0~12 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y41_N18
cycloneive_lcell_comb \ShiftRight0~14 (
// Equation(s):
// \ShiftRight0~14_combout  = (!\portb~62_combout  & ((\ShiftRight0~12_combout ) # ((\portb~60_combout  & \ShiftRight0~13_combout ))))

	.dataa(portb29),
	.datab(\ShiftRight0~12_combout ),
	.datac(portb28),
	.datad(\ShiftRight0~13_combout ),
	.cin(gnd),
	.combout(\ShiftRight0~14_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftRight0~14 .lut_mask = 16'h5444;
defparam \ShiftRight0~14 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X52_Y41_N30
cycloneive_lcell_comb \ShiftRight0~16 (
// Equation(s):
// \ShiftRight0~16_combout  = (\portb~58_combout  & ((\porta~94_combout ))) # (!\portb~58_combout  & (\porta~95_combout ))

	.dataa(gnd),
	.datab(porta11),
	.datac(porta10),
	.datad(portb27),
	.cin(gnd),
	.combout(\ShiftRight0~16_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftRight0~16 .lut_mask = 16'hF0CC;
defparam \ShiftRight0~16 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y41_N22
cycloneive_lcell_comb \ShiftRight0~18 (
// Equation(s):
// \ShiftRight0~18_combout  = (!\portb~64_combout  & ((\ShiftRight0~14_combout ) # ((\portb~62_combout  & \ShiftRight0~17_combout ))))

	.dataa(\ShiftRight0~14_combout ),
	.datab(portb29),
	.datac(portb30),
	.datad(\ShiftRight0~17_combout ),
	.cin(gnd),
	.combout(\ShiftRight0~18_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftRight0~18 .lut_mask = 16'h0E0A;
defparam \ShiftRight0~18 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y40_N30
cycloneive_lcell_comb \ShiftRight0~37 (
// Equation(s):
// \ShiftRight0~37_combout  = (\portb~58_combout  & ((\porta~117_combout ))) # (!\portb~58_combout  & (\porta~118_combout ))

	.dataa(gnd),
	.datab(portb27),
	.datac(porta34),
	.datad(porta33),
	.cin(gnd),
	.combout(\ShiftRight0~37_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftRight0~37 .lut_mask = 16'hFC30;
defparam \ShiftRight0~37 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X52_Y35_N10
cycloneive_lcell_comb \ShiftRight0~42 (
// Equation(s):
// \ShiftRight0~42_combout  = (!\portb~60_combout  & ((\portb~58_combout  & (\porta~57_combout )) # (!\portb~58_combout  & ((\porta~91_combout )))))

	.dataa(portb28),
	.datab(portb27),
	.datac(porta1),
	.datad(porta7),
	.cin(gnd),
	.combout(\ShiftRight0~42_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftRight0~42 .lut_mask = 16'h5140;
defparam \ShiftRight0~42 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y37_N26
cycloneive_lcell_comb \ShiftRight0~43 (
// Equation(s):
// \ShiftRight0~43_combout  = (\portb~58_combout  & ((\porta~61_combout ))) # (!\portb~58_combout  & (\porta~55_combout ))

	.dataa(portb27),
	.datab(gnd),
	.datac(porta),
	.datad(porta3),
	.cin(gnd),
	.combout(\ShiftRight0~43_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftRight0~43 .lut_mask = 16'hFA50;
defparam \ShiftRight0~43 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X52_Y35_N4
cycloneive_lcell_comb \ShiftRight0~44 (
// Equation(s):
// \ShiftRight0~44_combout  = (!\portb~62_combout  & ((\ShiftRight0~42_combout ) # ((\portb~60_combout  & \ShiftRight0~43_combout ))))

	.dataa(portb28),
	.datab(portb29),
	.datac(\ShiftRight0~43_combout ),
	.datad(\ShiftRight0~42_combout ),
	.cin(gnd),
	.combout(\ShiftRight0~44_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftRight0~44 .lut_mask = 16'h3320;
defparam \ShiftRight0~44 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X52_Y35_N30
cycloneive_lcell_comb \ShiftRight0~48 (
// Equation(s):
// \ShiftRight0~48_combout  = (!\portb~64_combout  & ((\ShiftRight0~44_combout ) # ((\portb~62_combout  & \ShiftRight0~47_combout ))))

	.dataa(portb30),
	.datab(portb29),
	.datac(\ShiftRight0~44_combout ),
	.datad(\ShiftRight0~47_combout ),
	.cin(gnd),
	.combout(\ShiftRight0~48_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftRight0~48 .lut_mask = 16'h5450;
defparam \ShiftRight0~48 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X52_Y40_N16
cycloneive_lcell_comb \Selector0~14 (
// Equation(s):
// \Selector0~14_combout  = (!plif_idexaluop_l_1 & (!plif_idexaluop_l_0 & (!plif_idexaluop_l_2 & !plif_idexaluop_l_3)))

	.dataa(plif_idexaluop_l_1),
	.datab(plif_idexaluop_l_0),
	.datac(plif_idexaluop_l_2),
	.datad(plif_idexaluop_l_3),
	.cin(gnd),
	.combout(\Selector0~14_combout ),
	.cout());
// synopsys translate_off
defparam \Selector0~14 .lut_mask = 16'h0001;
defparam \Selector0~14 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X52_Y40_N26
cycloneive_lcell_comb \Selector29~5 (
// Equation(s):
// \Selector29~5_combout  = (\ShiftRight0~74_combout  & (((\ShiftRight0~43_combout  & !\Selector3~1_combout )))) # (!\ShiftRight0~74_combout  & ((\ShiftRight0~85_combout ) # ((\Selector3~1_combout ))))

	.dataa(\ShiftRight0~74_combout ),
	.datab(\ShiftRight0~85_combout ),
	.datac(\ShiftRight0~43_combout ),
	.datad(\Selector3~1_combout ),
	.cin(gnd),
	.combout(\Selector29~5_combout ),
	.cout());
// synopsys translate_off
defparam \Selector29~5 .lut_mask = 16'h55E4;
defparam \Selector29~5 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y42_N22
cycloneive_lcell_comb \ShiftRight0~100 (
// Equation(s):
// \ShiftRight0~100_combout  = (\portb~62_combout  & ((\ShiftRight0~83_combout ))) # (!\portb~62_combout  & (\ShiftRight0~75_combout ))

	.dataa(gnd),
	.datab(portb29),
	.datac(\ShiftRight0~75_combout ),
	.datad(\ShiftRight0~83_combout ),
	.cin(gnd),
	.combout(\ShiftRight0~100_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftRight0~100 .lut_mask = 16'hFC30;
defparam \ShiftRight0~100 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y38_N20
cycloneive_lcell_comb \Selector20~2 (
// Equation(s):
// \Selector20~2_combout  = (\porta~101_combout  & ((\portb~44_combout  & (\Selector0~11_combout )) # (!\portb~44_combout  & ((\Selector0~13_combout ))))) # (!\porta~101_combout  & (((\Selector0~13_combout ) # (!\portb~44_combout ))))

	.dataa(\Selector0~11_combout ),
	.datab(\Selector0~13_combout ),
	.datac(porta17),
	.datad(portb20),
	.cin(gnd),
	.combout(\Selector20~2_combout ),
	.cout());
// synopsys translate_off
defparam \Selector20~2 .lut_mask = 16'hACCF;
defparam \Selector20~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X50_Y39_N12
cycloneive_lcell_comb \Selector21~3 (
// Equation(s):
// \Selector21~3_combout  = (\Selector0~13_combout  & (\porta~102_combout  $ (\portb~46_combout )))

	.dataa(\Selector0~13_combout ),
	.datab(porta18),
	.datac(gnd),
	.datad(portb21),
	.cin(gnd),
	.combout(\Selector21~3_combout ),
	.cout());
// synopsys translate_off
defparam \Selector21~3 .lut_mask = 16'h2288;
defparam \Selector21~3 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y38_N12
cycloneive_lcell_comb \Selector18~3 (
// Equation(s):
// \Selector18~3_combout  = (\ShiftRight0~74_combout  & (\portb~66_combout  & (plif_idexaluop_l_0 & \Selector1~3_combout )))

	.dataa(\ShiftRight0~74_combout ),
	.datab(portb31),
	.datac(plif_idexaluop_l_0),
	.datad(\Selector1~3_combout ),
	.cin(gnd),
	.combout(\Selector18~3_combout ),
	.cout());
// synopsys translate_off
defparam \Selector18~3 .lut_mask = 16'h8000;
defparam \Selector18~3 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X50_Y40_N22
cycloneive_lcell_comb \Selector19~2 (
// Equation(s):
// \Selector19~2_combout  = (\porta~100_combout  & (\Selector0~11_combout )) # (!\porta~100_combout  & ((\Selector0~12_combout )))

	.dataa(\Selector0~11_combout ),
	.datab(porta16),
	.datac(\Selector0~12_combout ),
	.datad(gnd),
	.cin(gnd),
	.combout(\Selector19~2_combout ),
	.cout());
// synopsys translate_off
defparam \Selector19~2 .lut_mask = 16'hB8B8;
defparam \Selector19~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X50_Y35_N22
cycloneive_lcell_comb \Selector14~1 (
// Equation(s):
// \Selector14~1_combout  = (\porta~118_combout  & (((\Selector0~10_combout )))) # (!\porta~118_combout  & (\Selector0~12_combout  & ((!\portb~32_combout ))))

	.dataa(\Selector0~12_combout ),
	.datab(\Selector0~10_combout ),
	.datac(porta34),
	.datad(portb14),
	.cin(gnd),
	.combout(\Selector14~1_combout ),
	.cout());
// synopsys translate_off
defparam \Selector14~1 .lut_mask = 16'hC0CA;
defparam \Selector14~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y37_N10
cycloneive_lcell_comb \Selector13~4 (
// Equation(s):
// \Selector13~4_combout  = (\Selector0~10_combout ) # ((\Selector0~11_combout  & \porta~117_combout ))

	.dataa(\Selector0~11_combout ),
	.datab(\Selector0~10_combout ),
	.datac(gnd),
	.datad(porta33),
	.cin(gnd),
	.combout(\Selector13~4_combout ),
	.cout());
// synopsys translate_off
defparam \Selector13~4 .lut_mask = 16'hEECC;
defparam \Selector13~4 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y40_N30
cycloneive_lcell_comb \Selector11~2 (
// Equation(s):
// \Selector11~2_combout  = (!plif_idexaluop_l_0 & (\ShiftLeft0~65_combout  & \Selector0~18_combout ))

	.dataa(gnd),
	.datab(plif_idexaluop_l_0),
	.datac(\ShiftLeft0~65_combout ),
	.datad(\Selector0~18_combout ),
	.cin(gnd),
	.combout(\Selector11~2_combout ),
	.cout());
// synopsys translate_off
defparam \Selector11~2 .lut_mask = 16'h3000;
defparam \Selector11~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X50_Y40_N26
cycloneive_lcell_comb \Selector8~6 (
// Equation(s):
// \Selector8~6_combout  = (\porta~112_combout  & (\Selector0~11_combout )) # (!\porta~112_combout  & ((\Selector0~12_combout )))

	.dataa(\Selector0~11_combout ),
	.datab(porta28),
	.datac(\Selector0~12_combout ),
	.datad(gnd),
	.cin(gnd),
	.combout(\Selector8~6_combout ),
	.cout());
// synopsys translate_off
defparam \Selector8~6 .lut_mask = 16'hB8B8;
defparam \Selector8~6 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y39_N0
cycloneive_lcell_comb \Selector9~3 (
// Equation(s):
// \Selector9~3_combout  = (\porta~113_combout  & (\Selector0~10_combout )) # (!\porta~113_combout  & (((\Selector0~12_combout  & !\portb~22_combout ))))

	.dataa(\Selector0~10_combout ),
	.datab(\Selector0~12_combout ),
	.datac(portb9),
	.datad(porta29),
	.cin(gnd),
	.combout(\Selector9~3_combout ),
	.cout());
// synopsys translate_off
defparam \Selector9~3 .lut_mask = 16'hAA0C;
defparam \Selector9~3 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y39_N10
cycloneive_lcell_comb \Selector9~4 (
// Equation(s):
// \Selector9~4_combout  = (\Selector9~3_combout ) # ((\Selector0~13_combout  & (\portb~22_combout  $ (\porta~113_combout ))))

	.dataa(\Selector0~13_combout ),
	.datab(\Selector9~3_combout ),
	.datac(portb9),
	.datad(porta29),
	.cin(gnd),
	.combout(\Selector9~4_combout ),
	.cout());
// synopsys translate_off
defparam \Selector9~4 .lut_mask = 16'hCEEC;
defparam \Selector9~4 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X52_Y36_N22
cycloneive_lcell_comb \ShiftLeft0~72 (
// Equation(s):
// \ShiftLeft0~72_combout  = (\portb~58_combout  & (\porta~112_combout )) # (!\portb~58_combout  & ((\porta~111_combout )))

	.dataa(porta28),
	.datab(gnd),
	.datac(porta27),
	.datad(portb27),
	.cin(gnd),
	.combout(\ShiftLeft0~72_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftLeft0~72 .lut_mask = 16'hAAF0;
defparam \ShiftLeft0~72 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X52_Y42_N4
cycloneive_lcell_comb \ShiftLeft0~79 (
// Equation(s):
// \ShiftLeft0~79_combout  = (\portb~58_combout  & (\porta~108_combout )) # (!\portb~58_combout  & ((\porta~107_combout )))

	.dataa(porta24),
	.datab(gnd),
	.datac(portb27),
	.datad(porta23),
	.cin(gnd),
	.combout(\ShiftLeft0~79_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftLeft0~79 .lut_mask = 16'hAFA0;
defparam \ShiftLeft0~79 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X52_Y39_N22
cycloneive_lcell_comb \WideOr1~5 (
// Equation(s):
// \WideOr1~5_combout  = (Selector29) # ((Selector28) # (Selector24))

	.dataa(Selector29),
	.datab(gnd),
	.datac(Selector28),
	.datad(Selector24),
	.cin(gnd),
	.combout(\WideOr1~5_combout ),
	.cout());
// synopsys translate_off
defparam \WideOr1~5 .lut_mask = 16'hFFFA;
defparam \WideOr1~5 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y39_N8
cycloneive_lcell_comb \Selector30~8 (
// Equation(s):
// Selector30 = (\Selector30~0_combout ) # (\Selector30~7_combout )

	.dataa(gnd),
	.datab(\Selector30~0_combout ),
	.datac(gnd),
	.datad(\Selector30~7_combout ),
	.cin(gnd),
	.combout(Selector30),
	.cout());
// synopsys translate_off
defparam \Selector30~8 .lut_mask = 16'hFFCC;
defparam \Selector30~8 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X50_Y39_N0
cycloneive_lcell_comb \Selector31~8 (
// Equation(s):
// Selector31 = (\Selector31~4_combout ) # ((\Selector31~7_combout ) # ((\Selector31~2_combout ) # (\Selector31~0_combout )))

	.dataa(\Selector31~4_combout ),
	.datab(\Selector31~7_combout ),
	.datac(\Selector31~2_combout ),
	.datad(\Selector31~0_combout ),
	.cin(gnd),
	.combout(Selector31),
	.cout());
// synopsys translate_off
defparam \Selector31~8 .lut_mask = 16'hFFFE;
defparam \Selector31~8 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X52_Y40_N20
cycloneive_lcell_comb \Selector28~10 (
// Equation(s):
// Selector28 = (\Selector28~4_combout ) # ((\Selector28~9_combout ) # ((\Selector23~1_combout  & \ShiftRight0~84_combout )))

	.dataa(\Selector23~1_combout ),
	.datab(\Selector28~4_combout ),
	.datac(\ShiftRight0~84_combout ),
	.datad(\Selector28~9_combout ),
	.cin(gnd),
	.combout(Selector28),
	.cout());
// synopsys translate_off
defparam \Selector28~10 .lut_mask = 16'hFFEC;
defparam \Selector28~10 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X52_Y40_N30
cycloneive_lcell_comb \Selector29~8 (
// Equation(s):
// Selector29 = (\Selector29~0_combout ) # ((\Selector29~7_combout ) # ((\Selector23~1_combout  & \ShiftRight0~93_combout )))

	.dataa(\Selector23~1_combout ),
	.datab(\Selector29~0_combout ),
	.datac(\ShiftRight0~93_combout ),
	.datad(\Selector29~7_combout ),
	.cin(gnd),
	.combout(Selector29),
	.cout());
// synopsys translate_off
defparam \Selector29~8 .lut_mask = 16'hFFEC;
defparam \Selector29~8 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X50_Y41_N24
cycloneive_lcell_comb \Selector26~8 (
// Equation(s):
// Selector26 = (\Selector26~5_combout ) # ((\Selector26~7_combout ) # ((\Selector26~0_combout ) # (\Selector26~4_combout )))

	.dataa(\Selector26~5_combout ),
	.datab(\Selector26~7_combout ),
	.datac(\Selector26~0_combout ),
	.datad(\Selector26~4_combout ),
	.cin(gnd),
	.combout(Selector26),
	.cout());
// synopsys translate_off
defparam \Selector26~8 .lut_mask = 16'hFFFE;
defparam \Selector26~8 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X50_Y38_N26
cycloneive_lcell_comb \Selector27~8 (
// Equation(s):
// Selector27 = (\Selector27~0_combout ) # ((\Selector27~5_combout ) # ((\Selector27~7_combout ) # (\Selector27~4_combout )))

	.dataa(\Selector27~0_combout ),
	.datab(\Selector27~5_combout ),
	.datac(\Selector27~7_combout ),
	.datad(\Selector27~4_combout ),
	.cin(gnd),
	.combout(Selector27),
	.cout());
// synopsys translate_off
defparam \Selector27~8 .lut_mask = 16'hFFFE;
defparam \Selector27~8 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y42_N4
cycloneive_lcell_comb \Selector24~9 (
// Equation(s):
// Selector24 = (\Selector24~6_combout ) # ((\Selector24~8_combout ) # ((\Selector24~5_combout ) # (\Selector24~1_combout )))

	.dataa(\Selector24~6_combout ),
	.datab(\Selector24~8_combout ),
	.datac(\Selector24~5_combout ),
	.datad(\Selector24~1_combout ),
	.cin(gnd),
	.combout(Selector24),
	.cout());
// synopsys translate_off
defparam \Selector24~9 .lut_mask = 16'hFFFE;
defparam \Selector24~9 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y39_N14
cycloneive_lcell_comb \Selector25~7 (
// Equation(s):
// Selector25 = (\Selector25~6_combout ) # ((\Selector25~3_combout ) # ((\Selector24~10_combout  & \ShiftLeft0~20_combout )))

	.dataa(\Selector24~10_combout ),
	.datab(\ShiftLeft0~20_combout ),
	.datac(\Selector25~6_combout ),
	.datad(\Selector25~3_combout ),
	.cin(gnd),
	.combout(Selector25),
	.cout());
// synopsys translate_off
defparam \Selector25~7 .lut_mask = 16'hFFF8;
defparam \Selector25~7 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y41_N12
cycloneive_lcell_comb \Selector22~8 (
// Equation(s):
// Selector22 = (\Selector22~1_combout ) # ((\Selector22~7_combout ) # ((\Selector0~9_combout  & \Add0~18_combout )))

	.dataa(\Selector0~9_combout ),
	.datab(\Add0~18_combout ),
	.datac(\Selector22~1_combout ),
	.datad(\Selector22~7_combout ),
	.cin(gnd),
	.combout(Selector22),
	.cout());
// synopsys translate_off
defparam \Selector22~8 .lut_mask = 16'hFFF8;
defparam \Selector22~8 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y40_N6
cycloneive_lcell_comb \Selector23~9 (
// Equation(s):
// Selector23 = (\Selector23~7_combout ) # ((\Selector23~8_combout ) # ((\Selector16~0_combout  & \ShiftLeft0~80_combout )))

	.dataa(\Selector16~0_combout ),
	.datab(\ShiftLeft0~80_combout ),
	.datac(\Selector23~7_combout ),
	.datad(\Selector23~8_combout ),
	.cin(gnd),
	.combout(Selector23),
	.cout());
// synopsys translate_off
defparam \Selector23~9 .lut_mask = 16'hFFF8;
defparam \Selector23~9 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y37_N4
cycloneive_lcell_comb \Selector20~9 (
// Equation(s):
// Selector20 = (\Selector20~8_combout ) # ((\Selector20~7_combout ) # ((\ShiftLeft0~32_combout  & \Selector16~0_combout )))

	.dataa(\ShiftLeft0~32_combout ),
	.datab(\Selector16~0_combout ),
	.datac(\Selector20~8_combout ),
	.datad(\Selector20~7_combout ),
	.cin(gnd),
	.combout(Selector20),
	.cout());
// synopsys translate_off
defparam \Selector20~9 .lut_mask = 16'hFFF8;
defparam \Selector20~9 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y37_N0
cycloneive_lcell_comb \Selector21~8 (
// Equation(s):
// Selector21 = (\Selector21~7_combout ) # ((\Selector21~6_combout ) # ((\ShiftLeft0~36_combout  & \Selector16~0_combout )))

	.dataa(\ShiftLeft0~36_combout ),
	.datab(\Selector16~0_combout ),
	.datac(\Selector21~7_combout ),
	.datad(\Selector21~6_combout ),
	.cin(gnd),
	.combout(Selector21),
	.cout());
// synopsys translate_off
defparam \Selector21~8 .lut_mask = 16'hFFF8;
defparam \Selector21~8 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y38_N0
cycloneive_lcell_comb \Selector18~9 (
// Equation(s):
// Selector18 = (\Selector18~8_combout ) # ((\Selector18~5_combout ) # ((\Selector0~9_combout  & \Add0~26_combout )))

	.dataa(\Selector0~9_combout ),
	.datab(\Selector18~8_combout ),
	.datac(\Add0~26_combout ),
	.datad(\Selector18~5_combout ),
	.cin(gnd),
	.combout(Selector18),
	.cout());
// synopsys translate_off
defparam \Selector18~9 .lut_mask = 16'hFFEC;
defparam \Selector18~9 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y40_N30
cycloneive_lcell_comb \Selector19~8 (
// Equation(s):
// Selector19 = (\Selector19~6_combout ) # ((\Selector19~0_combout ) # ((\Selector19~5_combout ) # (\Selector19~7_combout )))

	.dataa(\Selector19~6_combout ),
	.datab(\Selector19~0_combout ),
	.datac(\Selector19~5_combout ),
	.datad(\Selector19~7_combout ),
	.cin(gnd),
	.combout(Selector19),
	.cout());
// synopsys translate_off
defparam \Selector19~8 .lut_mask = 16'hFFFE;
defparam \Selector19~8 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X52_Y36_N26
cycloneive_lcell_comb \Selector16~10 (
// Equation(s):
// Selector16 = (\Selector16~4_combout ) # ((\Selector16~9_combout ) # ((\Selector0~8_combout  & \Add1~30_combout )))

	.dataa(\Selector0~8_combout ),
	.datab(\Add1~30_combout ),
	.datac(\Selector16~4_combout ),
	.datad(\Selector16~9_combout ),
	.cin(gnd),
	.combout(Selector16),
	.cout());
// synopsys translate_off
defparam \Selector16~10 .lut_mask = 16'hFFF8;
defparam \Selector16~10 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y39_N4
cycloneive_lcell_comb \Selector17~7 (
// Equation(s):
// Selector17 = (\Selector17~6_combout ) # ((\Selector17~3_combout ) # ((\Selector0~9_combout  & \Add0~28_combout )))

	.dataa(\Selector0~9_combout ),
	.datab(\Add0~28_combout ),
	.datac(\Selector17~6_combout ),
	.datad(\Selector17~3_combout ),
	.cin(gnd),
	.combout(Selector17),
	.cout());
// synopsys translate_off
defparam \Selector17~7 .lut_mask = 16'hFFF8;
defparam \Selector17~7 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y41_N14
cycloneive_lcell_comb \Selector14~8 (
// Equation(s):
// Selector14 = (\Selector14~7_combout ) # ((\Selector14~5_combout ) # ((\Selector0~9_combout  & \Add0~34_combout )))

	.dataa(\Selector14~7_combout ),
	.datab(\Selector0~9_combout ),
	.datac(\Add0~34_combout ),
	.datad(\Selector14~5_combout ),
	.cin(gnd),
	.combout(Selector14),
	.cout());
// synopsys translate_off
defparam \Selector14~8 .lut_mask = 16'hFFEA;
defparam \Selector14~8 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X52_Y35_N18
cycloneive_lcell_comb \Selector15~8 (
// Equation(s):
// Selector15 = (\Selector15~0_combout ) # ((\Selector15~7_combout ) # ((\Selector8~1_combout  & \ShiftRight0~70_combout )))

	.dataa(\Selector8~1_combout ),
	.datab(\Selector15~0_combout ),
	.datac(\ShiftRight0~70_combout ),
	.datad(\Selector15~7_combout ),
	.cin(gnd),
	.combout(Selector15),
	.cout());
// synopsys translate_off
defparam \Selector15~8 .lut_mask = 16'hFFEC;
defparam \Selector15~8 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y37_N28
cycloneive_lcell_comb \Selector12~10 (
// Equation(s):
// Selector12 = (\Selector12~9_combout ) # ((\Selector12~2_combout ) # ((\Selector12~7_combout ) # (\Selector12~8_combout )))

	.dataa(\Selector12~9_combout ),
	.datab(\Selector12~2_combout ),
	.datac(\Selector12~7_combout ),
	.datad(\Selector12~8_combout ),
	.cin(gnd),
	.combout(Selector12),
	.cout());
// synopsys translate_off
defparam \Selector12~10 .lut_mask = 16'hFFFE;
defparam \Selector12~10 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y37_N8
cycloneive_lcell_comb \Selector13~8 (
// Equation(s):
// Selector13 = (\Selector13~7_combout ) # ((\Selector13~0_combout ) # ((\Add1~36_combout  & \Selector0~8_combout )))

	.dataa(\Add1~36_combout ),
	.datab(\Selector0~8_combout ),
	.datac(\Selector13~7_combout ),
	.datad(\Selector13~0_combout ),
	.cin(gnd),
	.combout(Selector13),
	.cout());
// synopsys translate_off
defparam \Selector13~8 .lut_mask = 16'hFFF8;
defparam \Selector13~8 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y42_N28
cycloneive_lcell_comb \Selector10~8 (
// Equation(s):
// Selector10 = (\Selector10~1_combout ) # ((\Selector10~7_combout ) # ((\Selector0~9_combout  & \Add0~42_combout )))

	.dataa(\Selector0~9_combout ),
	.datab(\Selector10~1_combout ),
	.datac(\Add0~42_combout ),
	.datad(\Selector10~7_combout ),
	.cin(gnd),
	.combout(Selector10),
	.cout());
// synopsys translate_off
defparam \Selector10~8 .lut_mask = 16'hFFEC;
defparam \Selector10~8 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y39_N6
cycloneive_lcell_comb \Selector11~9 (
// Equation(s):
// Selector11 = (\Selector11~5_combout ) # ((\Selector11~8_combout ) # ((\Add0~40_combout  & \Selector0~9_combout )))

	.dataa(\Add0~40_combout ),
	.datab(\Selector0~9_combout ),
	.datac(\Selector11~5_combout ),
	.datad(\Selector11~8_combout ),
	.cin(gnd),
	.combout(Selector11),
	.cout());
// synopsys translate_off
defparam \Selector11~9 .lut_mask = 16'hFFF8;
defparam \Selector11~9 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X52_Y39_N14
cycloneive_lcell_comb \Selector8~10 (
// Equation(s):
// Selector8 = (\Selector8~9_combout ) # ((\Selector8~5_combout ) # ((\Add1~46_combout  & \Selector0~8_combout )))

	.dataa(\Selector8~9_combout ),
	.datab(\Add1~46_combout ),
	.datac(\Selector0~8_combout ),
	.datad(\Selector8~5_combout ),
	.cin(gnd),
	.combout(Selector8),
	.cout());
// synopsys translate_off
defparam \Selector8~10 .lut_mask = 16'hFFEA;
defparam \Selector8~10 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X52_Y39_N28
cycloneive_lcell_comb \Selector9~8 (
// Equation(s):
// Selector9 = (\Selector9~1_combout ) # ((\Selector9~7_combout ) # ((\Selector0~8_combout  & \Add1~44_combout )))

	.dataa(\Selector0~8_combout ),
	.datab(\Selector9~1_combout ),
	.datac(\Add1~44_combout ),
	.datad(\Selector9~7_combout ),
	.cin(gnd),
	.combout(Selector9),
	.cout());
// synopsys translate_off
defparam \Selector9~8 .lut_mask = 16'hFFEC;
defparam \Selector9~8 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y36_N0
cycloneive_lcell_comb \Selector6~8 (
// Equation(s):
// Selector6 = (\Selector6~7_combout ) # ((\Selector6~6_combout ) # ((\Selector0~6_combout  & \Add1~50_combout )))

	.dataa(\Selector0~6_combout ),
	.datab(\Add1~50_combout ),
	.datac(\Selector6~7_combout ),
	.datad(\Selector6~6_combout ),
	.cin(gnd),
	.combout(Selector6),
	.cout());
// synopsys translate_off
defparam \Selector6~8 .lut_mask = 16'hFFF8;
defparam \Selector6~8 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y35_N12
cycloneive_lcell_comb \Selector7~11 (
// Equation(s):
// Selector7 = (\Selector7~10_combout ) # ((\Selector7~7_combout ) # ((\Selector0~5_combout  & \Add0~48_combout )))

	.dataa(\Selector7~10_combout ),
	.datab(\Selector0~5_combout ),
	.datac(\Add0~48_combout ),
	.datad(\Selector7~7_combout ),
	.cin(gnd),
	.combout(Selector7),
	.cout());
// synopsys translate_off
defparam \Selector7~11 .lut_mask = 16'hFFEA;
defparam \Selector7~11 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y36_N30
cycloneive_lcell_comb \Selector4~10 (
// Equation(s):
// Selector4 = (\Selector4~9_combout ) # ((\Selector4~6_combout ) # ((\Selector0~6_combout  & \Add1~54_combout )))

	.dataa(\Selector0~6_combout ),
	.datab(\Selector4~9_combout ),
	.datac(\Add1~54_combout ),
	.datad(\Selector4~6_combout ),
	.cin(gnd),
	.combout(Selector4),
	.cout());
// synopsys translate_off
defparam \Selector4~10 .lut_mask = 16'hFFEC;
defparam \Selector4~10 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y36_N26
cycloneive_lcell_comb \Selector5~8 (
// Equation(s):
// Selector5 = (\Selector5~6_combout ) # ((\Selector5~7_combout ) # ((\Add0~52_combout  & \Selector0~5_combout )))

	.dataa(\Add0~52_combout ),
	.datab(\Selector0~5_combout ),
	.datac(\Selector5~6_combout ),
	.datad(\Selector5~7_combout ),
	.cin(gnd),
	.combout(Selector5),
	.cout());
// synopsys translate_off
defparam \Selector5~8 .lut_mask = 16'hFFF8;
defparam \Selector5~8 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X50_Y39_N20
cycloneive_lcell_comb \Selector2~11 (
// Equation(s):
// Selector2 = (\Selector2~10_combout ) # ((\Selector2~9_combout ) # ((\Selector0~8_combout  & \Add1~58_combout )))

	.dataa(\Selector0~8_combout ),
	.datab(\Add1~58_combout ),
	.datac(\Selector2~10_combout ),
	.datad(\Selector2~9_combout ),
	.cin(gnd),
	.combout(Selector2),
	.cout());
// synopsys translate_off
defparam \Selector2~11 .lut_mask = 16'hFFF8;
defparam \Selector2~11 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X50_Y39_N8
cycloneive_lcell_comb \Selector3~11 (
// Equation(s):
// Selector3 = (\Selector3~10_combout ) # ((\Selector3~9_combout ) # ((\Selector0~8_combout  & \Add1~56_combout )))

	.dataa(\Selector0~8_combout ),
	.datab(\Selector3~10_combout ),
	.datac(\Add1~56_combout ),
	.datad(\Selector3~9_combout ),
	.cin(gnd),
	.combout(Selector3),
	.cout());
// synopsys translate_off
defparam \Selector3~11 .lut_mask = 16'hFFEC;
defparam \Selector3~11 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X52_Y42_N24
cycloneive_lcell_comb \Selector0~34 (
// Equation(s):
// Selector0 = (\Selector0~23_combout ) # ((\Selector0~26_combout ) # ((\Selector0~33_combout ) # (\Selector0~22_combout )))

	.dataa(\Selector0~23_combout ),
	.datab(\Selector0~26_combout ),
	.datac(\Selector0~33_combout ),
	.datad(\Selector0~22_combout ),
	.cin(gnd),
	.combout(Selector0),
	.cout());
// synopsys translate_off
defparam \Selector0~34 .lut_mask = 16'hFFFE;
defparam \Selector0~34 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y42_N14
cycloneive_lcell_comb \Selector1~20 (
// Equation(s):
// Selector1 = (\Selector1~8_combout ) # ((\Selector1~19_combout ) # ((\Selector0~9_combout  & \Add0~60_combout )))

	.dataa(\Selector0~9_combout ),
	.datab(\Selector1~8_combout ),
	.datac(\Add0~60_combout ),
	.datad(\Selector1~19_combout ),
	.cin(gnd),
	.combout(Selector1),
	.cout());
// synopsys translate_off
defparam \Selector1~20 .lut_mask = 16'hFFEC;
defparam \Selector1~20 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y39_N6
cycloneive_lcell_comb WideOr1(
// Equation(s):
// WideOr11 = (!Selector1 & (!Selector0 & (!\WideOr1~0_combout  & !\WideOr1~11_combout )))

	.dataa(Selector1),
	.datab(Selector0),
	.datac(\WideOr1~0_combout ),
	.datad(\WideOr1~11_combout ),
	.cin(gnd),
	.combout(WideOr11),
	.cout());
// synopsys translate_off
defparam WideOr1.lut_mask = 16'h0001;
defparam WideOr1.sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y42_N24
cycloneive_lcell_comb \ShiftRight0~22 (
// Equation(s):
// \ShiftRight0~22_combout  = (\portb~58_combout  & (\porta~100_combout )) # (!\portb~58_combout  & ((\porta~101_combout )))

	.dataa(portb27),
	.datab(gnd),
	.datac(porta16),
	.datad(porta17),
	.cin(gnd),
	.combout(\ShiftRight0~22_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftRight0~22 .lut_mask = 16'hF5A0;
defparam \ShiftRight0~22 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X52_Y41_N28
cycloneive_lcell_comb \ShiftRight0~24 (
// Equation(s):
// \ShiftRight0~24_combout  = (\portb~60_combout  & ((\ShiftRight0~22_combout ))) # (!\portb~60_combout  & (\ShiftRight0~23_combout ))

	.dataa(\ShiftRight0~23_combout ),
	.datab(gnd),
	.datac(portb28),
	.datad(\ShiftRight0~22_combout ),
	.cin(gnd),
	.combout(\ShiftRight0~24_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftRight0~24 .lut_mask = 16'hFA0A;
defparam \ShiftRight0~24 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y41_N20
cycloneive_lcell_comb \ShiftRight0~25 (
// Equation(s):
// \ShiftRight0~25_combout  = (\portb~62_combout  & (\ShiftRight0~21_combout )) # (!\portb~62_combout  & ((\ShiftRight0~24_combout )))

	.dataa(\ShiftRight0~21_combout ),
	.datab(portb29),
	.datac(gnd),
	.datad(\ShiftRight0~24_combout ),
	.cin(gnd),
	.combout(\ShiftRight0~25_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftRight0~25 .lut_mask = 16'hBB88;
defparam \ShiftRight0~25 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y41_N6
cycloneive_lcell_comb \ShiftRight0~26 (
// Equation(s):
// \ShiftRight0~26_combout  = (!\portb~66_combout  & ((\ShiftRight0~18_combout ) # ((\portb~64_combout  & \ShiftRight0~25_combout ))))

	.dataa(\ShiftRight0~18_combout ),
	.datab(portb30),
	.datac(portb31),
	.datad(\ShiftRight0~25_combout ),
	.cin(gnd),
	.combout(\ShiftRight0~26_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftRight0~26 .lut_mask = 16'h0E0A;
defparam \ShiftRight0~26 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y38_N16
cycloneive_lcell_comb \ShiftRight0~10 (
// Equation(s):
// \ShiftRight0~10_combout  = (\portb~46_combout ) # ((\portb~50_combout ) # ((\portb~44_combout ) # (\portb~48_combout )))

	.dataa(portb21),
	.datab(portb23),
	.datac(portb20),
	.datad(portb22),
	.cin(gnd),
	.combout(\ShiftRight0~10_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftRight0~10 .lut_mask = 16'hFFFE;
defparam \ShiftRight0~10 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y38_N28
cycloneive_lcell_comb \ShiftRight0~11 (
// Equation(s):
// \ShiftRight0~11_combout  = (\portb~52_combout ) # ((\portb~54_combout ) # ((\portb~56_combout ) # (\ShiftRight0~10_combout )))

	.dataa(portb24),
	.datab(portb25),
	.datac(portb26),
	.datad(\ShiftRight0~10_combout ),
	.cin(gnd),
	.combout(\ShiftRight0~11_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftRight0~11 .lut_mask = 16'hFFFE;
defparam \ShiftRight0~11 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y38_N18
cycloneive_lcell_comb \ShiftRight0~9 (
// Equation(s):
// \ShiftRight0~9_combout  = (\portb~40_combout ) # ((\portb~36_combout ) # ((\portb~38_combout ) # (\portb~42_combout )))

	.dataa(portb18),
	.datab(portb16),
	.datac(portb17),
	.datad(portb19),
	.cin(gnd),
	.combout(\ShiftRight0~9_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftRight0~9 .lut_mask = 16'hFFFE;
defparam \ShiftRight0~9 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X52_Y40_N12
cycloneive_lcell_comb \Selector0~0 (
// Equation(s):
// \Selector0~0_combout  = (!plif_idexaluop_l_1 & (plif_idexaluop_l_0 & (!plif_idexaluop_l_2 & !plif_idexaluop_l_3)))

	.dataa(plif_idexaluop_l_1),
	.datab(plif_idexaluop_l_0),
	.datac(plif_idexaluop_l_2),
	.datad(plif_idexaluop_l_3),
	.cin(gnd),
	.combout(\Selector0~0_combout ),
	.cout());
// synopsys translate_off
defparam \Selector0~0 .lut_mask = 16'h0004;
defparam \Selector0~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y38_N10
cycloneive_lcell_comb \Selector24~0 (
// Equation(s):
// \Selector24~0_combout  = (!\ShiftRight0~8_combout  & (!\ShiftRight0~11_combout  & (!\ShiftRight0~9_combout  & \Selector0~0_combout )))

	.dataa(\ShiftRight0~8_combout ),
	.datab(\ShiftRight0~11_combout ),
	.datac(\ShiftRight0~9_combout ),
	.datad(\Selector0~0_combout ),
	.cin(gnd),
	.combout(\Selector24~0_combout ),
	.cout());
// synopsys translate_off
defparam \Selector24~0 .lut_mask = 16'h0100;
defparam \Selector24~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y41_N18
cycloneive_lcell_comb \ShiftRight0~27 (
// Equation(s):
// \ShiftRight0~27_combout  = (!\portb~58_combout  & ((\portb~60_combout  & (\porta~104_combout )) # (!\portb~60_combout  & ((\porta~105_combout )))))

	.dataa(porta20),
	.datab(portb27),
	.datac(porta21),
	.datad(portb28),
	.cin(gnd),
	.combout(\ShiftRight0~27_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftRight0~27 .lut_mask = 16'h2230;
defparam \ShiftRight0~27 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y41_N12
cycloneive_lcell_comb \ShiftRight0~28 (
// Equation(s):
// \ShiftRight0~28_combout  = (\ShiftRight0~27_combout ) # ((!\portb~60_combout  & (\portb~58_combout  & \porta~106_combout )))

	.dataa(portb28),
	.datab(portb27),
	.datac(porta22),
	.datad(\ShiftRight0~27_combout ),
	.cin(gnd),
	.combout(\ShiftRight0~28_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftRight0~28 .lut_mask = 16'hFF40;
defparam \ShiftRight0~28 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y42_N26
cycloneive_lcell_comb \ShiftRight0~30 (
// Equation(s):
// \ShiftRight0~30_combout  = (\portb~58_combout  & ((\porta~109_combout ))) # (!\portb~58_combout  & (\porta~110_combout ))

	.dataa(porta26),
	.datab(gnd),
	.datac(portb27),
	.datad(porta25),
	.cin(gnd),
	.combout(\ShiftRight0~30_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftRight0~30 .lut_mask = 16'hFA0A;
defparam \ShiftRight0~30 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y42_N20
cycloneive_lcell_comb \ShiftRight0~29 (
// Equation(s):
// \ShiftRight0~29_combout  = (\portb~58_combout  & ((\porta~107_combout ))) # (!\portb~58_combout  & (\porta~108_combout ))

	.dataa(gnd),
	.datab(portb27),
	.datac(porta24),
	.datad(porta23),
	.cin(gnd),
	.combout(\ShiftRight0~29_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftRight0~29 .lut_mask = 16'hFC30;
defparam \ShiftRight0~29 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y42_N8
cycloneive_lcell_comb \ShiftRight0~31 (
// Equation(s):
// \ShiftRight0~31_combout  = (\portb~60_combout  & ((\ShiftRight0~29_combout ))) # (!\portb~60_combout  & (\ShiftRight0~30_combout ))

	.dataa(portb28),
	.datab(gnd),
	.datac(\ShiftRight0~30_combout ),
	.datad(\ShiftRight0~29_combout ),
	.cin(gnd),
	.combout(\ShiftRight0~31_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftRight0~31 .lut_mask = 16'hFA50;
defparam \ShiftRight0~31 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y41_N16
cycloneive_lcell_comb \ShiftRight0~32 (
// Equation(s):
// \ShiftRight0~32_combout  = (\portb~62_combout  & (\ShiftRight0~28_combout )) # (!\portb~62_combout  & ((\ShiftRight0~31_combout )))

	.dataa(portb29),
	.datab(\ShiftRight0~28_combout ),
	.datac(gnd),
	.datad(\ShiftRight0~31_combout ),
	.cin(gnd),
	.combout(\ShiftRight0~32_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftRight0~32 .lut_mask = 16'hDD88;
defparam \ShiftRight0~32 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y40_N8
cycloneive_lcell_comb \ShiftRight0~36 (
// Equation(s):
// \ShiftRight0~36_combout  = (\portb~58_combout  & (\porta~115_combout )) # (!\portb~58_combout  & ((\porta~116_combout )))

	.dataa(gnd),
	.datab(portb27),
	.datac(porta31),
	.datad(porta32),
	.cin(gnd),
	.combout(\ShiftRight0~36_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftRight0~36 .lut_mask = 16'hF3C0;
defparam \ShiftRight0~36 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y40_N30
cycloneive_lcell_comb \ShiftRight0~38 (
// Equation(s):
// \ShiftRight0~38_combout  = (\portb~60_combout  & ((\ShiftRight0~36_combout ))) # (!\portb~60_combout  & (\ShiftRight0~37_combout ))

	.dataa(\ShiftRight0~37_combout ),
	.datab(gnd),
	.datac(\ShiftRight0~36_combout ),
	.datad(portb28),
	.cin(gnd),
	.combout(\ShiftRight0~38_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftRight0~38 .lut_mask = 16'hF0AA;
defparam \ShiftRight0~38 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y42_N4
cycloneive_lcell_comb \ShiftRight0~34 (
// Equation(s):
// \ShiftRight0~34_combout  = (\portb~58_combout  & ((\porta~113_combout ))) # (!\portb~58_combout  & (\porta~114_combout ))

	.dataa(gnd),
	.datab(porta30),
	.datac(portb27),
	.datad(porta29),
	.cin(gnd),
	.combout(\ShiftRight0~34_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftRight0~34 .lut_mask = 16'hFC0C;
defparam \ShiftRight0~34 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y42_N2
cycloneive_lcell_comb \ShiftRight0~33 (
// Equation(s):
// \ShiftRight0~33_combout  = (\portb~58_combout  & ((\porta~111_combout ))) # (!\portb~58_combout  & (\porta~112_combout ))

	.dataa(porta28),
	.datab(gnd),
	.datac(portb27),
	.datad(porta27),
	.cin(gnd),
	.combout(\ShiftRight0~33_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftRight0~33 .lut_mask = 16'hFA0A;
defparam \ShiftRight0~33 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y42_N30
cycloneive_lcell_comb \ShiftRight0~35 (
// Equation(s):
// \ShiftRight0~35_combout  = (\portb~60_combout  & ((\ShiftRight0~33_combout ))) # (!\portb~60_combout  & (\ShiftRight0~34_combout ))

	.dataa(portb28),
	.datab(gnd),
	.datac(\ShiftRight0~34_combout ),
	.datad(\ShiftRight0~33_combout ),
	.cin(gnd),
	.combout(\ShiftRight0~35_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftRight0~35 .lut_mask = 16'hFA50;
defparam \ShiftRight0~35 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y40_N28
cycloneive_lcell_comb \Selector22~0 (
// Equation(s):
// \Selector22~0_combout  = (\portb~62_combout  & ((\ShiftRight0~35_combout ))) # (!\portb~62_combout  & (\ShiftRight0~38_combout ))

	.dataa(gnd),
	.datab(portb29),
	.datac(\ShiftRight0~38_combout ),
	.datad(\ShiftRight0~35_combout ),
	.cin(gnd),
	.combout(\Selector22~0_combout ),
	.cout());
// synopsys translate_off
defparam \Selector22~0 .lut_mask = 16'hFC30;
defparam \Selector22~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y41_N0
cycloneive_lcell_comb \ShiftRight0~39 (
// Equation(s):
// \ShiftRight0~39_combout  = (\portb~64_combout  & (\ShiftRight0~32_combout )) # (!\portb~64_combout  & ((\Selector22~0_combout )))

	.dataa(gnd),
	.datab(\ShiftRight0~32_combout ),
	.datac(portb30),
	.datad(\Selector22~0_combout ),
	.cin(gnd),
	.combout(\ShiftRight0~39_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftRight0~39 .lut_mask = 16'hCFC0;
defparam \ShiftRight0~39 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y41_N30
cycloneive_lcell_comb \Selector30~0 (
// Equation(s):
// \Selector30~0_combout  = (\Selector24~0_combout  & ((\ShiftRight0~26_combout ) # ((\portb~66_combout  & \ShiftRight0~39_combout ))))

	.dataa(\ShiftRight0~26_combout ),
	.datab(portb31),
	.datac(\Selector24~0_combout ),
	.datad(\ShiftRight0~39_combout ),
	.cin(gnd),
	.combout(\Selector30~0_combout ),
	.cout());
// synopsys translate_off
defparam \Selector30~0 .lut_mask = 16'hE0A0;
defparam \Selector30~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y35_N18
cycloneive_lcell_comb \Selector0~3 (
// Equation(s):
// \Selector0~3_combout  = (plif_idexaluop_l_2 & (!plif_idexaluop_l_1 & (plif_idexaluop_l_0 & !plif_idexaluop_l_3)))

	.dataa(plif_idexaluop_l_2),
	.datab(plif_idexaluop_l_1),
	.datac(plif_idexaluop_l_0),
	.datad(plif_idexaluop_l_3),
	.cin(gnd),
	.combout(\Selector0~3_combout ),
	.cout());
// synopsys translate_off
defparam \Selector0~3 .lut_mask = 16'h0020;
defparam \Selector0~3 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y38_N6
cycloneive_lcell_comb \Selector0~7 (
// Equation(s):
// \Selector0~7_combout  = (plif_idexaluop_l_0 & (!plif_idexaluop_l_3 & (plif_idexaluop_l_1 & plif_idexaluop_l_2)))

	.dataa(plif_idexaluop_l_0),
	.datab(plif_idexaluop_l_3),
	.datac(plif_idexaluop_l_1),
	.datad(plif_idexaluop_l_2),
	.cin(gnd),
	.combout(\Selector0~7_combout ),
	.cout());
// synopsys translate_off
defparam \Selector0~7 .lut_mask = 16'h2000;
defparam \Selector0~7 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y41_N26
cycloneive_lcell_comb \Selector30~6 (
// Equation(s):
// \Selector30~6_combout  = (\porta~57_combout  & (\Selector0~3_combout )) # (!\porta~57_combout  & (((!\portb~60_combout  & \Selector0~7_combout ))))

	.dataa(porta1),
	.datab(\Selector0~3_combout ),
	.datac(portb28),
	.datad(\Selector0~7_combout ),
	.cin(gnd),
	.combout(\Selector30~6_combout ),
	.cout());
// synopsys translate_off
defparam \Selector30~6 .lut_mask = 16'h8D88;
defparam \Selector30~6 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y40_N6
cycloneive_lcell_comb \Selector0~4 (
// Equation(s):
// \Selector0~4_combout  = (plif_idexaluop_l_2 & (!plif_idexaluop_l_1 & (!plif_idexaluop_l_3 & !plif_idexaluop_l_0)))

	.dataa(plif_idexaluop_l_2),
	.datab(plif_idexaluop_l_1),
	.datac(plif_idexaluop_l_3),
	.datad(plif_idexaluop_l_0),
	.cin(gnd),
	.combout(\Selector0~4_combout ),
	.cout());
// synopsys translate_off
defparam \Selector0~4 .lut_mask = 16'h0002;
defparam \Selector0~4 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y41_N18
cycloneive_lcell_comb \Selector30~4 (
// Equation(s):
// \Selector30~4_combout  = (\portb~60_combout  & ((\Selector0~3_combout ) # ((\Selector0~4_combout  & \porta~57_combout ))))

	.dataa(\Selector0~3_combout ),
	.datab(portb28),
	.datac(\Selector0~4_combout ),
	.datad(porta1),
	.cin(gnd),
	.combout(\Selector30~4_combout ),
	.cout());
// synopsys translate_off
defparam \Selector30~4 .lut_mask = 16'hC888;
defparam \Selector30~4 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X52_Y40_N10
cycloneive_lcell_comb \Selector0~2 (
// Equation(s):
// \Selector0~2_combout  = (plif_idexaluop_l_1 & (!plif_idexaluop_l_0 & (plif_idexaluop_l_2 & !plif_idexaluop_l_3)))

	.dataa(plif_idexaluop_l_1),
	.datab(plif_idexaluop_l_0),
	.datac(plif_idexaluop_l_2),
	.datad(plif_idexaluop_l_3),
	.cin(gnd),
	.combout(\Selector0~2_combout ),
	.cout());
// synopsys translate_off
defparam \Selector0~2 .lut_mask = 16'h0020;
defparam \Selector0~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y41_N28
cycloneive_lcell_comb \ShiftLeft0~2 (
// Equation(s):
// \ShiftLeft0~2_combout  = (\portb~58_combout  & (\porta~91_combout )) # (!\portb~58_combout  & ((\porta~57_combout )))

	.dataa(gnd),
	.datab(portb27),
	.datac(porta7),
	.datad(porta1),
	.cin(gnd),
	.combout(\ShiftLeft0~2_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftLeft0~2 .lut_mask = 16'hF3C0;
defparam \ShiftLeft0~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y39_N6
cycloneive_lcell_comb \Selector1~0 (
// Equation(s):
// \Selector1~0_combout  = (\portb~60_combout ) # (\portb~62_combout )

	.dataa(portb28),
	.datab(gnd),
	.datac(gnd),
	.datad(portb29),
	.cin(gnd),
	.combout(\Selector1~0_combout ),
	.cout());
// synopsys translate_off
defparam \Selector1~0 .lut_mask = 16'hFFAA;
defparam \Selector1~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y38_N8
cycloneive_lcell_comb \Selector0~1 (
// Equation(s):
// \Selector0~1_combout  = (!plif_idexaluop_l_0 & (!plif_idexaluop_l_2 & (!plif_idexaluop_l_1 & !plif_idexaluop_l_3)))

	.dataa(plif_idexaluop_l_0),
	.datab(plif_idexaluop_l_2),
	.datac(plif_idexaluop_l_1),
	.datad(plif_idexaluop_l_3),
	.cin(gnd),
	.combout(\Selector0~1_combout ),
	.cout());
// synopsys translate_off
defparam \Selector0~1 .lut_mask = 16'h0001;
defparam \Selector0~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y38_N10
cycloneive_lcell_comb \ShiftRight0~40 (
// Equation(s):
// \ShiftRight0~40_combout  = (\portb~54_combout ) # ((\portb~56_combout ) # (\portb~52_combout ))

	.dataa(portb25),
	.datab(gnd),
	.datac(portb26),
	.datad(portb24),
	.cin(gnd),
	.combout(\ShiftRight0~40_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftRight0~40 .lut_mask = 16'hFFFA;
defparam \ShiftRight0~40 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y38_N22
cycloneive_lcell_comb \ShiftRight0~41 (
// Equation(s):
// \ShiftRight0~41_combout  = (\ShiftRight0~9_combout ) # ((\ShiftRight0~40_combout ) # (\ShiftRight0~10_combout ))

	.dataa(gnd),
	.datab(\ShiftRight0~9_combout ),
	.datac(\ShiftRight0~40_combout ),
	.datad(\ShiftRight0~10_combout ),
	.cin(gnd),
	.combout(\ShiftRight0~41_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftRight0~41 .lut_mask = 16'hFFFC;
defparam \ShiftRight0~41 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y41_N10
cycloneive_lcell_comb \Selector30~1 (
// Equation(s):
// \Selector30~1_combout  = (!\ShiftRight0~8_combout  & (\Selector0~1_combout  & (!\portb~66_combout  & !\ShiftRight0~41_combout )))

	.dataa(\ShiftRight0~8_combout ),
	.datab(\Selector0~1_combout ),
	.datac(portb31),
	.datad(\ShiftRight0~41_combout ),
	.cin(gnd),
	.combout(\Selector30~1_combout ),
	.cout());
// synopsys translate_off
defparam \Selector30~1 .lut_mask = 16'h0004;
defparam \Selector30~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y41_N6
cycloneive_lcell_comb \Selector30~2 (
// Equation(s):
// \Selector30~2_combout  = (!\portb~64_combout  & (\ShiftLeft0~2_combout  & (!\Selector1~0_combout  & \Selector30~1_combout )))

	.dataa(portb30),
	.datab(\ShiftLeft0~2_combout ),
	.datac(\Selector1~0_combout ),
	.datad(\Selector30~1_combout ),
	.cin(gnd),
	.combout(\Selector30~2_combout ),
	.cout());
// synopsys translate_off
defparam \Selector30~2 .lut_mask = 16'h0400;
defparam \Selector30~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y41_N0
cycloneive_lcell_comb \Selector30~3 (
// Equation(s):
// \Selector30~3_combout  = (\Selector30~2_combout ) # ((\Selector0~2_combout  & (\porta~57_combout  $ (\portb~60_combout ))))

	.dataa(porta1),
	.datab(portb28),
	.datac(\Selector0~2_combout ),
	.datad(\Selector30~2_combout ),
	.cin(gnd),
	.combout(\Selector30~3_combout ),
	.cout());
// synopsys translate_off
defparam \Selector30~3 .lut_mask = 16'hFF60;
defparam \Selector30~3 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X50_Y35_N0
cycloneive_lcell_comb \Selector0~5 (
// Equation(s):
// \Selector0~5_combout  = (!plif_idexaluop_l_3 & (plif_idexaluop_l_1 & (!plif_idexaluop_l_2 & !plif_idexaluop_l_0)))

	.dataa(plif_idexaluop_l_3),
	.datab(plif_idexaluop_l_1),
	.datac(plif_idexaluop_l_2),
	.datad(plif_idexaluop_l_0),
	.cin(gnd),
	.combout(\Selector0~5_combout ),
	.cout());
// synopsys translate_off
defparam \Selector0~5 .lut_mask = 16'h0004;
defparam \Selector0~5 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X50_Y35_N30
cycloneive_lcell_comb \Selector0~6 (
// Equation(s):
// \Selector0~6_combout  = (!plif_idexaluop_l_3 & (plif_idexaluop_l_1 & (!plif_idexaluop_l_2 & plif_idexaluop_l_0)))

	.dataa(plif_idexaluop_l_3),
	.datab(plif_idexaluop_l_1),
	.datac(plif_idexaluop_l_2),
	.datad(plif_idexaluop_l_0),
	.cin(gnd),
	.combout(\Selector0~6_combout ),
	.cout());
// synopsys translate_off
defparam \Selector0~6 .lut_mask = 16'h0400;
defparam \Selector0~6 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X52_Y38_N0
cycloneive_lcell_comb \Add0~0 (
// Equation(s):
// \Add0~0_combout  = (\porta~91_combout  & (\portb~58_combout  $ (VCC))) # (!\porta~91_combout  & (\portb~58_combout  & VCC))
// \Add0~1  = CARRY((\porta~91_combout  & \portb~58_combout ))

	.dataa(porta7),
	.datab(portb27),
	.datac(gnd),
	.datad(vcc),
	.cin(gnd),
	.combout(\Add0~0_combout ),
	.cout(\Add0~1 ));
// synopsys translate_off
defparam \Add0~0 .lut_mask = 16'h6688;
defparam \Add0~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X52_Y38_N2
cycloneive_lcell_comb \Add0~2 (
// Equation(s):
// \Add0~2_combout  = (\portb~60_combout  & ((\porta~57_combout  & (\Add0~1  & VCC)) # (!\porta~57_combout  & (!\Add0~1 )))) # (!\portb~60_combout  & ((\porta~57_combout  & (!\Add0~1 )) # (!\porta~57_combout  & ((\Add0~1 ) # (GND)))))
// \Add0~3  = CARRY((\portb~60_combout  & (!\porta~57_combout  & !\Add0~1 )) # (!\portb~60_combout  & ((!\Add0~1 ) # (!\porta~57_combout ))))

	.dataa(portb28),
	.datab(porta1),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add0~1 ),
	.combout(\Add0~2_combout ),
	.cout(\Add0~3 ));
// synopsys translate_off
defparam \Add0~2 .lut_mask = 16'h9617;
defparam \Add0~2 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X54_Y41_N24
cycloneive_lcell_comb \Selector30~5 (
// Equation(s):
// \Selector30~5_combout  = (\Add1~2_combout  & ((\Selector0~6_combout ) # ((\Selector0~5_combout  & \Add0~2_combout )))) # (!\Add1~2_combout  & (\Selector0~5_combout  & ((\Add0~2_combout ))))

	.dataa(\Add1~2_combout ),
	.datab(\Selector0~5_combout ),
	.datac(\Selector0~6_combout ),
	.datad(\Add0~2_combout ),
	.cin(gnd),
	.combout(\Selector30~5_combout ),
	.cout());
// synopsys translate_off
defparam \Selector30~5 .lut_mask = 16'hECA0;
defparam \Selector30~5 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y41_N20
cycloneive_lcell_comb \Selector30~7 (
// Equation(s):
// \Selector30~7_combout  = (\Selector30~6_combout ) # ((\Selector30~4_combout ) # ((\Selector30~3_combout ) # (\Selector30~5_combout )))

	.dataa(\Selector30~6_combout ),
	.datab(\Selector30~4_combout ),
	.datac(\Selector30~3_combout ),
	.datad(\Selector30~5_combout ),
	.cin(gnd),
	.combout(\Selector30~7_combout ),
	.cout());
// synopsys translate_off
defparam \Selector30~7 .lut_mask = 16'hFFFE;
defparam \Selector30~7 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X50_Y40_N24
cycloneive_lcell_comb \Selector31~3 (
// Equation(s):
// \Selector31~3_combout  = (\Add1~0_combout  & ((\Selector0~6_combout ) # ((\Selector0~3_combout  & \portb~58_combout )))) # (!\Add1~0_combout  & (\Selector0~3_combout  & ((\portb~58_combout ))))

	.dataa(\Add1~0_combout ),
	.datab(\Selector0~3_combout ),
	.datac(\Selector0~6_combout ),
	.datad(portb27),
	.cin(gnd),
	.combout(\Selector31~3_combout ),
	.cout());
// synopsys translate_off
defparam \Selector31~3 .lut_mask = 16'hECA0;
defparam \Selector31~3 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X50_Y40_N30
cycloneive_lcell_comb \Selector31~4 (
// Equation(s):
// \Selector31~4_combout  = (\Selector31~3_combout ) # ((\Add0~0_combout  & ((\Selector0~2_combout ) # (\Selector0~5_combout ))))

	.dataa(\Selector0~2_combout ),
	.datab(\Selector0~5_combout ),
	.datac(\Add0~0_combout ),
	.datad(\Selector31~3_combout ),
	.cin(gnd),
	.combout(\Selector31~4_combout ),
	.cout());
// synopsys translate_off
defparam \Selector31~4 .lut_mask = 16'hFFE0;
defparam \Selector31~4 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y37_N22
cycloneive_lcell_comb \ShiftRight0~71 (
// Equation(s):
// \ShiftRight0~71_combout  = (\portb~64_combout ) # ((\portb~62_combout ) # ((\portb~58_combout ) # (\portb~60_combout )))

	.dataa(portb30),
	.datab(portb29),
	.datac(portb27),
	.datad(portb28),
	.cin(gnd),
	.combout(\ShiftRight0~71_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftRight0~71 .lut_mask = 16'hFFFE;
defparam \ShiftRight0~71 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y41_N4
cycloneive_lcell_comb \Selector31~5 (
// Equation(s):
// \Selector31~5_combout  = (\Selector0~3_combout ) # ((\portb~58_combout  & \Selector0~4_combout ))

	.dataa(\Selector0~3_combout ),
	.datab(portb27),
	.datac(gnd),
	.datad(\Selector0~4_combout ),
	.cin(gnd),
	.combout(\Selector31~5_combout ),
	.cout());
// synopsys translate_off
defparam \Selector31~5 .lut_mask = 16'hEEAA;
defparam \Selector31~5 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y41_N30
cycloneive_lcell_comb \Selector31~6 (
// Equation(s):
// \Selector31~6_combout  = (\Selector31~5_combout ) # ((!\ShiftRight0~71_combout  & \Selector30~1_combout ))

	.dataa(gnd),
	.datab(\ShiftRight0~71_combout ),
	.datac(\Selector31~5_combout ),
	.datad(\Selector30~1_combout ),
	.cin(gnd),
	.combout(\Selector31~6_combout ),
	.cout());
// synopsys translate_off
defparam \Selector31~6 .lut_mask = 16'hF3F0;
defparam \Selector31~6 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y41_N8
cycloneive_lcell_comb \Selector31~7 (
// Equation(s):
// \Selector31~7_combout  = (\porta~91_combout  & (((\Selector31~6_combout )))) # (!\porta~91_combout  & (\Selector0~7_combout  & (!\portb~58_combout )))

	.dataa(\Selector0~7_combout ),
	.datab(portb27),
	.datac(\Selector31~6_combout ),
	.datad(porta7),
	.cin(gnd),
	.combout(\Selector31~7_combout ),
	.cout());
// synopsys translate_off
defparam \Selector31~7 .lut_mask = 16'hF022;
defparam \Selector31~7 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X50_Y35_N12
cycloneive_lcell_comb \Selector31~1 (
// Equation(s):
// \Selector31~1_combout  = (!plif_idexaluop_l_2 & (plif_idexaluop_l_3 & plif_idexaluop_l_1))

	.dataa(plif_idexaluop_l_2),
	.datab(plif_idexaluop_l_3),
	.datac(plif_idexaluop_l_1),
	.datad(gnd),
	.cin(gnd),
	.combout(\Selector31~1_combout ),
	.cout());
// synopsys translate_off
defparam \Selector31~1 .lut_mask = 16'h4040;
defparam \Selector31~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X49_Y38_N0
cycloneive_lcell_comb \LessThan0~1 (
// Equation(s):
// \LessThan0~1_cout  = CARRY((\portb~58_combout  & !\porta~91_combout ))

	.dataa(portb27),
	.datab(porta7),
	.datac(gnd),
	.datad(vcc),
	.cin(gnd),
	.combout(),
	.cout(\LessThan0~1_cout ));
// synopsys translate_off
defparam \LessThan0~1 .lut_mask = 16'h0022;
defparam \LessThan0~1 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X49_Y38_N2
cycloneive_lcell_comb \LessThan0~3 (
// Equation(s):
// \LessThan0~3_cout  = CARRY((\portb~60_combout  & (\porta~57_combout  & !\LessThan0~1_cout )) # (!\portb~60_combout  & ((\porta~57_combout ) # (!\LessThan0~1_cout ))))

	.dataa(portb28),
	.datab(porta1),
	.datac(gnd),
	.datad(vcc),
	.cin(\LessThan0~1_cout ),
	.combout(),
	.cout(\LessThan0~3_cout ));
// synopsys translate_off
defparam \LessThan0~3 .lut_mask = 16'h004D;
defparam \LessThan0~3 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X49_Y38_N4
cycloneive_lcell_comb \LessThan0~5 (
// Equation(s):
// \LessThan0~5_cout  = CARRY((\portb~62_combout  & ((!\LessThan0~3_cout ) # (!\porta~55_combout ))) # (!\portb~62_combout  & (!\porta~55_combout  & !\LessThan0~3_cout )))

	.dataa(portb29),
	.datab(porta),
	.datac(gnd),
	.datad(vcc),
	.cin(\LessThan0~3_cout ),
	.combout(),
	.cout(\LessThan0~5_cout ));
// synopsys translate_off
defparam \LessThan0~5 .lut_mask = 16'h002B;
defparam \LessThan0~5 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X49_Y38_N6
cycloneive_lcell_comb \LessThan0~7 (
// Equation(s):
// \LessThan0~7_cout  = CARRY((\porta~61_combout  & ((!\LessThan0~5_cout ) # (!\portb~64_combout ))) # (!\porta~61_combout  & (!\portb~64_combout  & !\LessThan0~5_cout )))

	.dataa(porta3),
	.datab(portb30),
	.datac(gnd),
	.datad(vcc),
	.cin(\LessThan0~5_cout ),
	.combout(),
	.cout(\LessThan0~7_cout ));
// synopsys translate_off
defparam \LessThan0~7 .lut_mask = 16'h002B;
defparam \LessThan0~7 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X49_Y38_N8
cycloneive_lcell_comb \LessThan0~9 (
// Equation(s):
// \LessThan0~9_cout  = CARRY((\portb~66_combout  & ((!\LessThan0~7_cout ) # (!\porta~59_combout ))) # (!\portb~66_combout  & (!\porta~59_combout  & !\LessThan0~7_cout )))

	.dataa(portb31),
	.datab(porta2),
	.datac(gnd),
	.datad(vcc),
	.cin(\LessThan0~7_cout ),
	.combout(),
	.cout(\LessThan0~9_cout ));
// synopsys translate_off
defparam \LessThan0~9 .lut_mask = 16'h002B;
defparam \LessThan0~9 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X49_Y38_N10
cycloneive_lcell_comb \LessThan0~11 (
// Equation(s):
// \LessThan0~11_cout  = CARRY((\porta~95_combout  & ((!\LessThan0~9_cout ) # (!\portb~56_combout ))) # (!\porta~95_combout  & (!\portb~56_combout  & !\LessThan0~9_cout )))

	.dataa(porta11),
	.datab(portb26),
	.datac(gnd),
	.datad(vcc),
	.cin(\LessThan0~9_cout ),
	.combout(),
	.cout(\LessThan0~11_cout ));
// synopsys translate_off
defparam \LessThan0~11 .lut_mask = 16'h002B;
defparam \LessThan0~11 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X49_Y38_N12
cycloneive_lcell_comb \LessThan0~13 (
// Equation(s):
// \LessThan0~13_cout  = CARRY((\porta~94_combout  & (\portb~54_combout  & !\LessThan0~11_cout )) # (!\porta~94_combout  & ((\portb~54_combout ) # (!\LessThan0~11_cout ))))

	.dataa(porta10),
	.datab(portb25),
	.datac(gnd),
	.datad(vcc),
	.cin(\LessThan0~11_cout ),
	.combout(),
	.cout(\LessThan0~13_cout ));
// synopsys translate_off
defparam \LessThan0~13 .lut_mask = 16'h004D;
defparam \LessThan0~13 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X49_Y38_N14
cycloneive_lcell_comb \LessThan0~15 (
// Equation(s):
// \LessThan0~15_cout  = CARRY((\portb~52_combout  & (\porta~93_combout  & !\LessThan0~13_cout )) # (!\portb~52_combout  & ((\porta~93_combout ) # (!\LessThan0~13_cout ))))

	.dataa(portb24),
	.datab(porta9),
	.datac(gnd),
	.datad(vcc),
	.cin(\LessThan0~13_cout ),
	.combout(),
	.cout(\LessThan0~15_cout ));
// synopsys translate_off
defparam \LessThan0~15 .lut_mask = 16'h004D;
defparam \LessThan0~15 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X49_Y38_N16
cycloneive_lcell_comb \LessThan0~17 (
// Equation(s):
// \LessThan0~17_cout  = CARRY((\porta~92_combout  & (\portb~50_combout  & !\LessThan0~15_cout )) # (!\porta~92_combout  & ((\portb~50_combout ) # (!\LessThan0~15_cout ))))

	.dataa(porta8),
	.datab(portb23),
	.datac(gnd),
	.datad(vcc),
	.cin(\LessThan0~15_cout ),
	.combout(),
	.cout(\LessThan0~17_cout ));
// synopsys translate_off
defparam \LessThan0~17 .lut_mask = 16'h004D;
defparam \LessThan0~17 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X49_Y38_N18
cycloneive_lcell_comb \LessThan0~19 (
// Equation(s):
// \LessThan0~19_cout  = CARRY((\portb~48_combout  & (\porta~103_combout  & !\LessThan0~17_cout )) # (!\portb~48_combout  & ((\porta~103_combout ) # (!\LessThan0~17_cout ))))

	.dataa(portb22),
	.datab(porta19),
	.datac(gnd),
	.datad(vcc),
	.cin(\LessThan0~17_cout ),
	.combout(),
	.cout(\LessThan0~19_cout ));
// synopsys translate_off
defparam \LessThan0~19 .lut_mask = 16'h004D;
defparam \LessThan0~19 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X49_Y38_N20
cycloneive_lcell_comb \LessThan0~21 (
// Equation(s):
// \LessThan0~21_cout  = CARRY((\portb~46_combout  & ((!\LessThan0~19_cout ) # (!\porta~102_combout ))) # (!\portb~46_combout  & (!\porta~102_combout  & !\LessThan0~19_cout )))

	.dataa(portb21),
	.datab(porta18),
	.datac(gnd),
	.datad(vcc),
	.cin(\LessThan0~19_cout ),
	.combout(),
	.cout(\LessThan0~21_cout ));
// synopsys translate_off
defparam \LessThan0~21 .lut_mask = 16'h002B;
defparam \LessThan0~21 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X49_Y38_N22
cycloneive_lcell_comb \LessThan0~23 (
// Equation(s):
// \LessThan0~23_cout  = CARRY((\portb~44_combout  & (\porta~101_combout  & !\LessThan0~21_cout )) # (!\portb~44_combout  & ((\porta~101_combout ) # (!\LessThan0~21_cout ))))

	.dataa(portb20),
	.datab(porta17),
	.datac(gnd),
	.datad(vcc),
	.cin(\LessThan0~21_cout ),
	.combout(),
	.cout(\LessThan0~23_cout ));
// synopsys translate_off
defparam \LessThan0~23 .lut_mask = 16'h004D;
defparam \LessThan0~23 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X49_Y38_N24
cycloneive_lcell_comb \LessThan0~25 (
// Equation(s):
// \LessThan0~25_cout  = CARRY((\portb~42_combout  & ((!\LessThan0~23_cout ) # (!\porta~100_combout ))) # (!\portb~42_combout  & (!\porta~100_combout  & !\LessThan0~23_cout )))

	.dataa(portb19),
	.datab(porta16),
	.datac(gnd),
	.datad(vcc),
	.cin(\LessThan0~23_cout ),
	.combout(),
	.cout(\LessThan0~25_cout ));
// synopsys translate_off
defparam \LessThan0~25 .lut_mask = 16'h002B;
defparam \LessThan0~25 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X49_Y38_N26
cycloneive_lcell_comb \LessThan0~27 (
// Equation(s):
// \LessThan0~27_cout  = CARRY((\portb~40_combout  & (\porta~99_combout  & !\LessThan0~25_cout )) # (!\portb~40_combout  & ((\porta~99_combout ) # (!\LessThan0~25_cout ))))

	.dataa(portb18),
	.datab(porta15),
	.datac(gnd),
	.datad(vcc),
	.cin(\LessThan0~25_cout ),
	.combout(),
	.cout(\LessThan0~27_cout ));
// synopsys translate_off
defparam \LessThan0~27 .lut_mask = 16'h004D;
defparam \LessThan0~27 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X49_Y38_N28
cycloneive_lcell_comb \LessThan0~29 (
// Equation(s):
// \LessThan0~29_cout  = CARRY((\portb~38_combout  & ((!\LessThan0~27_cout ) # (!\porta~98_combout ))) # (!\portb~38_combout  & (!\porta~98_combout  & !\LessThan0~27_cout )))

	.dataa(portb17),
	.datab(porta14),
	.datac(gnd),
	.datad(vcc),
	.cin(\LessThan0~27_cout ),
	.combout(),
	.cout(\LessThan0~29_cout ));
// synopsys translate_off
defparam \LessThan0~29 .lut_mask = 16'h002B;
defparam \LessThan0~29 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X49_Y38_N30
cycloneive_lcell_comb \LessThan0~31 (
// Equation(s):
// \LessThan0~31_cout  = CARRY((\porta~97_combout  & ((!\LessThan0~29_cout ) # (!\portb~36_combout ))) # (!\porta~97_combout  & (!\portb~36_combout  & !\LessThan0~29_cout )))

	.dataa(porta13),
	.datab(portb16),
	.datac(gnd),
	.datad(vcc),
	.cin(\LessThan0~29_cout ),
	.combout(),
	.cout(\LessThan0~31_cout ));
// synopsys translate_off
defparam \LessThan0~31 .lut_mask = 16'h002B;
defparam \LessThan0~31 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X49_Y37_N0
cycloneive_lcell_comb \LessThan0~33 (
// Equation(s):
// \LessThan0~33_cout  = CARRY((\porta~96_combout  & (\portb~34_combout  & !\LessThan0~31_cout )) # (!\porta~96_combout  & ((\portb~34_combout ) # (!\LessThan0~31_cout ))))

	.dataa(porta12),
	.datab(portb15),
	.datac(gnd),
	.datad(vcc),
	.cin(\LessThan0~31_cout ),
	.combout(),
	.cout(\LessThan0~33_cout ));
// synopsys translate_off
defparam \LessThan0~33 .lut_mask = 16'h004D;
defparam \LessThan0~33 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X49_Y37_N2
cycloneive_lcell_comb \LessThan0~35 (
// Equation(s):
// \LessThan0~35_cout  = CARRY((\portb~32_combout  & (\porta~118_combout  & !\LessThan0~33_cout )) # (!\portb~32_combout  & ((\porta~118_combout ) # (!\LessThan0~33_cout ))))

	.dataa(portb14),
	.datab(porta34),
	.datac(gnd),
	.datad(vcc),
	.cin(\LessThan0~33_cout ),
	.combout(),
	.cout(\LessThan0~35_cout ));
// synopsys translate_off
defparam \LessThan0~35 .lut_mask = 16'h004D;
defparam \LessThan0~35 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X49_Y37_N4
cycloneive_lcell_comb \LessThan0~37 (
// Equation(s):
// \LessThan0~37_cout  = CARRY((\portb~30_combout  & ((!\LessThan0~35_cout ) # (!\porta~117_combout ))) # (!\portb~30_combout  & (!\porta~117_combout  & !\LessThan0~35_cout )))

	.dataa(portb13),
	.datab(porta33),
	.datac(gnd),
	.datad(vcc),
	.cin(\LessThan0~35_cout ),
	.combout(),
	.cout(\LessThan0~37_cout ));
// synopsys translate_off
defparam \LessThan0~37 .lut_mask = 16'h002B;
defparam \LessThan0~37 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X49_Y37_N6
cycloneive_lcell_comb \LessThan0~39 (
// Equation(s):
// \LessThan0~39_cout  = CARRY((\portb~28_combout  & (\porta~116_combout  & !\LessThan0~37_cout )) # (!\portb~28_combout  & ((\porta~116_combout ) # (!\LessThan0~37_cout ))))

	.dataa(portb12),
	.datab(porta32),
	.datac(gnd),
	.datad(vcc),
	.cin(\LessThan0~37_cout ),
	.combout(),
	.cout(\LessThan0~39_cout ));
// synopsys translate_off
defparam \LessThan0~39 .lut_mask = 16'h004D;
defparam \LessThan0~39 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X49_Y37_N8
cycloneive_lcell_comb \LessThan0~41 (
// Equation(s):
// \LessThan0~41_cout  = CARRY((\porta~115_combout  & (\portb~26_combout  & !\LessThan0~39_cout )) # (!\porta~115_combout  & ((\portb~26_combout ) # (!\LessThan0~39_cout ))))

	.dataa(porta31),
	.datab(portb11),
	.datac(gnd),
	.datad(vcc),
	.cin(\LessThan0~39_cout ),
	.combout(),
	.cout(\LessThan0~41_cout ));
// synopsys translate_off
defparam \LessThan0~41 .lut_mask = 16'h004D;
defparam \LessThan0~41 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X49_Y37_N10
cycloneive_lcell_comb \LessThan0~43 (
// Equation(s):
// \LessThan0~43_cout  = CARRY((\portb~24_combout  & (\porta~114_combout  & !\LessThan0~41_cout )) # (!\portb~24_combout  & ((\porta~114_combout ) # (!\LessThan0~41_cout ))))

	.dataa(portb10),
	.datab(porta30),
	.datac(gnd),
	.datad(vcc),
	.cin(\LessThan0~41_cout ),
	.combout(),
	.cout(\LessThan0~43_cout ));
// synopsys translate_off
defparam \LessThan0~43 .lut_mask = 16'h004D;
defparam \LessThan0~43 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X49_Y37_N12
cycloneive_lcell_comb \LessThan0~45 (
// Equation(s):
// \LessThan0~45_cout  = CARRY((\porta~113_combout  & (\portb~22_combout  & !\LessThan0~43_cout )) # (!\porta~113_combout  & ((\portb~22_combout ) # (!\LessThan0~43_cout ))))

	.dataa(porta29),
	.datab(portb9),
	.datac(gnd),
	.datad(vcc),
	.cin(\LessThan0~43_cout ),
	.combout(),
	.cout(\LessThan0~45_cout ));
// synopsys translate_off
defparam \LessThan0~45 .lut_mask = 16'h004D;
defparam \LessThan0~45 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X49_Y37_N14
cycloneive_lcell_comb \LessThan0~47 (
// Equation(s):
// \LessThan0~47_cout  = CARRY((\portb~20_combout  & (\porta~112_combout  & !\LessThan0~45_cout )) # (!\portb~20_combout  & ((\porta~112_combout ) # (!\LessThan0~45_cout ))))

	.dataa(portb8),
	.datab(porta28),
	.datac(gnd),
	.datad(vcc),
	.cin(\LessThan0~45_cout ),
	.combout(),
	.cout(\LessThan0~47_cout ));
// synopsys translate_off
defparam \LessThan0~47 .lut_mask = 16'h004D;
defparam \LessThan0~47 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X49_Y37_N16
cycloneive_lcell_comb \LessThan0~49 (
// Equation(s):
// \LessThan0~49_cout  = CARRY((\portb~18_combout  & ((!\LessThan0~47_cout ) # (!\porta~111_combout ))) # (!\portb~18_combout  & (!\porta~111_combout  & !\LessThan0~47_cout )))

	.dataa(portb7),
	.datab(porta27),
	.datac(gnd),
	.datad(vcc),
	.cin(\LessThan0~47_cout ),
	.combout(),
	.cout(\LessThan0~49_cout ));
// synopsys translate_off
defparam \LessThan0~49 .lut_mask = 16'h002B;
defparam \LessThan0~49 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X49_Y37_N18
cycloneive_lcell_comb \LessThan0~51 (
// Equation(s):
// \LessThan0~51_cout  = CARRY((\porta~110_combout  & ((!\LessThan0~49_cout ) # (!\portb~16_combout ))) # (!\porta~110_combout  & (!\portb~16_combout  & !\LessThan0~49_cout )))

	.dataa(porta26),
	.datab(portb6),
	.datac(gnd),
	.datad(vcc),
	.cin(\LessThan0~49_cout ),
	.combout(),
	.cout(\LessThan0~51_cout ));
// synopsys translate_off
defparam \LessThan0~51 .lut_mask = 16'h002B;
defparam \LessThan0~51 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X49_Y37_N20
cycloneive_lcell_comb \LessThan0~53 (
// Equation(s):
// \LessThan0~53_cout  = CARRY((\porta~109_combout  & (\portb~14_combout  & !\LessThan0~51_cout )) # (!\porta~109_combout  & ((\portb~14_combout ) # (!\LessThan0~51_cout ))))

	.dataa(porta25),
	.datab(portb5),
	.datac(gnd),
	.datad(vcc),
	.cin(\LessThan0~51_cout ),
	.combout(),
	.cout(\LessThan0~53_cout ));
// synopsys translate_off
defparam \LessThan0~53 .lut_mask = 16'h004D;
defparam \LessThan0~53 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X49_Y37_N22
cycloneive_lcell_comb \LessThan0~55 (
// Equation(s):
// \LessThan0~55_cout  = CARRY((\porta~108_combout  & ((!\LessThan0~53_cout ) # (!\portb~12_combout ))) # (!\porta~108_combout  & (!\portb~12_combout  & !\LessThan0~53_cout )))

	.dataa(porta24),
	.datab(portb4),
	.datac(gnd),
	.datad(vcc),
	.cin(\LessThan0~53_cout ),
	.combout(),
	.cout(\LessThan0~55_cout ));
// synopsys translate_off
defparam \LessThan0~55 .lut_mask = 16'h002B;
defparam \LessThan0~55 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X49_Y37_N24
cycloneive_lcell_comb \LessThan0~57 (
// Equation(s):
// \LessThan0~57_cout  = CARRY((\porta~107_combout  & (\portb~10_combout  & !\LessThan0~55_cout )) # (!\porta~107_combout  & ((\portb~10_combout ) # (!\LessThan0~55_cout ))))

	.dataa(porta23),
	.datab(portb3),
	.datac(gnd),
	.datad(vcc),
	.cin(\LessThan0~55_cout ),
	.combout(),
	.cout(\LessThan0~57_cout ));
// synopsys translate_off
defparam \LessThan0~57 .lut_mask = 16'h004D;
defparam \LessThan0~57 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X49_Y37_N26
cycloneive_lcell_comb \LessThan0~59 (
// Equation(s):
// \LessThan0~59_cout  = CARRY((\porta~105_combout  & ((!\LessThan0~57_cout ) # (!\portb~8_combout ))) # (!\porta~105_combout  & (!\portb~8_combout  & !\LessThan0~57_cout )))

	.dataa(porta21),
	.datab(portb2),
	.datac(gnd),
	.datad(vcc),
	.cin(\LessThan0~57_cout ),
	.combout(),
	.cout(\LessThan0~59_cout ));
// synopsys translate_off
defparam \LessThan0~59 .lut_mask = 16'h002B;
defparam \LessThan0~59 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X49_Y37_N28
cycloneive_lcell_comb \LessThan0~61 (
// Equation(s):
// \LessThan0~61_cout  = CARRY((\porta~106_combout  & (\portb~6_combout  & !\LessThan0~59_cout )) # (!\porta~106_combout  & ((\portb~6_combout ) # (!\LessThan0~59_cout ))))

	.dataa(porta22),
	.datab(portb1),
	.datac(gnd),
	.datad(vcc),
	.cin(\LessThan0~59_cout ),
	.combout(),
	.cout(\LessThan0~61_cout ));
// synopsys translate_off
defparam \LessThan0~61 .lut_mask = 16'h004D;
defparam \LessThan0~61 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X49_Y37_N30
cycloneive_lcell_comb \LessThan0~62 (
// Equation(s):
// \LessThan0~62_combout  = (\portb~4_combout  & (\LessThan0~61_cout  & \porta~104_combout )) # (!\portb~4_combout  & ((\LessThan0~61_cout ) # (\porta~104_combout )))

	.dataa(portb),
	.datab(gnd),
	.datac(gnd),
	.datad(porta20),
	.cin(\LessThan0~61_cout ),
	.combout(\LessThan0~62_combout ),
	.cout());
// synopsys translate_off
defparam \LessThan0~62 .lut_mask = 16'hF550;
defparam \LessThan0~62 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X49_Y40_N0
cycloneive_lcell_comb \LessThan1~1 (
// Equation(s):
// \LessThan1~1_cout  = CARRY((\portb~58_combout  & !\porta~91_combout ))

	.dataa(portb27),
	.datab(porta7),
	.datac(gnd),
	.datad(vcc),
	.cin(gnd),
	.combout(),
	.cout(\LessThan1~1_cout ));
// synopsys translate_off
defparam \LessThan1~1 .lut_mask = 16'h0022;
defparam \LessThan1~1 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X49_Y40_N2
cycloneive_lcell_comb \LessThan1~3 (
// Equation(s):
// \LessThan1~3_cout  = CARRY((\porta~57_combout  & ((!\LessThan1~1_cout ) # (!\portb~60_combout ))) # (!\porta~57_combout  & (!\portb~60_combout  & !\LessThan1~1_cout )))

	.dataa(porta1),
	.datab(portb28),
	.datac(gnd),
	.datad(vcc),
	.cin(\LessThan1~1_cout ),
	.combout(),
	.cout(\LessThan1~3_cout ));
// synopsys translate_off
defparam \LessThan1~3 .lut_mask = 16'h002B;
defparam \LessThan1~3 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X49_Y40_N4
cycloneive_lcell_comb \LessThan1~5 (
// Equation(s):
// \LessThan1~5_cout  = CARRY((\portb~62_combout  & ((!\LessThan1~3_cout ) # (!\porta~55_combout ))) # (!\portb~62_combout  & (!\porta~55_combout  & !\LessThan1~3_cout )))

	.dataa(portb29),
	.datab(porta),
	.datac(gnd),
	.datad(vcc),
	.cin(\LessThan1~3_cout ),
	.combout(),
	.cout(\LessThan1~5_cout ));
// synopsys translate_off
defparam \LessThan1~5 .lut_mask = 16'h002B;
defparam \LessThan1~5 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X49_Y40_N6
cycloneive_lcell_comb \LessThan1~7 (
// Equation(s):
// \LessThan1~7_cout  = CARRY((\porta~61_combout  & ((!\LessThan1~5_cout ) # (!\portb~64_combout ))) # (!\porta~61_combout  & (!\portb~64_combout  & !\LessThan1~5_cout )))

	.dataa(porta3),
	.datab(portb30),
	.datac(gnd),
	.datad(vcc),
	.cin(\LessThan1~5_cout ),
	.combout(),
	.cout(\LessThan1~7_cout ));
// synopsys translate_off
defparam \LessThan1~7 .lut_mask = 16'h002B;
defparam \LessThan1~7 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X49_Y40_N8
cycloneive_lcell_comb \LessThan1~9 (
// Equation(s):
// \LessThan1~9_cout  = CARRY((\portb~66_combout  & ((!\LessThan1~7_cout ) # (!\porta~59_combout ))) # (!\portb~66_combout  & (!\porta~59_combout  & !\LessThan1~7_cout )))

	.dataa(portb31),
	.datab(porta2),
	.datac(gnd),
	.datad(vcc),
	.cin(\LessThan1~7_cout ),
	.combout(),
	.cout(\LessThan1~9_cout ));
// synopsys translate_off
defparam \LessThan1~9 .lut_mask = 16'h002B;
defparam \LessThan1~9 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X49_Y40_N10
cycloneive_lcell_comb \LessThan1~11 (
// Equation(s):
// \LessThan1~11_cout  = CARRY((\porta~95_combout  & ((!\LessThan1~9_cout ) # (!\portb~56_combout ))) # (!\porta~95_combout  & (!\portb~56_combout  & !\LessThan1~9_cout )))

	.dataa(porta11),
	.datab(portb26),
	.datac(gnd),
	.datad(vcc),
	.cin(\LessThan1~9_cout ),
	.combout(),
	.cout(\LessThan1~11_cout ));
// synopsys translate_off
defparam \LessThan1~11 .lut_mask = 16'h002B;
defparam \LessThan1~11 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X49_Y40_N12
cycloneive_lcell_comb \LessThan1~13 (
// Equation(s):
// \LessThan1~13_cout  = CARRY((\porta~94_combout  & (\portb~54_combout  & !\LessThan1~11_cout )) # (!\porta~94_combout  & ((\portb~54_combout ) # (!\LessThan1~11_cout ))))

	.dataa(porta10),
	.datab(portb25),
	.datac(gnd),
	.datad(vcc),
	.cin(\LessThan1~11_cout ),
	.combout(),
	.cout(\LessThan1~13_cout ));
// synopsys translate_off
defparam \LessThan1~13 .lut_mask = 16'h004D;
defparam \LessThan1~13 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X49_Y40_N14
cycloneive_lcell_comb \LessThan1~15 (
// Equation(s):
// \LessThan1~15_cout  = CARRY((\porta~93_combout  & ((!\LessThan1~13_cout ) # (!\portb~52_combout ))) # (!\porta~93_combout  & (!\portb~52_combout  & !\LessThan1~13_cout )))

	.dataa(porta9),
	.datab(portb24),
	.datac(gnd),
	.datad(vcc),
	.cin(\LessThan1~13_cout ),
	.combout(),
	.cout(\LessThan1~15_cout ));
// synopsys translate_off
defparam \LessThan1~15 .lut_mask = 16'h002B;
defparam \LessThan1~15 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X49_Y40_N16
cycloneive_lcell_comb \LessThan1~17 (
// Equation(s):
// \LessThan1~17_cout  = CARRY((\porta~92_combout  & (\portb~50_combout  & !\LessThan1~15_cout )) # (!\porta~92_combout  & ((\portb~50_combout ) # (!\LessThan1~15_cout ))))

	.dataa(porta8),
	.datab(portb23),
	.datac(gnd),
	.datad(vcc),
	.cin(\LessThan1~15_cout ),
	.combout(),
	.cout(\LessThan1~17_cout ));
// synopsys translate_off
defparam \LessThan1~17 .lut_mask = 16'h004D;
defparam \LessThan1~17 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X49_Y40_N18
cycloneive_lcell_comb \LessThan1~19 (
// Equation(s):
// \LessThan1~19_cout  = CARRY((\portb~48_combout  & (\porta~103_combout  & !\LessThan1~17_cout )) # (!\portb~48_combout  & ((\porta~103_combout ) # (!\LessThan1~17_cout ))))

	.dataa(portb22),
	.datab(porta19),
	.datac(gnd),
	.datad(vcc),
	.cin(\LessThan1~17_cout ),
	.combout(),
	.cout(\LessThan1~19_cout ));
// synopsys translate_off
defparam \LessThan1~19 .lut_mask = 16'h004D;
defparam \LessThan1~19 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X49_Y40_N20
cycloneive_lcell_comb \LessThan1~21 (
// Equation(s):
// \LessThan1~21_cout  = CARRY((\portb~46_combout  & ((!\LessThan1~19_cout ) # (!\porta~102_combout ))) # (!\portb~46_combout  & (!\porta~102_combout  & !\LessThan1~19_cout )))

	.dataa(portb21),
	.datab(porta18),
	.datac(gnd),
	.datad(vcc),
	.cin(\LessThan1~19_cout ),
	.combout(),
	.cout(\LessThan1~21_cout ));
// synopsys translate_off
defparam \LessThan1~21 .lut_mask = 16'h002B;
defparam \LessThan1~21 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X49_Y40_N22
cycloneive_lcell_comb \LessThan1~23 (
// Equation(s):
// \LessThan1~23_cout  = CARRY((\portb~44_combout  & (\porta~101_combout  & !\LessThan1~21_cout )) # (!\portb~44_combout  & ((\porta~101_combout ) # (!\LessThan1~21_cout ))))

	.dataa(portb20),
	.datab(porta17),
	.datac(gnd),
	.datad(vcc),
	.cin(\LessThan1~21_cout ),
	.combout(),
	.cout(\LessThan1~23_cout ));
// synopsys translate_off
defparam \LessThan1~23 .lut_mask = 16'h004D;
defparam \LessThan1~23 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X49_Y40_N24
cycloneive_lcell_comb \LessThan1~25 (
// Equation(s):
// \LessThan1~25_cout  = CARRY((\portb~42_combout  & ((!\LessThan1~23_cout ) # (!\porta~100_combout ))) # (!\portb~42_combout  & (!\porta~100_combout  & !\LessThan1~23_cout )))

	.dataa(portb19),
	.datab(porta16),
	.datac(gnd),
	.datad(vcc),
	.cin(\LessThan1~23_cout ),
	.combout(),
	.cout(\LessThan1~25_cout ));
// synopsys translate_off
defparam \LessThan1~25 .lut_mask = 16'h002B;
defparam \LessThan1~25 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X49_Y40_N26
cycloneive_lcell_comb \LessThan1~27 (
// Equation(s):
// \LessThan1~27_cout  = CARRY((\portb~40_combout  & (\porta~99_combout  & !\LessThan1~25_cout )) # (!\portb~40_combout  & ((\porta~99_combout ) # (!\LessThan1~25_cout ))))

	.dataa(portb18),
	.datab(porta15),
	.datac(gnd),
	.datad(vcc),
	.cin(\LessThan1~25_cout ),
	.combout(),
	.cout(\LessThan1~27_cout ));
// synopsys translate_off
defparam \LessThan1~27 .lut_mask = 16'h004D;
defparam \LessThan1~27 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X49_Y40_N28
cycloneive_lcell_comb \LessThan1~29 (
// Equation(s):
// \LessThan1~29_cout  = CARRY((\porta~98_combout  & (\portb~38_combout  & !\LessThan1~27_cout )) # (!\porta~98_combout  & ((\portb~38_combout ) # (!\LessThan1~27_cout ))))

	.dataa(porta14),
	.datab(portb17),
	.datac(gnd),
	.datad(vcc),
	.cin(\LessThan1~27_cout ),
	.combout(),
	.cout(\LessThan1~29_cout ));
// synopsys translate_off
defparam \LessThan1~29 .lut_mask = 16'h004D;
defparam \LessThan1~29 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X49_Y40_N30
cycloneive_lcell_comb \LessThan1~31 (
// Equation(s):
// \LessThan1~31_cout  = CARRY((\porta~97_combout  & ((!\LessThan1~29_cout ) # (!\portb~36_combout ))) # (!\porta~97_combout  & (!\portb~36_combout  & !\LessThan1~29_cout )))

	.dataa(porta13),
	.datab(portb16),
	.datac(gnd),
	.datad(vcc),
	.cin(\LessThan1~29_cout ),
	.combout(),
	.cout(\LessThan1~31_cout ));
// synopsys translate_off
defparam \LessThan1~31 .lut_mask = 16'h002B;
defparam \LessThan1~31 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X49_Y39_N0
cycloneive_lcell_comb \LessThan1~33 (
// Equation(s):
// \LessThan1~33_cout  = CARRY((\porta~96_combout  & (\portb~34_combout  & !\LessThan1~31_cout )) # (!\porta~96_combout  & ((\portb~34_combout ) # (!\LessThan1~31_cout ))))

	.dataa(porta12),
	.datab(portb15),
	.datac(gnd),
	.datad(vcc),
	.cin(\LessThan1~31_cout ),
	.combout(),
	.cout(\LessThan1~33_cout ));
// synopsys translate_off
defparam \LessThan1~33 .lut_mask = 16'h004D;
defparam \LessThan1~33 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X49_Y39_N2
cycloneive_lcell_comb \LessThan1~35 (
// Equation(s):
// \LessThan1~35_cout  = CARRY((\portb~32_combout  & (\porta~118_combout  & !\LessThan1~33_cout )) # (!\portb~32_combout  & ((\porta~118_combout ) # (!\LessThan1~33_cout ))))

	.dataa(portb14),
	.datab(porta34),
	.datac(gnd),
	.datad(vcc),
	.cin(\LessThan1~33_cout ),
	.combout(),
	.cout(\LessThan1~35_cout ));
// synopsys translate_off
defparam \LessThan1~35 .lut_mask = 16'h004D;
defparam \LessThan1~35 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X49_Y39_N4
cycloneive_lcell_comb \LessThan1~37 (
// Equation(s):
// \LessThan1~37_cout  = CARRY((\porta~117_combout  & (\portb~30_combout  & !\LessThan1~35_cout )) # (!\porta~117_combout  & ((\portb~30_combout ) # (!\LessThan1~35_cout ))))

	.dataa(porta33),
	.datab(portb13),
	.datac(gnd),
	.datad(vcc),
	.cin(\LessThan1~35_cout ),
	.combout(),
	.cout(\LessThan1~37_cout ));
// synopsys translate_off
defparam \LessThan1~37 .lut_mask = 16'h004D;
defparam \LessThan1~37 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X49_Y39_N6
cycloneive_lcell_comb \LessThan1~39 (
// Equation(s):
// \LessThan1~39_cout  = CARRY((\portb~28_combout  & (\porta~116_combout  & !\LessThan1~37_cout )) # (!\portb~28_combout  & ((\porta~116_combout ) # (!\LessThan1~37_cout ))))

	.dataa(portb12),
	.datab(porta32),
	.datac(gnd),
	.datad(vcc),
	.cin(\LessThan1~37_cout ),
	.combout(),
	.cout(\LessThan1~39_cout ));
// synopsys translate_off
defparam \LessThan1~39 .lut_mask = 16'h004D;
defparam \LessThan1~39 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X49_Y39_N8
cycloneive_lcell_comb \LessThan1~41 (
// Equation(s):
// \LessThan1~41_cout  = CARRY((\portb~26_combout  & ((!\LessThan1~39_cout ) # (!\porta~115_combout ))) # (!\portb~26_combout  & (!\porta~115_combout  & !\LessThan1~39_cout )))

	.dataa(portb11),
	.datab(porta31),
	.datac(gnd),
	.datad(vcc),
	.cin(\LessThan1~39_cout ),
	.combout(),
	.cout(\LessThan1~41_cout ));
// synopsys translate_off
defparam \LessThan1~41 .lut_mask = 16'h002B;
defparam \LessThan1~41 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X49_Y39_N10
cycloneive_lcell_comb \LessThan1~43 (
// Equation(s):
// \LessThan1~43_cout  = CARRY((\porta~114_combout  & ((!\LessThan1~41_cout ) # (!\portb~24_combout ))) # (!\porta~114_combout  & (!\portb~24_combout  & !\LessThan1~41_cout )))

	.dataa(porta30),
	.datab(portb10),
	.datac(gnd),
	.datad(vcc),
	.cin(\LessThan1~41_cout ),
	.combout(),
	.cout(\LessThan1~43_cout ));
// synopsys translate_off
defparam \LessThan1~43 .lut_mask = 16'h002B;
defparam \LessThan1~43 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X49_Y39_N12
cycloneive_lcell_comb \LessThan1~45 (
// Equation(s):
// \LessThan1~45_cout  = CARRY((\porta~113_combout  & (\portb~22_combout  & !\LessThan1~43_cout )) # (!\porta~113_combout  & ((\portb~22_combout ) # (!\LessThan1~43_cout ))))

	.dataa(porta29),
	.datab(portb9),
	.datac(gnd),
	.datad(vcc),
	.cin(\LessThan1~43_cout ),
	.combout(),
	.cout(\LessThan1~45_cout ));
// synopsys translate_off
defparam \LessThan1~45 .lut_mask = 16'h004D;
defparam \LessThan1~45 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X49_Y39_N14
cycloneive_lcell_comb \LessThan1~47 (
// Equation(s):
// \LessThan1~47_cout  = CARRY((\porta~112_combout  & ((!\LessThan1~45_cout ) # (!\portb~20_combout ))) # (!\porta~112_combout  & (!\portb~20_combout  & !\LessThan1~45_cout )))

	.dataa(porta28),
	.datab(portb8),
	.datac(gnd),
	.datad(vcc),
	.cin(\LessThan1~45_cout ),
	.combout(),
	.cout(\LessThan1~47_cout ));
// synopsys translate_off
defparam \LessThan1~47 .lut_mask = 16'h002B;
defparam \LessThan1~47 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X49_Y39_N16
cycloneive_lcell_comb \LessThan1~49 (
// Equation(s):
// \LessThan1~49_cout  = CARRY((\portb~18_combout  & ((!\LessThan1~47_cout ) # (!\porta~111_combout ))) # (!\portb~18_combout  & (!\porta~111_combout  & !\LessThan1~47_cout )))

	.dataa(portb7),
	.datab(porta27),
	.datac(gnd),
	.datad(vcc),
	.cin(\LessThan1~47_cout ),
	.combout(),
	.cout(\LessThan1~49_cout ));
// synopsys translate_off
defparam \LessThan1~49 .lut_mask = 16'h002B;
defparam \LessThan1~49 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X49_Y39_N18
cycloneive_lcell_comb \LessThan1~51 (
// Equation(s):
// \LessThan1~51_cout  = CARRY((\porta~110_combout  & ((!\LessThan1~49_cout ) # (!\portb~16_combout ))) # (!\porta~110_combout  & (!\portb~16_combout  & !\LessThan1~49_cout )))

	.dataa(porta26),
	.datab(portb6),
	.datac(gnd),
	.datad(vcc),
	.cin(\LessThan1~49_cout ),
	.combout(),
	.cout(\LessThan1~51_cout ));
// synopsys translate_off
defparam \LessThan1~51 .lut_mask = 16'h002B;
defparam \LessThan1~51 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X49_Y39_N20
cycloneive_lcell_comb \LessThan1~53 (
// Equation(s):
// \LessThan1~53_cout  = CARRY((\porta~109_combout  & (\portb~14_combout  & !\LessThan1~51_cout )) # (!\porta~109_combout  & ((\portb~14_combout ) # (!\LessThan1~51_cout ))))

	.dataa(porta25),
	.datab(portb5),
	.datac(gnd),
	.datad(vcc),
	.cin(\LessThan1~51_cout ),
	.combout(),
	.cout(\LessThan1~53_cout ));
// synopsys translate_off
defparam \LessThan1~53 .lut_mask = 16'h004D;
defparam \LessThan1~53 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X49_Y39_N22
cycloneive_lcell_comb \LessThan1~55 (
// Equation(s):
// \LessThan1~55_cout  = CARRY((\portb~12_combout  & (\porta~108_combout  & !\LessThan1~53_cout )) # (!\portb~12_combout  & ((\porta~108_combout ) # (!\LessThan1~53_cout ))))

	.dataa(portb4),
	.datab(porta24),
	.datac(gnd),
	.datad(vcc),
	.cin(\LessThan1~53_cout ),
	.combout(),
	.cout(\LessThan1~55_cout ));
// synopsys translate_off
defparam \LessThan1~55 .lut_mask = 16'h004D;
defparam \LessThan1~55 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X49_Y39_N24
cycloneive_lcell_comb \LessThan1~57 (
// Equation(s):
// \LessThan1~57_cout  = CARRY((\portb~10_combout  & ((!\LessThan1~55_cout ) # (!\porta~107_combout ))) # (!\portb~10_combout  & (!\porta~107_combout  & !\LessThan1~55_cout )))

	.dataa(portb3),
	.datab(porta23),
	.datac(gnd),
	.datad(vcc),
	.cin(\LessThan1~55_cout ),
	.combout(),
	.cout(\LessThan1~57_cout ));
// synopsys translate_off
defparam \LessThan1~57 .lut_mask = 16'h002B;
defparam \LessThan1~57 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X49_Y39_N26
cycloneive_lcell_comb \LessThan1~59 (
// Equation(s):
// \LessThan1~59_cout  = CARRY((\porta~105_combout  & ((!\LessThan1~57_cout ) # (!\portb~8_combout ))) # (!\porta~105_combout  & (!\portb~8_combout  & !\LessThan1~57_cout )))

	.dataa(porta21),
	.datab(portb2),
	.datac(gnd),
	.datad(vcc),
	.cin(\LessThan1~57_cout ),
	.combout(),
	.cout(\LessThan1~59_cout ));
// synopsys translate_off
defparam \LessThan1~59 .lut_mask = 16'h002B;
defparam \LessThan1~59 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X49_Y39_N28
cycloneive_lcell_comb \LessThan1~61 (
// Equation(s):
// \LessThan1~61_cout  = CARRY((\porta~106_combout  & (\portb~6_combout  & !\LessThan1~59_cout )) # (!\porta~106_combout  & ((\portb~6_combout ) # (!\LessThan1~59_cout ))))

	.dataa(porta22),
	.datab(portb1),
	.datac(gnd),
	.datad(vcc),
	.cin(\LessThan1~59_cout ),
	.combout(),
	.cout(\LessThan1~61_cout ));
// synopsys translate_off
defparam \LessThan1~61 .lut_mask = 16'h004D;
defparam \LessThan1~61 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X49_Y39_N30
cycloneive_lcell_comb \LessThan1~62 (
// Equation(s):
// \LessThan1~62_combout  = (\portb~4_combout  & ((\LessThan1~61_cout ) # (!\porta~104_combout ))) # (!\portb~4_combout  & (\LessThan1~61_cout  & !\porta~104_combout ))

	.dataa(gnd),
	.datab(portb),
	.datac(gnd),
	.datad(porta20),
	.cin(\LessThan1~61_cout ),
	.combout(\LessThan1~62_combout ),
	.cout());
// synopsys translate_off
defparam \LessThan1~62 .lut_mask = 16'hC0FC;
defparam \LessThan1~62 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X50_Y39_N30
cycloneive_lcell_comb \Selector31~2 (
// Equation(s):
// \Selector31~2_combout  = (\Selector31~1_combout  & ((plif_idexaluop_l_0 & ((\LessThan1~62_combout ))) # (!plif_idexaluop_l_0 & (\LessThan0~62_combout ))))

	.dataa(plif_idexaluop_l_0),
	.datab(\Selector31~1_combout ),
	.datac(\LessThan0~62_combout ),
	.datad(\LessThan1~62_combout ),
	.cin(gnd),
	.combout(\Selector31~2_combout ),
	.cout());
// synopsys translate_off
defparam \Selector31~2 .lut_mask = 16'hC840;
defparam \Selector31~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y36_N8
cycloneive_lcell_comb \ShiftRight0~60 (
// Equation(s):
// \ShiftRight0~60_combout  = (\portb~58_combout  & (\porta~108_combout )) # (!\portb~58_combout  & ((\porta~109_combout )))

	.dataa(porta24),
	.datab(porta25),
	.datac(gnd),
	.datad(portb27),
	.cin(gnd),
	.combout(\ShiftRight0~60_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftRight0~60 .lut_mask = 16'hAACC;
defparam \ShiftRight0~60 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y36_N22
cycloneive_lcell_comb \ShiftRight0~61 (
// Equation(s):
// \ShiftRight0~61_combout  = (\portb~58_combout  & (\porta~110_combout )) # (!\portb~58_combout  & ((\porta~111_combout )))

	.dataa(gnd),
	.datab(portb27),
	.datac(porta26),
	.datad(porta27),
	.cin(gnd),
	.combout(\ShiftRight0~61_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftRight0~61 .lut_mask = 16'hF3C0;
defparam \ShiftRight0~61 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y36_N0
cycloneive_lcell_comb \ShiftRight0~62 (
// Equation(s):
// \ShiftRight0~62_combout  = (\portb~60_combout  & (\ShiftRight0~60_combout )) # (!\portb~60_combout  & ((\ShiftRight0~61_combout )))

	.dataa(portb28),
	.datab(\ShiftRight0~60_combout ),
	.datac(\ShiftRight0~61_combout ),
	.datad(gnd),
	.cin(gnd),
	.combout(\ShiftRight0~62_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftRight0~62 .lut_mask = 16'hD8D8;
defparam \ShiftRight0~62 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y39_N2
cycloneive_lcell_comb \ShiftRight0~58 (
// Equation(s):
// \ShiftRight0~58_combout  = (\portb~58_combout  & ((\porta~105_combout ))) # (!\portb~58_combout  & (\porta~107_combout ))

	.dataa(porta23),
	.datab(portb27),
	.datac(gnd),
	.datad(porta21),
	.cin(gnd),
	.combout(\ShiftRight0~58_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftRight0~58 .lut_mask = 16'hEE22;
defparam \ShiftRight0~58 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y39_N20
cycloneive_lcell_comb \ShiftRight0~57 (
// Equation(s):
// \ShiftRight0~57_combout  = (\portb~58_combout  & (\porta~104_combout )) # (!\portb~58_combout  & ((\porta~106_combout )))

	.dataa(porta20),
	.datab(portb27),
	.datac(gnd),
	.datad(porta22),
	.cin(gnd),
	.combout(\ShiftRight0~57_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftRight0~57 .lut_mask = 16'hBB88;
defparam \ShiftRight0~57 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y39_N0
cycloneive_lcell_comb \ShiftRight0~59 (
// Equation(s):
// \ShiftRight0~59_combout  = (\portb~60_combout  & ((\ShiftRight0~57_combout ))) # (!\portb~60_combout  & (\ShiftRight0~58_combout ))

	.dataa(gnd),
	.datab(portb28),
	.datac(\ShiftRight0~58_combout ),
	.datad(\ShiftRight0~57_combout ),
	.cin(gnd),
	.combout(\ShiftRight0~59_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftRight0~59 .lut_mask = 16'hFC30;
defparam \ShiftRight0~59 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y40_N22
cycloneive_lcell_comb \ShiftRight0~63 (
// Equation(s):
// \ShiftRight0~63_combout  = (\portb~62_combout  & ((\ShiftRight0~59_combout ))) # (!\portb~62_combout  & (\ShiftRight0~62_combout ))

	.dataa(portb29),
	.datab(gnd),
	.datac(\ShiftRight0~62_combout ),
	.datad(\ShiftRight0~59_combout ),
	.cin(gnd),
	.combout(\ShiftRight0~63_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftRight0~63 .lut_mask = 16'hFA50;
defparam \ShiftRight0~63 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y36_N28
cycloneive_lcell_comb \ShiftRight0~68 (
// Equation(s):
// \ShiftRight0~68_combout  = (\portb~58_combout  & ((\porta~118_combout ))) # (!\portb~58_combout  & (\porta~96_combout ))

	.dataa(gnd),
	.datab(porta12),
	.datac(porta34),
	.datad(portb27),
	.cin(gnd),
	.combout(\ShiftRight0~68_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftRight0~68 .lut_mask = 16'hF0CC;
defparam \ShiftRight0~68 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y36_N20
cycloneive_lcell_comb \ShiftRight0~67 (
// Equation(s):
// \ShiftRight0~67_combout  = (\portb~58_combout  & (\porta~116_combout )) # (!\portb~58_combout  & ((\porta~117_combout )))

	.dataa(porta32),
	.datab(gnd),
	.datac(porta33),
	.datad(portb27),
	.cin(gnd),
	.combout(\ShiftRight0~67_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftRight0~67 .lut_mask = 16'hAAF0;
defparam \ShiftRight0~67 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X52_Y35_N14
cycloneive_lcell_comb \ShiftRight0~69 (
// Equation(s):
// \ShiftRight0~69_combout  = (\portb~60_combout  & ((\ShiftRight0~67_combout ))) # (!\portb~60_combout  & (\ShiftRight0~68_combout ))

	.dataa(portb28),
	.datab(gnd),
	.datac(\ShiftRight0~68_combout ),
	.datad(\ShiftRight0~67_combout ),
	.cin(gnd),
	.combout(\ShiftRight0~69_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftRight0~69 .lut_mask = 16'hFA50;
defparam \ShiftRight0~69 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y36_N2
cycloneive_lcell_comb \ShiftRight0~65 (
// Equation(s):
// \ShiftRight0~65_combout  = (\portb~58_combout  & (\porta~114_combout )) # (!\portb~58_combout  & ((\porta~115_combout )))

	.dataa(gnd),
	.datab(portb27),
	.datac(porta30),
	.datad(porta31),
	.cin(gnd),
	.combout(\ShiftRight0~65_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftRight0~65 .lut_mask = 16'hF3C0;
defparam \ShiftRight0~65 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y39_N24
cycloneive_lcell_comb \ShiftRight0~64 (
// Equation(s):
// \ShiftRight0~64_combout  = (\portb~58_combout  & ((\porta~112_combout ))) # (!\portb~58_combout  & (\porta~113_combout ))

	.dataa(gnd),
	.datab(porta29),
	.datac(portb27),
	.datad(porta28),
	.cin(gnd),
	.combout(\ShiftRight0~64_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftRight0~64 .lut_mask = 16'hFC0C;
defparam \ShiftRight0~64 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y36_N26
cycloneive_lcell_comb \ShiftRight0~66 (
// Equation(s):
// \ShiftRight0~66_combout  = (\portb~60_combout  & ((\ShiftRight0~64_combout ))) # (!\portb~60_combout  & (\ShiftRight0~65_combout ))

	.dataa(gnd),
	.datab(\ShiftRight0~65_combout ),
	.datac(portb28),
	.datad(\ShiftRight0~64_combout ),
	.cin(gnd),
	.combout(\ShiftRight0~66_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftRight0~66 .lut_mask = 16'hFC0C;
defparam \ShiftRight0~66 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X52_Y35_N16
cycloneive_lcell_comb \Selector23~0 (
// Equation(s):
// \Selector23~0_combout  = (\portb~62_combout  & ((\ShiftRight0~66_combout ))) # (!\portb~62_combout  & (\ShiftRight0~69_combout ))

	.dataa(gnd),
	.datab(portb29),
	.datac(\ShiftRight0~69_combout ),
	.datad(\ShiftRight0~66_combout ),
	.cin(gnd),
	.combout(\Selector23~0_combout ),
	.cout());
// synopsys translate_off
defparam \Selector23~0 .lut_mask = 16'hFC30;
defparam \Selector23~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X52_Y35_N26
cycloneive_lcell_comb \ShiftRight0~70 (
// Equation(s):
// \ShiftRight0~70_combout  = (\portb~64_combout  & (\ShiftRight0~63_combout )) # (!\portb~64_combout  & ((\Selector23~0_combout )))

	.dataa(portb30),
	.datab(gnd),
	.datac(\ShiftRight0~63_combout ),
	.datad(\Selector23~0_combout ),
	.cin(gnd),
	.combout(\ShiftRight0~70_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftRight0~70 .lut_mask = 16'hF5A0;
defparam \ShiftRight0~70 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y36_N24
cycloneive_lcell_comb \ShiftRight0~50 (
// Equation(s):
// \ShiftRight0~50_combout  = (\portb~58_combout  & (\porta~99_combout )) # (!\portb~58_combout  & ((\porta~100_combout )))

	.dataa(portb27),
	.datab(gnd),
	.datac(porta15),
	.datad(porta16),
	.cin(gnd),
	.combout(\ShiftRight0~50_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftRight0~50 .lut_mask = 16'hF5A0;
defparam \ShiftRight0~50 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y36_N6
cycloneive_lcell_comb \ShiftRight0~49 (
// Equation(s):
// \ShiftRight0~49_combout  = (\portb~58_combout  & (\porta~97_combout )) # (!\portb~58_combout  & ((\porta~98_combout )))

	.dataa(porta13),
	.datab(gnd),
	.datac(porta14),
	.datad(portb27),
	.cin(gnd),
	.combout(\ShiftRight0~49_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftRight0~49 .lut_mask = 16'hAAF0;
defparam \ShiftRight0~49 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y36_N14
cycloneive_lcell_comb \ShiftRight0~51 (
// Equation(s):
// \ShiftRight0~51_combout  = (\portb~60_combout  & ((\ShiftRight0~49_combout ))) # (!\portb~60_combout  & (\ShiftRight0~50_combout ))

	.dataa(gnd),
	.datab(\ShiftRight0~50_combout ),
	.datac(portb28),
	.datad(\ShiftRight0~49_combout ),
	.cin(gnd),
	.combout(\ShiftRight0~51_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftRight0~51 .lut_mask = 16'hFC0C;
defparam \ShiftRight0~51 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y36_N0
cycloneive_lcell_comb \ShiftRight0~52 (
// Equation(s):
// \ShiftRight0~52_combout  = (\portb~58_combout  & ((\porta~101_combout ))) # (!\portb~58_combout  & (\porta~102_combout ))

	.dataa(porta18),
	.datab(gnd),
	.datac(portb27),
	.datad(porta17),
	.cin(gnd),
	.combout(\ShiftRight0~52_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftRight0~52 .lut_mask = 16'hFA0A;
defparam \ShiftRight0~52 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X52_Y41_N16
cycloneive_lcell_comb \ShiftRight0~53 (
// Equation(s):
// \ShiftRight0~53_combout  = (\portb~58_combout  & (\porta~103_combout )) # (!\portb~58_combout  & ((\porta~92_combout )))

	.dataa(portb27),
	.datab(gnd),
	.datac(porta19),
	.datad(porta8),
	.cin(gnd),
	.combout(\ShiftRight0~53_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftRight0~53 .lut_mask = 16'hF5A0;
defparam \ShiftRight0~53 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y36_N10
cycloneive_lcell_comb \ShiftRight0~54 (
// Equation(s):
// \ShiftRight0~54_combout  = (\portb~60_combout  & (\ShiftRight0~52_combout )) # (!\portb~60_combout  & ((\ShiftRight0~53_combout )))

	.dataa(gnd),
	.datab(\ShiftRight0~52_combout ),
	.datac(portb28),
	.datad(\ShiftRight0~53_combout ),
	.cin(gnd),
	.combout(\ShiftRight0~54_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftRight0~54 .lut_mask = 16'hCFC0;
defparam \ShiftRight0~54 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y36_N12
cycloneive_lcell_comb \ShiftRight0~55 (
// Equation(s):
// \ShiftRight0~55_combout  = (\portb~62_combout  & (\ShiftRight0~51_combout )) # (!\portb~62_combout  & ((\ShiftRight0~54_combout )))

	.dataa(portb29),
	.datab(gnd),
	.datac(\ShiftRight0~51_combout ),
	.datad(\ShiftRight0~54_combout ),
	.cin(gnd),
	.combout(\ShiftRight0~55_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftRight0~55 .lut_mask = 16'hF5A0;
defparam \ShiftRight0~55 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X52_Y35_N20
cycloneive_lcell_comb \ShiftRight0~56 (
// Equation(s):
// \ShiftRight0~56_combout  = (!\portb~66_combout  & ((\ShiftRight0~48_combout ) # ((\portb~64_combout  & \ShiftRight0~55_combout ))))

	.dataa(\ShiftRight0~48_combout ),
	.datab(portb30),
	.datac(portb31),
	.datad(\ShiftRight0~55_combout ),
	.cin(gnd),
	.combout(\ShiftRight0~56_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftRight0~56 .lut_mask = 16'h0E0A;
defparam \ShiftRight0~56 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X52_Y35_N28
cycloneive_lcell_comb \Selector31~0 (
// Equation(s):
// \Selector31~0_combout  = (\Selector24~0_combout  & ((\ShiftRight0~56_combout ) # ((\portb~66_combout  & \ShiftRight0~70_combout ))))

	.dataa(portb31),
	.datab(\Selector24~0_combout ),
	.datac(\ShiftRight0~70_combout ),
	.datad(\ShiftRight0~56_combout ),
	.cin(gnd),
	.combout(\Selector31~0_combout ),
	.cout());
// synopsys translate_off
defparam \Selector31~0 .lut_mask = 16'hCC80;
defparam \Selector31~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y38_N14
cycloneive_lcell_comb \ShiftRight0~5 (
// Equation(s):
// \ShiftRight0~5_combout  = (\portb~14_combout ) # ((\portb~12_combout ) # ((\portb~16_combout ) # (\portb~18_combout )))

	.dataa(portb5),
	.datab(portb4),
	.datac(portb6),
	.datad(portb7),
	.cin(gnd),
	.combout(\ShiftRight0~5_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftRight0~5 .lut_mask = 16'hFFFE;
defparam \ShiftRight0~5 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y38_N4
cycloneive_lcell_comb \ShiftRight0~4 (
// Equation(s):
// \ShiftRight0~4_combout  = (\portb~10_combout ) # ((\portb~6_combout ) # ((\portb~8_combout ) # (\portb~4_combout )))

	.dataa(portb3),
	.datab(portb1),
	.datac(portb2),
	.datad(portb),
	.cin(gnd),
	.combout(\ShiftRight0~4_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftRight0~4 .lut_mask = 16'hFFFE;
defparam \ShiftRight0~4 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y38_N20
cycloneive_lcell_comb \ShiftRight0~6 (
// Equation(s):
// \ShiftRight0~6_combout  = (\portb~26_combout ) # ((\portb~20_combout ) # ((\portb~24_combout ) # (\portb~22_combout )))

	.dataa(portb11),
	.datab(portb8),
	.datac(portb10),
	.datad(portb9),
	.cin(gnd),
	.combout(\ShiftRight0~6_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftRight0~6 .lut_mask = 16'hFFFE;
defparam \ShiftRight0~6 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y38_N16
cycloneive_lcell_comb \ShiftRight0~8 (
// Equation(s):
// \ShiftRight0~8_combout  = (\ShiftRight0~7_combout ) # ((\ShiftRight0~5_combout ) # ((\ShiftRight0~4_combout ) # (\ShiftRight0~6_combout )))

	.dataa(\ShiftRight0~7_combout ),
	.datab(\ShiftRight0~5_combout ),
	.datac(\ShiftRight0~4_combout ),
	.datad(\ShiftRight0~6_combout ),
	.cin(gnd),
	.combout(\ShiftRight0~8_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftRight0~8 .lut_mask = 16'hFFFE;
defparam \ShiftRight0~8 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y38_N26
cycloneive_lcell_comb \Selector0~15 (
// Equation(s):
// \Selector0~15_combout  = (!plif_idexaluop_l_1 & (!plif_idexaluop_l_2 & (!\ShiftRight0~41_combout  & !\ShiftRight0~8_combout )))

	.dataa(plif_idexaluop_l_1),
	.datab(plif_idexaluop_l_2),
	.datac(\ShiftRight0~41_combout ),
	.datad(\ShiftRight0~8_combout ),
	.cin(gnd),
	.combout(\Selector0~15_combout ),
	.cout());
// synopsys translate_off
defparam \Selector0~15 .lut_mask = 16'h0001;
defparam \Selector0~15 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y40_N20
cycloneive_lcell_comb \Selector23~1 (
// Equation(s):
// \Selector23~1_combout  = (!plif_idexaluop_l_3 & (\portb~66_combout  & (\Selector0~15_combout  & plif_idexaluop_l_0)))

	.dataa(plif_idexaluop_l_3),
	.datab(portb31),
	.datac(\Selector0~15_combout ),
	.datad(plif_idexaluop_l_0),
	.cin(gnd),
	.combout(\Selector23~1_combout ),
	.cout());
// synopsys translate_off
defparam \Selector23~1 .lut_mask = 16'h4000;
defparam \Selector23~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y38_N24
cycloneive_lcell_comb \ShiftRight0~72 (
// Equation(s):
// \ShiftRight0~72_combout  = (\ShiftRight0~10_combout ) # ((\ShiftRight0~9_combout ) # ((\ShiftRight0~40_combout ) # (\ShiftRight0~8_combout )))

	.dataa(\ShiftRight0~10_combout ),
	.datab(\ShiftRight0~9_combout ),
	.datac(\ShiftRight0~40_combout ),
	.datad(\ShiftRight0~8_combout ),
	.cin(gnd),
	.combout(\ShiftRight0~72_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftRight0~72 .lut_mask = 16'hFFFE;
defparam \ShiftRight0~72 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X52_Y40_N6
cycloneive_lcell_comb \Selector3~0 (
// Equation(s):
// \Selector3~0_combout  = (plif_idexaluop_l_3) # ((plif_idexaluop_l_2) # ((\portb~66_combout  & !\ShiftRight0~72_combout )))

	.dataa(portb31),
	.datab(plif_idexaluop_l_3),
	.datac(plif_idexaluop_l_2),
	.datad(\ShiftRight0~72_combout ),
	.cin(gnd),
	.combout(\Selector3~0_combout ),
	.cout());
// synopsys translate_off
defparam \Selector3~0 .lut_mask = 16'hFCFE;
defparam \Selector3~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X52_Y40_N24
cycloneive_lcell_comb \Selector28~1 (
// Equation(s):
// \Selector28~1_combout  = (!\ShiftRight0~72_combout  & (plif_idexaluop_l_0 & (!plif_idexaluop_l_1 & !\Selector3~0_combout )))

	.dataa(\ShiftRight0~72_combout ),
	.datab(plif_idexaluop_l_0),
	.datac(plif_idexaluop_l_1),
	.datad(\Selector3~0_combout ),
	.cin(gnd),
	.combout(\Selector28~1_combout ),
	.cout());
// synopsys translate_off
defparam \Selector28~1 .lut_mask = 16'h0004;
defparam \Selector28~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X50_Y37_N28
cycloneive_lcell_comb \Selector3~1 (
// Equation(s):
// \Selector3~1_combout  = (\portb~64_combout ) # ((\portb~60_combout  & !\portb~62_combout ))

	.dataa(portb28),
	.datab(gnd),
	.datac(portb30),
	.datad(portb29),
	.cin(gnd),
	.combout(\Selector3~1_combout ),
	.cout());
// synopsys translate_off
defparam \Selector3~1 .lut_mask = 16'hF0FA;
defparam \Selector3~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y41_N16
cycloneive_lcell_comb \ShiftRight0~13 (
// Equation(s):
// \ShiftRight0~13_combout  = (\portb~58_combout  & (\porta~59_combout )) # (!\portb~58_combout  & ((\porta~61_combout )))

	.dataa(portb27),
	.datab(porta2),
	.datac(gnd),
	.datad(porta3),
	.cin(gnd),
	.combout(\ShiftRight0~13_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftRight0~13 .lut_mask = 16'hDD88;
defparam \ShiftRight0~13 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X52_Y41_N8
cycloneive_lcell_comb \ShiftRight0~15 (
// Equation(s):
// \ShiftRight0~15_combout  = (\portb~58_combout  & ((\porta~92_combout ))) # (!\portb~58_combout  & (\porta~93_combout ))

	.dataa(porta9),
	.datab(porta8),
	.datac(gnd),
	.datad(portb27),
	.cin(gnd),
	.combout(\ShiftRight0~15_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftRight0~15 .lut_mask = 16'hCCAA;
defparam \ShiftRight0~15 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X52_Y41_N6
cycloneive_lcell_comb \ShiftRight0~23 (
// Equation(s):
// \ShiftRight0~23_combout  = (\portb~58_combout  & ((\porta~102_combout ))) # (!\portb~58_combout  & (\porta~103_combout ))

	.dataa(gnd),
	.datab(porta19),
	.datac(porta18),
	.datad(portb27),
	.cin(gnd),
	.combout(\ShiftRight0~23_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftRight0~23 .lut_mask = 16'hF0CC;
defparam \ShiftRight0~23 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X52_Y41_N14
cycloneive_lcell_comb \ShiftRight0~73 (
// Equation(s):
// \ShiftRight0~73_combout  = (\portb~60_combout  & ((\ShiftRight0~23_combout ))) # (!\portb~60_combout  & (\ShiftRight0~15_combout ))

	.dataa(gnd),
	.datab(portb28),
	.datac(\ShiftRight0~15_combout ),
	.datad(\ShiftRight0~23_combout ),
	.cin(gnd),
	.combout(\ShiftRight0~73_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftRight0~73 .lut_mask = 16'hFC30;
defparam \ShiftRight0~73 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X52_Y40_N22
cycloneive_lcell_comb \Selector28~2 (
// Equation(s):
// \Selector28~2_combout  = (\ShiftRight0~74_combout  & (!\Selector3~1_combout  & (\ShiftRight0~13_combout ))) # (!\ShiftRight0~74_combout  & ((\Selector3~1_combout ) # ((\ShiftRight0~73_combout ))))

	.dataa(\ShiftRight0~74_combout ),
	.datab(\Selector3~1_combout ),
	.datac(\ShiftRight0~13_combout ),
	.datad(\ShiftRight0~73_combout ),
	.cin(gnd),
	.combout(\Selector28~2_combout ),
	.cout());
// synopsys translate_off
defparam \Selector28~2 .lut_mask = 16'h7564;
defparam \Selector28~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y40_N20
cycloneive_lcell_comb \ShiftRight0~19 (
// Equation(s):
// \ShiftRight0~19_combout  = (\portb~58_combout  & ((\porta~96_combout ))) # (!\portb~58_combout  & (\porta~97_combout ))

	.dataa(gnd),
	.datab(portb27),
	.datac(porta13),
	.datad(porta12),
	.cin(gnd),
	.combout(\ShiftRight0~19_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftRight0~19 .lut_mask = 16'hFC30;
defparam \ShiftRight0~19 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y40_N28
cycloneive_lcell_comb \ShiftRight0~75 (
// Equation(s):
// \ShiftRight0~75_combout  = (\portb~60_combout  & (\ShiftRight0~37_combout )) # (!\portb~60_combout  & ((\ShiftRight0~19_combout )))

	.dataa(\ShiftRight0~37_combout ),
	.datab(gnd),
	.datac(portb28),
	.datad(\ShiftRight0~19_combout ),
	.cin(gnd),
	.combout(\ShiftRight0~75_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftRight0~75 .lut_mask = 16'hAFA0;
defparam \ShiftRight0~75 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y42_N14
cycloneive_lcell_comb \ShiftRight0~20 (
// Equation(s):
// \ShiftRight0~20_combout  = (\portb~58_combout  & ((\porta~98_combout ))) # (!\portb~58_combout  & (\porta~99_combout ))

	.dataa(porta15),
	.datab(gnd),
	.datac(portb27),
	.datad(porta14),
	.cin(gnd),
	.combout(\ShiftRight0~20_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftRight0~20 .lut_mask = 16'hFA0A;
defparam \ShiftRight0~20 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y42_N10
cycloneive_lcell_comb \ShiftRight0~76 (
// Equation(s):
// \ShiftRight0~76_combout  = (\portb~60_combout  & (\ShiftRight0~20_combout )) # (!\portb~60_combout  & ((\ShiftRight0~22_combout )))

	.dataa(gnd),
	.datab(portb28),
	.datac(\ShiftRight0~20_combout ),
	.datad(\ShiftRight0~22_combout ),
	.cin(gnd),
	.combout(\ShiftRight0~76_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftRight0~76 .lut_mask = 16'hF3C0;
defparam \ShiftRight0~76 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y42_N20
cycloneive_lcell_comb \ShiftRight0~77 (
// Equation(s):
// \ShiftRight0~77_combout  = (\portb~62_combout  & (\ShiftRight0~75_combout )) # (!\portb~62_combout  & ((\ShiftRight0~76_combout )))

	.dataa(gnd),
	.datab(portb29),
	.datac(\ShiftRight0~75_combout ),
	.datad(\ShiftRight0~76_combout ),
	.cin(gnd),
	.combout(\ShiftRight0~77_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftRight0~77 .lut_mask = 16'hF3C0;
defparam \ShiftRight0~77 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X52_Y40_N4
cycloneive_lcell_comb \Selector28~3 (
// Equation(s):
// \Selector28~3_combout  = (\Selector3~1_combout  & ((\Selector28~2_combout  & ((\ShiftRight0~77_combout ))) # (!\Selector28~2_combout  & (\ShiftRight0~16_combout )))) # (!\Selector3~1_combout  & (((\Selector28~2_combout ))))

	.dataa(\ShiftRight0~16_combout ),
	.datab(\Selector3~1_combout ),
	.datac(\Selector28~2_combout ),
	.datad(\ShiftRight0~77_combout ),
	.cin(gnd),
	.combout(\Selector28~3_combout ),
	.cout());
// synopsys translate_off
defparam \Selector28~3 .lut_mask = 16'hF838;
defparam \Selector28~3 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X50_Y35_N24
cycloneive_lcell_comb \Selector0~9 (
// Equation(s):
// \Selector0~9_combout  = (!plif_idexaluop_l_2 & (!plif_idexaluop_l_3 & (plif_idexaluop_l_1 & !plif_idexaluop_l_0)))

	.dataa(plif_idexaluop_l_2),
	.datab(plif_idexaluop_l_3),
	.datac(plif_idexaluop_l_1),
	.datad(plif_idexaluop_l_0),
	.cin(gnd),
	.combout(\Selector0~9_combout ),
	.cout());
// synopsys translate_off
defparam \Selector0~9 .lut_mask = 16'h0010;
defparam \Selector0~9 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y40_N4
cycloneive_lcell_comb \Add1~4 (
// Equation(s):
// \Add1~4_combout  = ((\porta~55_combout  $ (\portb~62_combout  $ (\Add1~3 )))) # (GND)
// \Add1~5  = CARRY((\porta~55_combout  & ((!\Add1~3 ) # (!\portb~62_combout ))) # (!\porta~55_combout  & (!\portb~62_combout  & !\Add1~3 )))

	.dataa(porta),
	.datab(portb29),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add1~3 ),
	.combout(\Add1~4_combout ),
	.cout(\Add1~5 ));
// synopsys translate_off
defparam \Add1~4 .lut_mask = 16'h962B;
defparam \Add1~4 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X57_Y40_N6
cycloneive_lcell_comb \Add1~6 (
// Equation(s):
// \Add1~6_combout  = (\portb~64_combout  & ((\porta~61_combout  & (!\Add1~5 )) # (!\porta~61_combout  & ((\Add1~5 ) # (GND))))) # (!\portb~64_combout  & ((\porta~61_combout  & (\Add1~5  & VCC)) # (!\porta~61_combout  & (!\Add1~5 ))))
// \Add1~7  = CARRY((\portb~64_combout  & ((!\Add1~5 ) # (!\porta~61_combout ))) # (!\portb~64_combout  & (!\porta~61_combout  & !\Add1~5 )))

	.dataa(portb30),
	.datab(porta3),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add1~5 ),
	.combout(\Add1~6_combout ),
	.cout(\Add1~7 ));
// synopsys translate_off
defparam \Add1~6 .lut_mask = 16'h692B;
defparam \Add1~6 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X52_Y38_N4
cycloneive_lcell_comb \Add0~4 (
// Equation(s):
// \Add0~4_combout  = ((\porta~55_combout  $ (\portb~62_combout  $ (!\Add0~3 )))) # (GND)
// \Add0~5  = CARRY((\porta~55_combout  & ((\portb~62_combout ) # (!\Add0~3 ))) # (!\porta~55_combout  & (\portb~62_combout  & !\Add0~3 )))

	.dataa(porta),
	.datab(portb29),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add0~3 ),
	.combout(\Add0~4_combout ),
	.cout(\Add0~5 ));
// synopsys translate_off
defparam \Add0~4 .lut_mask = 16'h698E;
defparam \Add0~4 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X52_Y38_N6
cycloneive_lcell_comb \Add0~6 (
// Equation(s):
// \Add0~6_combout  = (\portb~64_combout  & ((\porta~61_combout  & (\Add0~5  & VCC)) # (!\porta~61_combout  & (!\Add0~5 )))) # (!\portb~64_combout  & ((\porta~61_combout  & (!\Add0~5 )) # (!\porta~61_combout  & ((\Add0~5 ) # (GND)))))
// \Add0~7  = CARRY((\portb~64_combout  & (!\porta~61_combout  & !\Add0~5 )) # (!\portb~64_combout  & ((!\Add0~5 ) # (!\porta~61_combout ))))

	.dataa(portb30),
	.datab(porta3),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add0~5 ),
	.combout(\Add0~6_combout ),
	.cout(\Add0~7 ));
// synopsys translate_off
defparam \Add0~6 .lut_mask = 16'h9617;
defparam \Add0~6 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X52_Y40_N28
cycloneive_lcell_comb \Selector28~0 (
// Equation(s):
// \Selector28~0_combout  = (\Selector0~8_combout  & ((\Add1~6_combout ) # ((\Selector0~9_combout  & \Add0~6_combout )))) # (!\Selector0~8_combout  & (\Selector0~9_combout  & ((\Add0~6_combout ))))

	.dataa(\Selector0~8_combout ),
	.datab(\Selector0~9_combout ),
	.datac(\Add1~6_combout ),
	.datad(\Add0~6_combout ),
	.cin(gnd),
	.combout(\Selector28~0_combout ),
	.cout());
// synopsys translate_off
defparam \Selector28~0 .lut_mask = 16'hECA0;
defparam \Selector28~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X52_Y40_N2
cycloneive_lcell_comb \Selector28~4 (
// Equation(s):
// \Selector28~4_combout  = (\Selector28~0_combout ) # ((\Selector28~1_combout  & \Selector28~3_combout ))

	.dataa(gnd),
	.datab(\Selector28~1_combout ),
	.datac(\Selector28~3_combout ),
	.datad(\Selector28~0_combout ),
	.cin(gnd),
	.combout(\Selector28~4_combout ),
	.cout());
// synopsys translate_off
defparam \Selector28~4 .lut_mask = 16'hFFC0;
defparam \Selector28~4 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y38_N24
cycloneive_lcell_comb \ShiftRight0~78 (
// Equation(s):
// \ShiftRight0~78_combout  = (\porta~104_combout  & (!\portb~60_combout  & !\portb~58_combout ))

	.dataa(porta20),
	.datab(portb28),
	.datac(portb27),
	.datad(gnd),
	.cin(gnd),
	.combout(\ShiftRight0~78_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftRight0~78 .lut_mask = 16'h0202;
defparam \ShiftRight0~78 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y42_N16
cycloneive_lcell_comb \ShiftRight0~79 (
// Equation(s):
// \ShiftRight0~79_combout  = (\portb~60_combout  & ((\portb~58_combout  & ((\porta~106_combout ))) # (!\portb~58_combout  & (\porta~105_combout ))))

	.dataa(portb28),
	.datab(portb27),
	.datac(porta21),
	.datad(porta22),
	.cin(gnd),
	.combout(\ShiftRight0~79_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftRight0~79 .lut_mask = 16'hA820;
defparam \ShiftRight0~79 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y42_N6
cycloneive_lcell_comb \ShiftRight0~80 (
// Equation(s):
// \ShiftRight0~80_combout  = (\ShiftRight0~79_combout ) # ((\ShiftRight0~29_combout  & !\portb~60_combout ))

	.dataa(gnd),
	.datab(\ShiftRight0~29_combout ),
	.datac(portb28),
	.datad(\ShiftRight0~79_combout ),
	.cin(gnd),
	.combout(\ShiftRight0~80_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftRight0~80 .lut_mask = 16'hFF0C;
defparam \ShiftRight0~80 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y38_N22
cycloneive_lcell_comb \ShiftRight0~81 (
// Equation(s):
// \ShiftRight0~81_combout  = (\portb~62_combout  & (\ShiftRight0~78_combout )) # (!\portb~62_combout  & ((\ShiftRight0~80_combout )))

	.dataa(gnd),
	.datab(\ShiftRight0~78_combout ),
	.datac(portb29),
	.datad(\ShiftRight0~80_combout ),
	.cin(gnd),
	.combout(\ShiftRight0~81_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftRight0~81 .lut_mask = 16'hCFC0;
defparam \ShiftRight0~81 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y42_N14
cycloneive_lcell_comb \ShiftRight0~83 (
// Equation(s):
// \ShiftRight0~83_combout  = (\portb~60_combout  & (\ShiftRight0~34_combout )) # (!\portb~60_combout  & ((\ShiftRight0~36_combout )))

	.dataa(portb28),
	.datab(gnd),
	.datac(\ShiftRight0~34_combout ),
	.datad(\ShiftRight0~36_combout ),
	.cin(gnd),
	.combout(\ShiftRight0~83_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftRight0~83 .lut_mask = 16'hF5A0;
defparam \ShiftRight0~83 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y42_N24
cycloneive_lcell_comb \ShiftRight0~82 (
// Equation(s):
// \ShiftRight0~82_combout  = (\portb~60_combout  & (\ShiftRight0~30_combout )) # (!\portb~60_combout  & ((\ShiftRight0~33_combout )))

	.dataa(portb28),
	.datab(gnd),
	.datac(\ShiftRight0~30_combout ),
	.datad(\ShiftRight0~33_combout ),
	.cin(gnd),
	.combout(\ShiftRight0~82_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftRight0~82 .lut_mask = 16'hF5A0;
defparam \ShiftRight0~82 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y42_N28
cycloneive_lcell_comb \Selector20~0 (
// Equation(s):
// \Selector20~0_combout  = (\portb~62_combout  & ((\ShiftRight0~82_combout ))) # (!\portb~62_combout  & (\ShiftRight0~83_combout ))

	.dataa(portb29),
	.datab(gnd),
	.datac(\ShiftRight0~83_combout ),
	.datad(\ShiftRight0~82_combout ),
	.cin(gnd),
	.combout(\Selector20~0_combout ),
	.cout());
// synopsys translate_off
defparam \Selector20~0 .lut_mask = 16'hFA50;
defparam \Selector20~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y40_N2
cycloneive_lcell_comb \ShiftRight0~84 (
// Equation(s):
// \ShiftRight0~84_combout  = (\portb~64_combout  & (\ShiftRight0~81_combout )) # (!\portb~64_combout  & ((\Selector20~0_combout )))

	.dataa(portb30),
	.datab(gnd),
	.datac(\ShiftRight0~81_combout ),
	.datad(\Selector20~0_combout ),
	.cin(gnd),
	.combout(\ShiftRight0~84_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftRight0~84 .lut_mask = 16'hF5A0;
defparam \ShiftRight0~84 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y37_N20
cycloneive_lcell_comb \ShiftLeft0~3 (
// Equation(s):
// \ShiftLeft0~3_combout  = (\portb~58_combout  & (\porta~55_combout )) # (!\portb~58_combout  & ((\porta~61_combout )))

	.dataa(portb27),
	.datab(gnd),
	.datac(porta),
	.datad(porta3),
	.cin(gnd),
	.combout(\ShiftLeft0~3_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftLeft0~3 .lut_mask = 16'hF5A0;
defparam \ShiftLeft0~3 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y37_N30
cycloneive_lcell_comb \ShiftLeft0~4 (
// Equation(s):
// \ShiftLeft0~4_combout  = (\portb~60_combout  & ((\ShiftLeft0~2_combout ))) # (!\portb~60_combout  & (\ShiftLeft0~3_combout ))

	.dataa(gnd),
	.datab(\ShiftLeft0~3_combout ),
	.datac(portb28),
	.datad(\ShiftLeft0~2_combout ),
	.cin(gnd),
	.combout(\ShiftLeft0~4_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftLeft0~4 .lut_mask = 16'hFC0C;
defparam \ShiftLeft0~4 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X50_Y35_N26
cycloneive_lcell_comb \Selector0~12 (
// Equation(s):
// \Selector0~12_combout  = (plif_idexaluop_l_2 & (!plif_idexaluop_l_3 & (plif_idexaluop_l_1 & plif_idexaluop_l_0)))

	.dataa(plif_idexaluop_l_2),
	.datab(plif_idexaluop_l_3),
	.datac(plif_idexaluop_l_1),
	.datad(plif_idexaluop_l_0),
	.cin(gnd),
	.combout(\Selector0~12_combout ),
	.cout());
// synopsys translate_off
defparam \Selector0~12 .lut_mask = 16'h2000;
defparam \Selector0~12 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X50_Y36_N24
cycloneive_lcell_comb \Selector28~6 (
// Equation(s):
// \Selector28~6_combout  = (\porta~61_combout  & (\Selector0~10_combout )) # (!\porta~61_combout  & (((!\portb~64_combout  & \Selector0~12_combout ))))

	.dataa(\Selector0~10_combout ),
	.datab(portb30),
	.datac(porta3),
	.datad(\Selector0~12_combout ),
	.cin(gnd),
	.combout(\Selector28~6_combout ),
	.cout());
// synopsys translate_off
defparam \Selector28~6 .lut_mask = 16'hA3A0;
defparam \Selector28~6 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X50_Y36_N22
cycloneive_lcell_comb \Selector28~7 (
// Equation(s):
// \Selector28~7_combout  = (\Selector28~6_combout ) # ((\Selector0~13_combout  & (\portb~64_combout  $ (\porta~61_combout ))))

	.dataa(\Selector0~13_combout ),
	.datab(portb30),
	.datac(porta3),
	.datad(\Selector28~6_combout ),
	.cin(gnd),
	.combout(\Selector28~7_combout ),
	.cout());
// synopsys translate_off
defparam \Selector28~7 .lut_mask = 16'hFF28;
defparam \Selector28~7 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X50_Y38_N28
cycloneive_lcell_comb \ShiftRight0~74 (
// Equation(s):
// \ShiftRight0~74_combout  = (!\portb~64_combout  & !\portb~62_combout )

	.dataa(gnd),
	.datab(portb30),
	.datac(gnd),
	.datad(portb29),
	.cin(gnd),
	.combout(\ShiftRight0~74_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftRight0~74 .lut_mask = 16'h0033;
defparam \ShiftRight0~74 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y37_N4
cycloneive_lcell_comb \Selector28~8 (
// Equation(s):
// \Selector28~8_combout  = (\Selector0~14_combout  & (!\portb~66_combout  & (!\ShiftRight0~72_combout  & \ShiftRight0~74_combout )))

	.dataa(\Selector0~14_combout ),
	.datab(portb31),
	.datac(\ShiftRight0~72_combout ),
	.datad(\ShiftRight0~74_combout ),
	.cin(gnd),
	.combout(\Selector28~8_combout ),
	.cout());
// synopsys translate_off
defparam \Selector28~8 .lut_mask = 16'h0200;
defparam \Selector28~8 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X50_Y35_N18
cycloneive_lcell_comb \Selector0~10 (
// Equation(s):
// \Selector0~10_combout  = (plif_idexaluop_l_2 & (!plif_idexaluop_l_3 & (!plif_idexaluop_l_1 & plif_idexaluop_l_0)))

	.dataa(plif_idexaluop_l_2),
	.datab(plif_idexaluop_l_3),
	.datac(plif_idexaluop_l_1),
	.datad(plif_idexaluop_l_0),
	.cin(gnd),
	.combout(\Selector0~10_combout ),
	.cout());
// synopsys translate_off
defparam \Selector0~10 .lut_mask = 16'h0200;
defparam \Selector0~10 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X50_Y35_N16
cycloneive_lcell_comb \Selector0~11 (
// Equation(s):
// \Selector0~11_combout  = (plif_idexaluop_l_2 & (!plif_idexaluop_l_3 & (!plif_idexaluop_l_1 & !plif_idexaluop_l_0)))

	.dataa(plif_idexaluop_l_2),
	.datab(plif_idexaluop_l_3),
	.datac(plif_idexaluop_l_1),
	.datad(plif_idexaluop_l_0),
	.cin(gnd),
	.combout(\Selector0~11_combout ),
	.cout());
// synopsys translate_off
defparam \Selector0~11 .lut_mask = 16'h0002;
defparam \Selector0~11 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y37_N26
cycloneive_lcell_comb \Selector28~5 (
// Equation(s):
// \Selector28~5_combout  = (\portb~64_combout  & ((\Selector0~10_combout ) # ((\Selector0~11_combout  & \porta~61_combout ))))

	.dataa(portb30),
	.datab(\Selector0~10_combout ),
	.datac(\Selector0~11_combout ),
	.datad(porta3),
	.cin(gnd),
	.combout(\Selector28~5_combout ),
	.cout());
// synopsys translate_off
defparam \Selector28~5 .lut_mask = 16'hA888;
defparam \Selector28~5 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y37_N18
cycloneive_lcell_comb \Selector28~9 (
// Equation(s):
// \Selector28~9_combout  = (\Selector28~7_combout ) # ((\Selector28~5_combout ) # ((\ShiftLeft0~4_combout  & \Selector28~8_combout )))

	.dataa(\ShiftLeft0~4_combout ),
	.datab(\Selector28~7_combout ),
	.datac(\Selector28~8_combout ),
	.datad(\Selector28~5_combout ),
	.cin(gnd),
	.combout(\Selector28~9_combout ),
	.cout());
// synopsys translate_off
defparam \Selector28~9 .lut_mask = 16'hFFEC;
defparam \Selector28~9 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y38_N0
cycloneive_lcell_comb \Selector16~0 (
// Equation(s):
// \Selector16~0_combout  = (\Selector0~14_combout  & (!\portb~66_combout  & (!\ShiftRight0~41_combout  & !\ShiftRight0~8_combout )))

	.dataa(\Selector0~14_combout ),
	.datab(portb31),
	.datac(\ShiftRight0~41_combout ),
	.datad(\ShiftRight0~8_combout ),
	.cin(gnd),
	.combout(\Selector16~0_combout ),
	.cout());
// synopsys translate_off
defparam \Selector16~0 .lut_mask = 16'h0002;
defparam \Selector16~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y41_N4
cycloneive_lcell_comb \ShiftLeft0~5 (
// Equation(s):
// \ShiftLeft0~5_combout  = (!\portb~58_combout  & ((\portb~60_combout  & ((\porta~91_combout ))) # (!\portb~60_combout  & (\porta~55_combout ))))

	.dataa(porta),
	.datab(portb27),
	.datac(porta7),
	.datad(portb28),
	.cin(gnd),
	.combout(\ShiftLeft0~5_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftLeft0~5 .lut_mask = 16'h3022;
defparam \ShiftLeft0~5 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y41_N10
cycloneive_lcell_comb \ShiftLeft0~6 (
// Equation(s):
// \ShiftLeft0~6_combout  = (\ShiftLeft0~5_combout ) # ((\porta~57_combout  & (\portb~58_combout  & !\portb~60_combout )))

	.dataa(porta1),
	.datab(portb27),
	.datac(\ShiftLeft0~5_combout ),
	.datad(portb28),
	.cin(gnd),
	.combout(\ShiftLeft0~6_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftLeft0~6 .lut_mask = 16'hF0F8;
defparam \ShiftLeft0~6 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X52_Y40_N14
cycloneive_lcell_comb \Selector29~0 (
// Equation(s):
// \Selector29~0_combout  = (!\portb~64_combout  & (!\portb~62_combout  & (\Selector16~0_combout  & \ShiftLeft0~6_combout )))

	.dataa(portb30),
	.datab(portb29),
	.datac(\Selector16~0_combout ),
	.datad(\ShiftLeft0~6_combout ),
	.cin(gnd),
	.combout(\Selector29~0_combout ),
	.cout());
// synopsys translate_off
defparam \Selector29~0 .lut_mask = 16'h1000;
defparam \Selector29~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y36_N16
cycloneive_lcell_comb \ShiftRight0~92 (
// Equation(s):
// \ShiftRight0~92_combout  = (\portb~60_combout  & ((\ShiftRight0~65_combout ))) # (!\portb~60_combout  & (\ShiftRight0~67_combout ))

	.dataa(gnd),
	.datab(\ShiftRight0~67_combout ),
	.datac(portb28),
	.datad(\ShiftRight0~65_combout ),
	.cin(gnd),
	.combout(\ShiftRight0~92_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftRight0~92 .lut_mask = 16'hFC0C;
defparam \ShiftRight0~92 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y39_N28
cycloneive_lcell_comb \ShiftRight0~91 (
// Equation(s):
// \ShiftRight0~91_combout  = (\portb~60_combout  & ((\ShiftRight0~61_combout ))) # (!\portb~60_combout  & (\ShiftRight0~64_combout ))

	.dataa(gnd),
	.datab(portb28),
	.datac(\ShiftRight0~64_combout ),
	.datad(\ShiftRight0~61_combout ),
	.cin(gnd),
	.combout(\ShiftRight0~91_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftRight0~91 .lut_mask = 16'hFC30;
defparam \ShiftRight0~91 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y39_N26
cycloneive_lcell_comb \Selector21~0 (
// Equation(s):
// \Selector21~0_combout  = (\portb~62_combout  & ((\ShiftRight0~91_combout ))) # (!\portb~62_combout  & (\ShiftRight0~92_combout ))

	.dataa(portb29),
	.datab(gnd),
	.datac(\ShiftRight0~92_combout ),
	.datad(\ShiftRight0~91_combout ),
	.cin(gnd),
	.combout(\Selector21~0_combout ),
	.cout());
// synopsys translate_off
defparam \Selector21~0 .lut_mask = 16'hFA50;
defparam \Selector21~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y39_N10
cycloneive_lcell_comb \ShiftRight0~89 (
// Equation(s):
// \ShiftRight0~89_combout  = (\portb~60_combout  & ((\ShiftRight0~58_combout ))) # (!\portb~60_combout  & (\ShiftRight0~60_combout ))

	.dataa(gnd),
	.datab(portb28),
	.datac(\ShiftRight0~60_combout ),
	.datad(\ShiftRight0~58_combout ),
	.cin(gnd),
	.combout(\ShiftRight0~89_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftRight0~89 .lut_mask = 16'hFC30;
defparam \ShiftRight0~89 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y40_N28
cycloneive_lcell_comb \ShiftRight0~90 (
// Equation(s):
// \ShiftRight0~90_combout  = (\portb~62_combout  & (!\portb~60_combout  & ((\ShiftRight0~57_combout )))) # (!\portb~62_combout  & (((\ShiftRight0~89_combout ))))

	.dataa(portb28),
	.datab(portb29),
	.datac(\ShiftRight0~89_combout ),
	.datad(\ShiftRight0~57_combout ),
	.cin(gnd),
	.combout(\ShiftRight0~90_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftRight0~90 .lut_mask = 16'h7430;
defparam \ShiftRight0~90 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y37_N14
cycloneive_lcell_comb \ShiftRight0~93 (
// Equation(s):
// \ShiftRight0~93_combout  = (\portb~64_combout  & ((\ShiftRight0~90_combout ))) # (!\portb~64_combout  & (\Selector21~0_combout ))

	.dataa(gnd),
	.datab(portb30),
	.datac(\Selector21~0_combout ),
	.datad(\ShiftRight0~90_combout ),
	.cin(gnd),
	.combout(\ShiftRight0~93_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftRight0~93 .lut_mask = 16'hFC30;
defparam \ShiftRight0~93 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X50_Y35_N28
cycloneive_lcell_comb \Selector0~13 (
// Equation(s):
// \Selector0~13_combout  = (plif_idexaluop_l_2 & (!plif_idexaluop_l_3 & (plif_idexaluop_l_1 & !plif_idexaluop_l_0)))

	.dataa(plif_idexaluop_l_2),
	.datab(plif_idexaluop_l_3),
	.datac(plif_idexaluop_l_1),
	.datad(plif_idexaluop_l_0),
	.cin(gnd),
	.combout(\Selector0~13_combout ),
	.cout());
// synopsys translate_off
defparam \Selector0~13 .lut_mask = 16'h0020;
defparam \Selector0~13 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X50_Y36_N8
cycloneive_lcell_comb \Selector29~2 (
// Equation(s):
// \Selector29~2_combout  = (\porta~55_combout  & (\Selector0~11_combout )) # (!\porta~55_combout  & ((\Selector0~12_combout )))

	.dataa(\Selector0~11_combout ),
	.datab(\Selector0~12_combout ),
	.datac(porta),
	.datad(gnd),
	.cin(gnd),
	.combout(\Selector29~2_combout ),
	.cout());
// synopsys translate_off
defparam \Selector29~2 .lut_mask = 16'hACAC;
defparam \Selector29~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X50_Y36_N18
cycloneive_lcell_comb \Selector29~3 (
// Equation(s):
// \Selector29~3_combout  = (\porta~55_combout  & ((\Selector0~10_combout ) # (!\portb~62_combout ))) # (!\porta~55_combout  & ((\portb~62_combout )))

	.dataa(\Selector0~10_combout ),
	.datab(gnd),
	.datac(porta),
	.datad(portb29),
	.cin(gnd),
	.combout(\Selector29~3_combout ),
	.cout());
// synopsys translate_off
defparam \Selector29~3 .lut_mask = 16'hAFF0;
defparam \Selector29~3 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X50_Y36_N20
cycloneive_lcell_comb \Selector29~4 (
// Equation(s):
// \Selector29~4_combout  = (\Selector29~3_combout  & ((\Selector0~10_combout ) # ((\Selector0~13_combout )))) # (!\Selector29~3_combout  & (((\Selector29~2_combout ))))

	.dataa(\Selector0~10_combout ),
	.datab(\Selector0~13_combout ),
	.datac(\Selector29~2_combout ),
	.datad(\Selector29~3_combout ),
	.cin(gnd),
	.combout(\Selector29~4_combout ),
	.cout());
// synopsys translate_off
defparam \Selector29~4 .lut_mask = 16'hEEF0;
defparam \Selector29~4 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X52_Y41_N4
cycloneive_lcell_comb \ShiftRight0~46 (
// Equation(s):
// \ShiftRight0~46_combout  = (\portb~58_combout  & (\porta~95_combout )) # (!\portb~58_combout  & ((\porta~59_combout )))

	.dataa(portb27),
	.datab(gnd),
	.datac(porta11),
	.datad(porta2),
	.cin(gnd),
	.combout(\ShiftRight0~46_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftRight0~46 .lut_mask = 16'hF5A0;
defparam \ShiftRight0~46 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y36_N8
cycloneive_lcell_comb \ShiftRight0~87 (
// Equation(s):
// \ShiftRight0~87_combout  = (\portb~60_combout  & (\ShiftRight0~50_combout )) # (!\portb~60_combout  & ((\ShiftRight0~52_combout )))

	.dataa(gnd),
	.datab(\ShiftRight0~50_combout ),
	.datac(portb28),
	.datad(\ShiftRight0~52_combout ),
	.cin(gnd),
	.combout(\ShiftRight0~87_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftRight0~87 .lut_mask = 16'hCFC0;
defparam \ShiftRight0~87 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y36_N18
cycloneive_lcell_comb \ShiftRight0~86 (
// Equation(s):
// \ShiftRight0~86_combout  = (\portb~60_combout  & (\ShiftRight0~68_combout )) # (!\portb~60_combout  & ((\ShiftRight0~49_combout )))

	.dataa(gnd),
	.datab(\ShiftRight0~68_combout ),
	.datac(portb28),
	.datad(\ShiftRight0~49_combout ),
	.cin(gnd),
	.combout(\ShiftRight0~86_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftRight0~86 .lut_mask = 16'hCFC0;
defparam \ShiftRight0~86 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y36_N26
cycloneive_lcell_comb \ShiftRight0~88 (
// Equation(s):
// \ShiftRight0~88_combout  = (\portb~62_combout  & ((\ShiftRight0~86_combout ))) # (!\portb~62_combout  & (\ShiftRight0~87_combout ))

	.dataa(portb29),
	.datab(gnd),
	.datac(\ShiftRight0~87_combout ),
	.datad(\ShiftRight0~86_combout ),
	.cin(gnd),
	.combout(\ShiftRight0~88_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftRight0~88 .lut_mask = 16'hFA50;
defparam \ShiftRight0~88 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X52_Y40_N8
cycloneive_lcell_comb \Selector29~6 (
// Equation(s):
// \Selector29~6_combout  = (\Selector29~5_combout  & (((\ShiftRight0~88_combout ) # (!\Selector3~1_combout )))) # (!\Selector29~5_combout  & (\ShiftRight0~46_combout  & ((\Selector3~1_combout ))))

	.dataa(\Selector29~5_combout ),
	.datab(\ShiftRight0~46_combout ),
	.datac(\ShiftRight0~88_combout ),
	.datad(\Selector3~1_combout ),
	.cin(gnd),
	.combout(\Selector29~6_combout ),
	.cout());
// synopsys translate_off
defparam \Selector29~6 .lut_mask = 16'hE4AA;
defparam \Selector29~6 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X52_Y40_N0
cycloneive_lcell_comb \Selector29~1 (
// Equation(s):
// \Selector29~1_combout  = (\Selector0~8_combout  & ((\Add1~4_combout ) # ((\Selector0~9_combout  & \Add0~4_combout )))) # (!\Selector0~8_combout  & (\Selector0~9_combout  & ((\Add0~4_combout ))))

	.dataa(\Selector0~8_combout ),
	.datab(\Selector0~9_combout ),
	.datac(\Add1~4_combout ),
	.datad(\Add0~4_combout ),
	.cin(gnd),
	.combout(\Selector29~1_combout ),
	.cout());
// synopsys translate_off
defparam \Selector29~1 .lut_mask = 16'hECA0;
defparam \Selector29~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X52_Y40_N18
cycloneive_lcell_comb \Selector29~7 (
// Equation(s):
// \Selector29~7_combout  = (\Selector29~4_combout ) # ((\Selector29~1_combout ) # ((\Selector28~1_combout  & \Selector29~6_combout )))

	.dataa(\Selector29~4_combout ),
	.datab(\Selector28~1_combout ),
	.datac(\Selector29~6_combout ),
	.datad(\Selector29~1_combout ),
	.cin(gnd),
	.combout(\Selector29~7_combout ),
	.cout());
// synopsys translate_off
defparam \Selector29~7 .lut_mask = 16'hFFEA;
defparam \Selector29~7 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X50_Y41_N26
cycloneive_lcell_comb \Selector26~5 (
// Equation(s):
// \Selector26~5_combout  = (\portb~56_combout  & ((\Selector0~3_combout ) # ((\Selector0~4_combout  & \porta~95_combout ))))

	.dataa(portb26),
	.datab(\Selector0~4_combout ),
	.datac(porta11),
	.datad(\Selector0~3_combout ),
	.cin(gnd),
	.combout(\Selector26~5_combout ),
	.cout());
// synopsys translate_off
defparam \Selector26~5 .lut_mask = 16'hAA80;
defparam \Selector26~5 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y42_N24
cycloneive_lcell_comb \Selector26~6 (
// Equation(s):
// \Selector26~6_combout  = (\porta~95_combout  & (((\Selector0~3_combout )))) # (!\porta~95_combout  & (\Selector0~7_combout  & (!\portb~56_combout )))

	.dataa(\Selector0~7_combout ),
	.datab(porta11),
	.datac(portb26),
	.datad(\Selector0~3_combout ),
	.cin(gnd),
	.combout(\Selector26~6_combout ),
	.cout());
// synopsys translate_off
defparam \Selector26~6 .lut_mask = 16'hCE02;
defparam \Selector26~6 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y42_N30
cycloneive_lcell_comb \Selector26~7 (
// Equation(s):
// \Selector26~7_combout  = (\Selector26~6_combout ) # ((\Selector0~2_combout  & (\porta~95_combout  $ (\portb~56_combout ))))

	.dataa(porta11),
	.datab(\Selector0~2_combout ),
	.datac(portb26),
	.datad(\Selector26~6_combout ),
	.cin(gnd),
	.combout(\Selector26~7_combout ),
	.cout());
// synopsys translate_off
defparam \Selector26~7 .lut_mask = 16'hFF48;
defparam \Selector26~7 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y38_N0
cycloneive_lcell_comb \Selector1~1 (
// Equation(s):
// \Selector1~1_combout  = (\ShiftRight0~8_combout ) # ((\ShiftRight0~9_combout ) # ((\portb~66_combout ) # (\ShiftRight0~11_combout )))

	.dataa(\ShiftRight0~8_combout ),
	.datab(\ShiftRight0~9_combout ),
	.datac(portb31),
	.datad(\ShiftRight0~11_combout ),
	.cin(gnd),
	.combout(\Selector1~1_combout ),
	.cout());
// synopsys translate_off
defparam \Selector1~1 .lut_mask = 16'hFFFE;
defparam \Selector1~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y37_N0
cycloneive_lcell_comb \ShiftLeft0~7 (
// Equation(s):
// \ShiftLeft0~7_combout  = (\portb~58_combout  & ((\porta~59_combout ))) # (!\portb~58_combout  & (\porta~95_combout ))

	.dataa(gnd),
	.datab(portb27),
	.datac(porta11),
	.datad(porta2),
	.cin(gnd),
	.combout(\ShiftLeft0~7_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftLeft0~7 .lut_mask = 16'hFC30;
defparam \ShiftLeft0~7 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y38_N4
cycloneive_lcell_comb \ShiftLeft0~8 (
// Equation(s):
// \ShiftLeft0~8_combout  = (\portb~60_combout  & ((\ShiftLeft0~3_combout ))) # (!\portb~60_combout  & (\ShiftLeft0~7_combout ))

	.dataa(portb28),
	.datab(\ShiftLeft0~7_combout ),
	.datac(gnd),
	.datad(\ShiftLeft0~3_combout ),
	.cin(gnd),
	.combout(\ShiftLeft0~8_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftLeft0~8 .lut_mask = 16'hEE44;
defparam \ShiftLeft0~8 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y38_N2
cycloneive_lcell_comb \ShiftLeft0~9 (
// Equation(s):
// \ShiftLeft0~9_combout  = (\portb~62_combout  & (\ShiftLeft0~2_combout  & ((!\portb~60_combout )))) # (!\portb~62_combout  & (((\ShiftLeft0~8_combout ))))

	.dataa(portb29),
	.datab(\ShiftLeft0~2_combout ),
	.datac(\ShiftLeft0~8_combout ),
	.datad(portb28),
	.cin(gnd),
	.combout(\ShiftLeft0~9_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftLeft0~9 .lut_mask = 16'h50D8;
defparam \ShiftLeft0~9 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X50_Y41_N14
cycloneive_lcell_comb \Selector26~0 (
// Equation(s):
// \Selector26~0_combout  = (!\portb~64_combout  & (\Selector0~1_combout  & (!\Selector1~1_combout  & \ShiftLeft0~9_combout )))

	.dataa(portb30),
	.datab(\Selector0~1_combout ),
	.datac(\Selector1~1_combout ),
	.datad(\ShiftLeft0~9_combout ),
	.cin(gnd),
	.combout(\Selector26~0_combout ),
	.cout());
// synopsys translate_off
defparam \Selector26~0 .lut_mask = 16'h0400;
defparam \Selector26~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y40_N8
cycloneive_lcell_comb \Add1~8 (
// Equation(s):
// \Add1~8_combout  = ((\porta~59_combout  $ (\portb~66_combout  $ (\Add1~7 )))) # (GND)
// \Add1~9  = CARRY((\porta~59_combout  & ((!\Add1~7 ) # (!\portb~66_combout ))) # (!\porta~59_combout  & (!\portb~66_combout  & !\Add1~7 )))

	.dataa(porta2),
	.datab(portb31),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add1~7 ),
	.combout(\Add1~8_combout ),
	.cout(\Add1~9 ));
// synopsys translate_off
defparam \Add1~8 .lut_mask = 16'h962B;
defparam \Add1~8 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X57_Y40_N10
cycloneive_lcell_comb \Add1~10 (
// Equation(s):
// \Add1~10_combout  = (\porta~95_combout  & ((\portb~56_combout  & (!\Add1~9 )) # (!\portb~56_combout  & (\Add1~9  & VCC)))) # (!\porta~95_combout  & ((\portb~56_combout  & ((\Add1~9 ) # (GND))) # (!\portb~56_combout  & (!\Add1~9 ))))
// \Add1~11  = CARRY((\porta~95_combout  & (\portb~56_combout  & !\Add1~9 )) # (!\porta~95_combout  & ((\portb~56_combout ) # (!\Add1~9 ))))

	.dataa(porta11),
	.datab(portb26),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add1~9 ),
	.combout(\Add1~10_combout ),
	.cout(\Add1~11 ));
// synopsys translate_off
defparam \Add1~10 .lut_mask = 16'h694D;
defparam \Add1~10 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X52_Y38_N8
cycloneive_lcell_comb \Add0~8 (
// Equation(s):
// \Add0~8_combout  = ((\portb~66_combout  $ (\porta~59_combout  $ (!\Add0~7 )))) # (GND)
// \Add0~9  = CARRY((\portb~66_combout  & ((\porta~59_combout ) # (!\Add0~7 ))) # (!\portb~66_combout  & (\porta~59_combout  & !\Add0~7 )))

	.dataa(portb31),
	.datab(porta2),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add0~7 ),
	.combout(\Add0~8_combout ),
	.cout(\Add0~9 ));
// synopsys translate_off
defparam \Add0~8 .lut_mask = 16'h698E;
defparam \Add0~8 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X52_Y38_N10
cycloneive_lcell_comb \Add0~10 (
// Equation(s):
// \Add0~10_combout  = (\portb~56_combout  & ((\porta~95_combout  & (\Add0~9  & VCC)) # (!\porta~95_combout  & (!\Add0~9 )))) # (!\portb~56_combout  & ((\porta~95_combout  & (!\Add0~9 )) # (!\porta~95_combout  & ((\Add0~9 ) # (GND)))))
// \Add0~11  = CARRY((\portb~56_combout  & (!\porta~95_combout  & !\Add0~9 )) # (!\portb~56_combout  & ((!\Add0~9 ) # (!\porta~95_combout ))))

	.dataa(portb26),
	.datab(porta11),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add0~9 ),
	.combout(\Add0~10_combout ),
	.cout(\Add0~11 ));
// synopsys translate_off
defparam \Add0~10 .lut_mask = 16'h9617;
defparam \Add0~10 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X50_Y41_N8
cycloneive_lcell_comb \Selector26~1 (
// Equation(s):
// \Selector26~1_combout  = (\Selector0~5_combout  & ((\Add0~10_combout ) # ((\Add1~10_combout  & \Selector0~6_combout )))) # (!\Selector0~5_combout  & (\Add1~10_combout  & (\Selector0~6_combout )))

	.dataa(\Selector0~5_combout ),
	.datab(\Add1~10_combout ),
	.datac(\Selector0~6_combout ),
	.datad(\Add0~10_combout ),
	.cin(gnd),
	.combout(\Selector26~1_combout ),
	.cout());
// synopsys translate_off
defparam \Selector26~1 .lut_mask = 16'hEAC0;
defparam \Selector26~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X52_Y41_N24
cycloneive_lcell_comb \ShiftRight0~17 (
// Equation(s):
// \ShiftRight0~17_combout  = (\portb~60_combout  & ((\ShiftRight0~15_combout ))) # (!\portb~60_combout  & (\ShiftRight0~16_combout ))

	.dataa(\ShiftRight0~16_combout ),
	.datab(\ShiftRight0~15_combout ),
	.datac(portb28),
	.datad(gnd),
	.cin(gnd),
	.combout(\ShiftRight0~17_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftRight0~17 .lut_mask = 16'hCACA;
defparam \ShiftRight0~17 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y40_N4
cycloneive_lcell_comb \Selector7~0 (
// Equation(s):
// \Selector7~0_combout  = (\portb~64_combout ) # (\portb~66_combout )

	.dataa(portb30),
	.datab(gnd),
	.datac(gnd),
	.datad(portb31),
	.cin(gnd),
	.combout(\Selector7~0_combout ),
	.cout());
// synopsys translate_off
defparam \Selector7~0 .lut_mask = 16'hFFAA;
defparam \Selector7~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X52_Y41_N22
cycloneive_lcell_comb \Selector26~2 (
// Equation(s):
// \Selector26~2_combout  = (\Selector7~1_combout  & (((\Selector7~0_combout ) # (\ShiftRight0~24_combout )))) # (!\Selector7~1_combout  & (\ShiftRight0~17_combout  & (!\Selector7~0_combout )))

	.dataa(\Selector7~1_combout ),
	.datab(\ShiftRight0~17_combout ),
	.datac(\Selector7~0_combout ),
	.datad(\ShiftRight0~24_combout ),
	.cin(gnd),
	.combout(\Selector26~2_combout ),
	.cout());
// synopsys translate_off
defparam \Selector26~2 .lut_mask = 16'hAEA4;
defparam \Selector26~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y41_N22
cycloneive_lcell_comb \ShiftRight0~95 (
// Equation(s):
// \ShiftRight0~95_combout  = (!\portb~62_combout  & ((\portb~64_combout  & ((\ShiftRight0~28_combout ))) # (!\portb~64_combout  & (\ShiftRight0~35_combout ))))

	.dataa(portb30),
	.datab(portb29),
	.datac(\ShiftRight0~35_combout ),
	.datad(\ShiftRight0~28_combout ),
	.cin(gnd),
	.combout(\ShiftRight0~95_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftRight0~95 .lut_mask = 16'h3210;
defparam \ShiftRight0~95 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y41_N4
cycloneive_lcell_comb \ShiftRight0~96 (
// Equation(s):
// \ShiftRight0~96_combout  = (\ShiftRight0~95_combout ) # ((!\portb~64_combout  & (\portb~62_combout  & \ShiftRight0~31_combout )))

	.dataa(portb30),
	.datab(portb29),
	.datac(\ShiftRight0~95_combout ),
	.datad(\ShiftRight0~31_combout ),
	.cin(gnd),
	.combout(\ShiftRight0~96_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftRight0~96 .lut_mask = 16'hF4F0;
defparam \ShiftRight0~96 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y38_N10
cycloneive_lcell_comb \ShiftRight0~21 (
// Equation(s):
// \ShiftRight0~21_combout  = (\portb~60_combout  & (\ShiftRight0~19_combout )) # (!\portb~60_combout  & ((\ShiftRight0~20_combout )))

	.dataa(portb28),
	.datab(gnd),
	.datac(\ShiftRight0~19_combout ),
	.datad(\ShiftRight0~20_combout ),
	.cin(gnd),
	.combout(\ShiftRight0~21_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftRight0~21 .lut_mask = 16'hF5A0;
defparam \ShiftRight0~21 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y38_N28
cycloneive_lcell_comb \ShiftRight0~94 (
// Equation(s):
// \ShiftRight0~94_combout  = (\portb~62_combout  & (\ShiftRight0~38_combout )) # (!\portb~62_combout  & ((\ShiftRight0~21_combout )))

	.dataa(portb29),
	.datab(\ShiftRight0~38_combout ),
	.datac(gnd),
	.datad(\ShiftRight0~21_combout ),
	.cin(gnd),
	.combout(\ShiftRight0~94_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftRight0~94 .lut_mask = 16'hDD88;
defparam \ShiftRight0~94 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X50_Y41_N6
cycloneive_lcell_comb \Selector26~3 (
// Equation(s):
// \Selector26~3_combout  = (\Selector7~0_combout  & ((\Selector26~2_combout  & (\ShiftRight0~96_combout )) # (!\Selector26~2_combout  & ((\ShiftRight0~94_combout ))))) # (!\Selector7~0_combout  & (\Selector26~2_combout ))

	.dataa(\Selector7~0_combout ),
	.datab(\Selector26~2_combout ),
	.datac(\ShiftRight0~96_combout ),
	.datad(\ShiftRight0~94_combout ),
	.cin(gnd),
	.combout(\Selector26~3_combout ),
	.cout());
// synopsys translate_off
defparam \Selector26~3 .lut_mask = 16'hE6C4;
defparam \Selector26~3 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X50_Y41_N12
cycloneive_lcell_comb \Selector26~4 (
// Equation(s):
// \Selector26~4_combout  = (\Selector26~1_combout ) # ((\Selector24~0_combout  & \Selector26~3_combout ))

	.dataa(\Selector24~0_combout ),
	.datab(gnd),
	.datac(\Selector26~1_combout ),
	.datad(\Selector26~3_combout ),
	.cin(gnd),
	.combout(\Selector26~4_combout ),
	.cout());
// synopsys translate_off
defparam \Selector26~4 .lut_mask = 16'hFAF0;
defparam \Selector26~4 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y40_N14
cycloneive_lcell_comb \ShiftLeft0~10 (
// Equation(s):
// \ShiftLeft0~10_combout  = (!\portb~58_combout  & (!\portb~60_combout  & \porta~91_combout ))

	.dataa(gnd),
	.datab(portb27),
	.datac(portb28),
	.datad(porta7),
	.cin(gnd),
	.combout(\ShiftLeft0~10_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftLeft0~10 .lut_mask = 16'h0300;
defparam \ShiftLeft0~10 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y40_N2
cycloneive_lcell_comb \ShiftLeft0~12 (
// Equation(s):
// \ShiftLeft0~12_combout  = (\portb~58_combout  & ((\porta~61_combout ))) # (!\portb~58_combout  & (\porta~59_combout ))

	.dataa(gnd),
	.datab(portb27),
	.datac(porta2),
	.datad(porta3),
	.cin(gnd),
	.combout(\ShiftLeft0~12_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftLeft0~12 .lut_mask = 16'hFC30;
defparam \ShiftLeft0~12 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y40_N20
cycloneive_lcell_comb \ShiftLeft0~11 (
// Equation(s):
// \ShiftLeft0~11_combout  = (\portb~60_combout  & ((\portb~58_combout  & ((\porta~57_combout ))) # (!\portb~58_combout  & (\porta~55_combout ))))

	.dataa(portb28),
	.datab(portb27),
	.datac(porta),
	.datad(porta1),
	.cin(gnd),
	.combout(\ShiftLeft0~11_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftLeft0~11 .lut_mask = 16'hA820;
defparam \ShiftLeft0~11 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y40_N12
cycloneive_lcell_comb \ShiftLeft0~13 (
// Equation(s):
// \ShiftLeft0~13_combout  = (\ShiftLeft0~11_combout ) # ((\ShiftLeft0~12_combout  & !\portb~60_combout ))

	.dataa(gnd),
	.datab(\ShiftLeft0~12_combout ),
	.datac(portb28),
	.datad(\ShiftLeft0~11_combout ),
	.cin(gnd),
	.combout(\ShiftLeft0~13_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftLeft0~13 .lut_mask = 16'hFF0C;
defparam \ShiftLeft0~13 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y40_N26
cycloneive_lcell_comb \ShiftLeft0~14 (
// Equation(s):
// \ShiftLeft0~14_combout  = (\portb~62_combout  & (\ShiftLeft0~10_combout )) # (!\portb~62_combout  & ((\ShiftLeft0~13_combout )))

	.dataa(gnd),
	.datab(portb29),
	.datac(\ShiftLeft0~10_combout ),
	.datad(\ShiftLeft0~13_combout ),
	.cin(gnd),
	.combout(\ShiftLeft0~14_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftLeft0~14 .lut_mask = 16'hF3C0;
defparam \ShiftLeft0~14 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X50_Y38_N30
cycloneive_lcell_comb \Selector27~0 (
// Equation(s):
// \Selector27~0_combout  = (\ShiftLeft0~14_combout  & (!\portb~64_combout  & (\Selector0~1_combout  & !\Selector1~1_combout )))

	.dataa(\ShiftLeft0~14_combout ),
	.datab(portb30),
	.datac(\Selector0~1_combout ),
	.datad(\Selector1~1_combout ),
	.cin(gnd),
	.combout(\Selector27~0_combout ),
	.cout());
// synopsys translate_off
defparam \Selector27~0 .lut_mask = 16'h0020;
defparam \Selector27~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X50_Y38_N8
cycloneive_lcell_comb \Selector27~5 (
// Equation(s):
// \Selector27~5_combout  = (\portb~66_combout  & ((\Selector0~3_combout ) # ((\Selector0~4_combout  & \porta~59_combout ))))

	.dataa(\Selector0~4_combout ),
	.datab(portb31),
	.datac(porta2),
	.datad(\Selector0~3_combout ),
	.cin(gnd),
	.combout(\Selector27~5_combout ),
	.cout());
// synopsys translate_off
defparam \Selector27~5 .lut_mask = 16'hCC80;
defparam \Selector27~5 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y42_N20
cycloneive_lcell_comb \Selector27~6 (
// Equation(s):
// \Selector27~6_combout  = (\porta~59_combout  & (((\Selector0~3_combout )))) # (!\porta~59_combout  & (\Selector0~7_combout  & (!\portb~66_combout )))

	.dataa(\Selector0~7_combout ),
	.datab(portb31),
	.datac(\Selector0~3_combout ),
	.datad(porta2),
	.cin(gnd),
	.combout(\Selector27~6_combout ),
	.cout());
// synopsys translate_off
defparam \Selector27~6 .lut_mask = 16'hF022;
defparam \Selector27~6 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y42_N6
cycloneive_lcell_comb \Selector27~7 (
// Equation(s):
// \Selector27~7_combout  = (\Selector27~6_combout ) # ((\Selector0~2_combout  & (\portb~66_combout  $ (\porta~59_combout ))))

	.dataa(\Selector27~6_combout ),
	.datab(\Selector0~2_combout ),
	.datac(portb31),
	.datad(porta2),
	.cin(gnd),
	.combout(\Selector27~7_combout ),
	.cout());
// synopsys translate_off
defparam \Selector27~7 .lut_mask = 16'hAEEA;
defparam \Selector27~7 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X50_Y38_N4
cycloneive_lcell_comb \Selector27~1 (
// Equation(s):
// \Selector27~1_combout  = (\Selector0~5_combout  & ((\Add0~8_combout ) # ((\Selector0~6_combout  & \Add1~8_combout )))) # (!\Selector0~5_combout  & (\Selector0~6_combout  & ((\Add1~8_combout ))))

	.dataa(\Selector0~5_combout ),
	.datab(\Selector0~6_combout ),
	.datac(\Add0~8_combout ),
	.datad(\Add1~8_combout ),
	.cin(gnd),
	.combout(\Selector27~1_combout ),
	.cout());
// synopsys translate_off
defparam \Selector27~1 .lut_mask = 16'hECA0;
defparam \Selector27~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y40_N26
cycloneive_lcell_comb \Selector7~1 (
// Equation(s):
// \Selector7~1_combout  = (\portb~66_combout ) # ((\portb~62_combout  & !\portb~64_combout ))

	.dataa(gnd),
	.datab(portb31),
	.datac(portb29),
	.datad(portb30),
	.cin(gnd),
	.combout(\Selector7~1_combout ),
	.cout());
// synopsys translate_off
defparam \Selector7~1 .lut_mask = 16'hCCFC;
defparam \Selector7~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y36_N18
cycloneive_lcell_comb \ShiftRight0~98 (
// Equation(s):
// \ShiftRight0~98_combout  = (!\portb~64_combout  & ((\portb~62_combout  & ((\ShiftRight0~62_combout ))) # (!\portb~62_combout  & (\ShiftRight0~66_combout ))))

	.dataa(portb29),
	.datab(portb30),
	.datac(\ShiftRight0~66_combout ),
	.datad(\ShiftRight0~62_combout ),
	.cin(gnd),
	.combout(\ShiftRight0~98_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftRight0~98 .lut_mask = 16'h3210;
defparam \ShiftRight0~98 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y36_N16
cycloneive_lcell_comb \ShiftRight0~99 (
// Equation(s):
// \ShiftRight0~99_combout  = (\ShiftRight0~98_combout ) # ((\ShiftRight0~59_combout  & (\portb~64_combout  & !\portb~62_combout )))

	.dataa(\ShiftRight0~59_combout ),
	.datab(portb30),
	.datac(portb29),
	.datad(\ShiftRight0~98_combout ),
	.cin(gnd),
	.combout(\ShiftRight0~99_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftRight0~99 .lut_mask = 16'hFF08;
defparam \ShiftRight0~99 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X52_Y41_N2
cycloneive_lcell_comb \ShiftRight0~45 (
// Equation(s):
// \ShiftRight0~45_combout  = (\portb~58_combout  & (\porta~93_combout )) # (!\portb~58_combout  & ((\porta~94_combout )))

	.dataa(porta9),
	.datab(gnd),
	.datac(porta10),
	.datad(portb27),
	.cin(gnd),
	.combout(\ShiftRight0~45_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftRight0~45 .lut_mask = 16'hAAF0;
defparam \ShiftRight0~45 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X52_Y41_N18
cycloneive_lcell_comb \ShiftRight0~47 (
// Equation(s):
// \ShiftRight0~47_combout  = (\portb~60_combout  & ((\ShiftRight0~45_combout ))) # (!\portb~60_combout  & (\ShiftRight0~46_combout ))

	.dataa(gnd),
	.datab(portb28),
	.datac(\ShiftRight0~46_combout ),
	.datad(\ShiftRight0~45_combout ),
	.cin(gnd),
	.combout(\ShiftRight0~47_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftRight0~47 .lut_mask = 16'hFC30;
defparam \ShiftRight0~47 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y40_N12
cycloneive_lcell_comb \ShiftRight0~97 (
// Equation(s):
// \ShiftRight0~97_combout  = (\portb~62_combout  & ((\ShiftRight0~69_combout ))) # (!\portb~62_combout  & (\ShiftRight0~51_combout ))

	.dataa(gnd),
	.datab(portb29),
	.datac(\ShiftRight0~51_combout ),
	.datad(\ShiftRight0~69_combout ),
	.cin(gnd),
	.combout(\ShiftRight0~97_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftRight0~97 .lut_mask = 16'hFC30;
defparam \ShiftRight0~97 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X50_Y38_N18
cycloneive_lcell_comb \Selector27~2 (
// Equation(s):
// \Selector27~2_combout  = (\Selector7~0_combout  & ((\Selector7~1_combout ) # ((\ShiftRight0~97_combout )))) # (!\Selector7~0_combout  & (!\Selector7~1_combout  & (\ShiftRight0~47_combout )))

	.dataa(\Selector7~0_combout ),
	.datab(\Selector7~1_combout ),
	.datac(\ShiftRight0~47_combout ),
	.datad(\ShiftRight0~97_combout ),
	.cin(gnd),
	.combout(\Selector27~2_combout ),
	.cout());
// synopsys translate_off
defparam \Selector27~2 .lut_mask = 16'hBA98;
defparam \Selector27~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X50_Y38_N0
cycloneive_lcell_comb \Selector27~3 (
// Equation(s):
// \Selector27~3_combout  = (\Selector7~1_combout  & ((\Selector27~2_combout  & ((\ShiftRight0~99_combout ))) # (!\Selector27~2_combout  & (\ShiftRight0~54_combout )))) # (!\Selector7~1_combout  & (((\Selector27~2_combout ))))

	.dataa(\ShiftRight0~54_combout ),
	.datab(\Selector7~1_combout ),
	.datac(\ShiftRight0~99_combout ),
	.datad(\Selector27~2_combout ),
	.cin(gnd),
	.combout(\Selector27~3_combout ),
	.cout());
// synopsys translate_off
defparam \Selector27~3 .lut_mask = 16'hF388;
defparam \Selector27~3 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X50_Y38_N2
cycloneive_lcell_comb \Selector27~4 (
// Equation(s):
// \Selector27~4_combout  = (\Selector27~1_combout ) # ((\Selector24~0_combout  & \Selector27~3_combout ))

	.dataa(\Selector24~0_combout ),
	.datab(gnd),
	.datac(\Selector27~1_combout ),
	.datad(\Selector27~3_combout ),
	.cin(gnd),
	.combout(\Selector27~4_combout ),
	.cout());
// synopsys translate_off
defparam \Selector27~4 .lut_mask = 16'hFAF0;
defparam \Selector27~4 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y42_N12
cycloneive_lcell_comb \Selector24~6 (
// Equation(s):
// \Selector24~6_combout  = (\portb~52_combout  & ((\Selector0~3_combout ) # ((\porta~93_combout  & \Selector0~4_combout ))))

	.dataa(\Selector0~3_combout ),
	.datab(porta9),
	.datac(\Selector0~4_combout ),
	.datad(portb24),
	.cin(gnd),
	.combout(\Selector24~6_combout ),
	.cout());
// synopsys translate_off
defparam \Selector24~6 .lut_mask = 16'hEA00;
defparam \Selector24~6 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y42_N22
cycloneive_lcell_comb \Selector24~7 (
// Equation(s):
// \Selector24~7_combout  = (\porta~93_combout  & (((\Selector0~3_combout )))) # (!\porta~93_combout  & (\Selector0~7_combout  & ((!\portb~52_combout ))))

	.dataa(\Selector0~7_combout ),
	.datab(porta9),
	.datac(\Selector0~3_combout ),
	.datad(portb24),
	.cin(gnd),
	.combout(\Selector24~7_combout ),
	.cout());
// synopsys translate_off
defparam \Selector24~7 .lut_mask = 16'hC0E2;
defparam \Selector24~7 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y42_N28
cycloneive_lcell_comb \Selector24~8 (
// Equation(s):
// \Selector24~8_combout  = (\Selector24~7_combout ) # ((\Selector0~2_combout  & (\porta~93_combout  $ (\portb~52_combout ))))

	.dataa(\Selector24~7_combout ),
	.datab(\Selector0~2_combout ),
	.datac(porta9),
	.datad(portb24),
	.cin(gnd),
	.combout(\Selector24~8_combout ),
	.cout());
// synopsys translate_off
defparam \Selector24~8 .lut_mask = 16'hAEEA;
defparam \Selector24~8 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y40_N12
cycloneive_lcell_comb \Add1~12 (
// Equation(s):
// \Add1~12_combout  = ((\porta~94_combout  $ (\portb~54_combout  $ (\Add1~11 )))) # (GND)
// \Add1~13  = CARRY((\porta~94_combout  & ((!\Add1~11 ) # (!\portb~54_combout ))) # (!\porta~94_combout  & (!\portb~54_combout  & !\Add1~11 )))

	.dataa(porta10),
	.datab(portb25),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add1~11 ),
	.combout(\Add1~12_combout ),
	.cout(\Add1~13 ));
// synopsys translate_off
defparam \Add1~12 .lut_mask = 16'h962B;
defparam \Add1~12 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X57_Y40_N14
cycloneive_lcell_comb \Add1~14 (
// Equation(s):
// \Add1~14_combout  = (\porta~93_combout  & ((\portb~52_combout  & (!\Add1~13 )) # (!\portb~52_combout  & (\Add1~13  & VCC)))) # (!\porta~93_combout  & ((\portb~52_combout  & ((\Add1~13 ) # (GND))) # (!\portb~52_combout  & (!\Add1~13 ))))
// \Add1~15  = CARRY((\porta~93_combout  & (\portb~52_combout  & !\Add1~13 )) # (!\porta~93_combout  & ((\portb~52_combout ) # (!\Add1~13 ))))

	.dataa(porta9),
	.datab(portb24),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add1~13 ),
	.combout(\Add1~14_combout ),
	.cout(\Add1~15 ));
// synopsys translate_off
defparam \Add1~14 .lut_mask = 16'h694D;
defparam \Add1~14 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X53_Y42_N28
cycloneive_lcell_comb \Selector24~2 (
// Equation(s):
// \Selector24~2_combout  = (\Add0~14_combout  & ((\Selector0~5_combout ) # ((\Add1~14_combout  & \Selector0~6_combout )))) # (!\Add0~14_combout  & (\Add1~14_combout  & (\Selector0~6_combout )))

	.dataa(\Add0~14_combout ),
	.datab(\Add1~14_combout ),
	.datac(\Selector0~6_combout ),
	.datad(\Selector0~5_combout ),
	.cin(gnd),
	.combout(\Selector24~2_combout ),
	.cout());
// synopsys translate_off
defparam \Selector24~2 .lut_mask = 16'hEAC0;
defparam \Selector24~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y42_N18
cycloneive_lcell_comb \ShiftRight0~101 (
// Equation(s):
// \ShiftRight0~101_combout  = (\portb~64_combout  & (!\portb~62_combout  & ((\ShiftRight0~78_combout )))) # (!\portb~64_combout  & (\portb~62_combout  & (\ShiftRight0~80_combout )))

	.dataa(portb30),
	.datab(portb29),
	.datac(\ShiftRight0~80_combout ),
	.datad(\ShiftRight0~78_combout ),
	.cin(gnd),
	.combout(\ShiftRight0~101_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftRight0~101 .lut_mask = 16'h6240;
defparam \ShiftRight0~101 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y42_N30
cycloneive_lcell_comb \ShiftRight0~105 (
// Equation(s):
// \ShiftRight0~105_combout  = (\ShiftRight0~101_combout ) # ((!\portb~64_combout  & (!\portb~62_combout  & \ShiftRight0~82_combout )))

	.dataa(portb30),
	.datab(portb29),
	.datac(\ShiftRight0~82_combout ),
	.datad(\ShiftRight0~101_combout ),
	.cin(gnd),
	.combout(\ShiftRight0~105_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftRight0~105 .lut_mask = 16'hFF10;
defparam \ShiftRight0~105 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y42_N12
cycloneive_lcell_comb \Selector24~3 (
// Equation(s):
// \Selector24~3_combout  = (\Selector7~1_combout  & ((\ShiftRight0~76_combout ) # ((\Selector7~0_combout )))) # (!\Selector7~1_combout  & (((!\Selector7~0_combout  & \ShiftRight0~73_combout ))))

	.dataa(\ShiftRight0~76_combout ),
	.datab(\Selector7~1_combout ),
	.datac(\Selector7~0_combout ),
	.datad(\ShiftRight0~73_combout ),
	.cin(gnd),
	.combout(\Selector24~3_combout ),
	.cout());
// synopsys translate_off
defparam \Selector24~3 .lut_mask = 16'hCBC8;
defparam \Selector24~3 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y42_N8
cycloneive_lcell_comb \Selector24~4 (
// Equation(s):
// \Selector24~4_combout  = (\Selector7~0_combout  & ((\Selector24~3_combout  & ((\ShiftRight0~105_combout ))) # (!\Selector24~3_combout  & (\ShiftRight0~100_combout )))) # (!\Selector7~0_combout  & (((\Selector24~3_combout ))))

	.dataa(\ShiftRight0~100_combout ),
	.datab(\Selector7~0_combout ),
	.datac(\ShiftRight0~105_combout ),
	.datad(\Selector24~3_combout ),
	.cin(gnd),
	.combout(\Selector24~4_combout ),
	.cout());
// synopsys translate_off
defparam \Selector24~4 .lut_mask = 16'hF388;
defparam \Selector24~4 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y42_N26
cycloneive_lcell_comb \Selector24~5 (
// Equation(s):
// \Selector24~5_combout  = (\Selector24~2_combout ) # ((\Selector24~0_combout  & \Selector24~4_combout ))

	.dataa(gnd),
	.datab(\Selector24~2_combout ),
	.datac(\Selector24~0_combout ),
	.datad(\Selector24~4_combout ),
	.cin(gnd),
	.combout(\Selector24~5_combout ),
	.cout());
// synopsys translate_off
defparam \Selector24~5 .lut_mask = 16'hFCCC;
defparam \Selector24~5 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y37_N8
cycloneive_lcell_comb \ShiftLeft0~16 (
// Equation(s):
// \ShiftLeft0~16_combout  = (\portb~60_combout  & ((\ShiftLeft0~7_combout ))) # (!\portb~60_combout  & (\ShiftLeft0~15_combout ))

	.dataa(\ShiftLeft0~15_combout ),
	.datab(\ShiftLeft0~7_combout ),
	.datac(gnd),
	.datad(portb28),
	.cin(gnd),
	.combout(\ShiftLeft0~16_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftLeft0~16 .lut_mask = 16'hCCAA;
defparam \ShiftLeft0~16 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X52_Y36_N14
cycloneive_lcell_comb \ShiftLeft0~17 (
// Equation(s):
// \ShiftLeft0~17_combout  = (\portb~62_combout  & ((\ShiftLeft0~4_combout ))) # (!\portb~62_combout  & (\ShiftLeft0~16_combout ))

	.dataa(portb29),
	.datab(\ShiftLeft0~16_combout ),
	.datac(\ShiftLeft0~4_combout ),
	.datad(gnd),
	.cin(gnd),
	.combout(\ShiftLeft0~17_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftLeft0~17 .lut_mask = 16'hE4E4;
defparam \ShiftLeft0~17 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y42_N2
cycloneive_lcell_comb \Selector24~1 (
// Equation(s):
// \Selector24~1_combout  = (!\portb~64_combout  & (\Selector0~1_combout  & (!\Selector1~1_combout  & \ShiftLeft0~17_combout )))

	.dataa(portb30),
	.datab(\Selector0~1_combout ),
	.datac(\Selector1~1_combout ),
	.datad(\ShiftLeft0~17_combout ),
	.cin(gnd),
	.combout(\Selector24~1_combout ),
	.cout());
// synopsys translate_off
defparam \Selector24~1 .lut_mask = 16'h0400;
defparam \Selector24~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y38_N26
cycloneive_lcell_comb \Selector24~10 (
// Equation(s):
// \Selector24~10_combout  = (!\ShiftRight0~72_combout  & (!\portb~66_combout  & (\Selector0~1_combout  & !\portb~64_combout )))

	.dataa(\ShiftRight0~72_combout ),
	.datab(portb31),
	.datac(\Selector0~1_combout ),
	.datad(portb30),
	.cin(gnd),
	.combout(\Selector24~10_combout ),
	.cout());
// synopsys translate_off
defparam \Selector24~10 .lut_mask = 16'h0010;
defparam \Selector24~10 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y41_N20
cycloneive_lcell_comb \ShiftLeft0~18 (
// Equation(s):
// \ShiftLeft0~18_combout  = (\portb~58_combout  & (\porta~95_combout )) # (!\portb~58_combout  & ((\porta~94_combout )))

	.dataa(gnd),
	.datab(portb27),
	.datac(porta11),
	.datad(porta10),
	.cin(gnd),
	.combout(\ShiftLeft0~18_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftLeft0~18 .lut_mask = 16'hF3C0;
defparam \ShiftLeft0~18 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y41_N22
cycloneive_lcell_comb \ShiftLeft0~19 (
// Equation(s):
// \ShiftLeft0~19_combout  = (\portb~60_combout  & ((\ShiftLeft0~12_combout ))) # (!\portb~60_combout  & (\ShiftLeft0~18_combout ))

	.dataa(gnd),
	.datab(\ShiftLeft0~18_combout ),
	.datac(portb28),
	.datad(\ShiftLeft0~12_combout ),
	.cin(gnd),
	.combout(\ShiftLeft0~19_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftLeft0~19 .lut_mask = 16'hFC0C;
defparam \ShiftLeft0~19 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y41_N8
cycloneive_lcell_comb \ShiftLeft0~20 (
// Equation(s):
// \ShiftLeft0~20_combout  = (\portb~62_combout  & ((\ShiftLeft0~6_combout ))) # (!\portb~62_combout  & (\ShiftLeft0~19_combout ))

	.dataa(portb29),
	.datab(gnd),
	.datac(\ShiftLeft0~19_combout ),
	.datad(\ShiftLeft0~6_combout ),
	.cin(gnd),
	.combout(\ShiftLeft0~20_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftLeft0~20 .lut_mask = 16'hFA50;
defparam \ShiftLeft0~20 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y42_N8
cycloneive_lcell_comb \Selector25~5 (
// Equation(s):
// \Selector25~5_combout  = (\porta~94_combout  & ((\Selector0~3_combout ) # (!\portb~54_combout ))) # (!\porta~94_combout  & ((\portb~54_combout )))

	.dataa(\Selector0~3_combout ),
	.datab(gnd),
	.datac(porta10),
	.datad(portb25),
	.cin(gnd),
	.combout(\Selector25~5_combout ),
	.cout());
// synopsys translate_off
defparam \Selector25~5 .lut_mask = 16'hAFF0;
defparam \Selector25~5 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y42_N18
cycloneive_lcell_comb \Selector25~4 (
// Equation(s):
// \Selector25~4_combout  = (\porta~94_combout  & (\Selector0~4_combout )) # (!\porta~94_combout  & ((\Selector0~7_combout )))

	.dataa(porta10),
	.datab(gnd),
	.datac(\Selector0~4_combout ),
	.datad(\Selector0~7_combout ),
	.cin(gnd),
	.combout(\Selector25~4_combout ),
	.cout());
// synopsys translate_off
defparam \Selector25~4 .lut_mask = 16'hF5A0;
defparam \Selector25~4 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y42_N2
cycloneive_lcell_comb \Selector25~6 (
// Equation(s):
// \Selector25~6_combout  = (\Selector25~5_combout  & ((\Selector0~2_combout ) # ((\Selector0~3_combout )))) # (!\Selector25~5_combout  & (((\Selector25~4_combout ))))

	.dataa(\Selector0~2_combout ),
	.datab(\Selector25~5_combout ),
	.datac(\Selector0~3_combout ),
	.datad(\Selector25~4_combout ),
	.cin(gnd),
	.combout(\Selector25~6_combout ),
	.cout());
// synopsys translate_off
defparam \Selector25~6 .lut_mask = 16'hFBC8;
defparam \Selector25~6 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X52_Y38_N12
cycloneive_lcell_comb \Add0~12 (
// Equation(s):
// \Add0~12_combout  = ((\porta~94_combout  $ (\portb~54_combout  $ (!\Add0~11 )))) # (GND)
// \Add0~13  = CARRY((\porta~94_combout  & ((\portb~54_combout ) # (!\Add0~11 ))) # (!\porta~94_combout  & (\portb~54_combout  & !\Add0~11 )))

	.dataa(porta10),
	.datab(portb25),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add0~11 ),
	.combout(\Add0~12_combout ),
	.cout(\Add0~13 ));
// synopsys translate_off
defparam \Add0~12 .lut_mask = 16'h698E;
defparam \Add0~12 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X55_Y39_N4
cycloneive_lcell_comb \Selector25~0 (
// Equation(s):
// \Selector25~0_combout  = (\Selector0~6_combout  & ((\Add1~12_combout ) # ((\Selector0~5_combout  & \Add0~12_combout )))) # (!\Selector0~6_combout  & (\Selector0~5_combout  & (\Add0~12_combout )))

	.dataa(\Selector0~6_combout ),
	.datab(\Selector0~5_combout ),
	.datac(\Add0~12_combout ),
	.datad(\Add1~12_combout ),
	.cin(gnd),
	.combout(\Selector25~0_combout ),
	.cout());
// synopsys translate_off
defparam \Selector25~0 .lut_mask = 16'hEAC0;
defparam \Selector25~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y39_N22
cycloneive_lcell_comb \ShiftRight0~103 (
// Equation(s):
// \ShiftRight0~103_combout  = (\portb~64_combout  & (!\portb~60_combout  & (!\portb~62_combout  & \ShiftRight0~57_combout )))

	.dataa(portb30),
	.datab(portb28),
	.datac(portb29),
	.datad(\ShiftRight0~57_combout ),
	.cin(gnd),
	.combout(\ShiftRight0~103_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftRight0~103 .lut_mask = 16'h0200;
defparam \ShiftRight0~103 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y39_N8
cycloneive_lcell_comb \ShiftRight0~104 (
// Equation(s):
// \ShiftRight0~104_combout  = (\ShiftRight0~103_combout ) # ((!\portb~64_combout  & (\portb~62_combout  & \ShiftRight0~89_combout )))

	.dataa(portb30),
	.datab(\ShiftRight0~103_combout ),
	.datac(portb29),
	.datad(\ShiftRight0~89_combout ),
	.cin(gnd),
	.combout(\ShiftRight0~104_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftRight0~104 .lut_mask = 16'hDCCC;
defparam \ShiftRight0~104 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y39_N30
cycloneive_lcell_comb \ShiftRight0~106 (
// Equation(s):
// \ShiftRight0~106_combout  = (\ShiftRight0~104_combout ) # ((!\portb~64_combout  & (!\portb~62_combout  & \ShiftRight0~91_combout )))

	.dataa(portb30),
	.datab(\ShiftRight0~104_combout ),
	.datac(portb29),
	.datad(\ShiftRight0~91_combout ),
	.cin(gnd),
	.combout(\ShiftRight0~106_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftRight0~106 .lut_mask = 16'hCDCC;
defparam \ShiftRight0~106 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X52_Y41_N20
cycloneive_lcell_comb \ShiftRight0~85 (
// Equation(s):
// \ShiftRight0~85_combout  = (\portb~60_combout  & ((\ShiftRight0~53_combout ))) # (!\portb~60_combout  & (\ShiftRight0~45_combout ))

	.dataa(gnd),
	.datab(\ShiftRight0~45_combout ),
	.datac(portb28),
	.datad(\ShiftRight0~53_combout ),
	.cin(gnd),
	.combout(\ShiftRight0~85_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftRight0~85 .lut_mask = 16'hFC0C;
defparam \ShiftRight0~85 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y36_N30
cycloneive_lcell_comb \ShiftRight0~102 (
// Equation(s):
// \ShiftRight0~102_combout  = (\portb~62_combout  & (\ShiftRight0~92_combout )) # (!\portb~62_combout  & ((\ShiftRight0~86_combout )))

	.dataa(gnd),
	.datab(\ShiftRight0~92_combout ),
	.datac(portb29),
	.datad(\ShiftRight0~86_combout ),
	.cin(gnd),
	.combout(\ShiftRight0~102_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftRight0~102 .lut_mask = 16'hCFC0;
defparam \ShiftRight0~102 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X52_Y41_N10
cycloneive_lcell_comb \Selector25~1 (
// Equation(s):
// \Selector25~1_combout  = (\Selector7~1_combout  & (((\Selector7~0_combout )))) # (!\Selector7~1_combout  & ((\Selector7~0_combout  & ((\ShiftRight0~102_combout ))) # (!\Selector7~0_combout  & (\ShiftRight0~85_combout ))))

	.dataa(\Selector7~1_combout ),
	.datab(\ShiftRight0~85_combout ),
	.datac(\Selector7~0_combout ),
	.datad(\ShiftRight0~102_combout ),
	.cin(gnd),
	.combout(\Selector25~1_combout ),
	.cout());
// synopsys translate_off
defparam \Selector25~1 .lut_mask = 16'hF4A4;
defparam \Selector25~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y39_N6
cycloneive_lcell_comb \Selector25~2 (
// Equation(s):
// \Selector25~2_combout  = (\Selector7~1_combout  & ((\Selector25~1_combout  & ((\ShiftRight0~106_combout ))) # (!\Selector25~1_combout  & (\ShiftRight0~87_combout )))) # (!\Selector7~1_combout  & (((\Selector25~1_combout ))))

	.dataa(\ShiftRight0~87_combout ),
	.datab(\Selector7~1_combout ),
	.datac(\ShiftRight0~106_combout ),
	.datad(\Selector25~1_combout ),
	.cin(gnd),
	.combout(\Selector25~2_combout ),
	.cout());
// synopsys translate_off
defparam \Selector25~2 .lut_mask = 16'hF388;
defparam \Selector25~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y39_N16
cycloneive_lcell_comb \Selector25~3 (
// Equation(s):
// \Selector25~3_combout  = (\Selector25~0_combout ) # ((\Selector24~0_combout  & \Selector25~2_combout ))

	.dataa(gnd),
	.datab(\Selector24~0_combout ),
	.datac(\Selector25~0_combout ),
	.datad(\Selector25~2_combout ),
	.cin(gnd),
	.combout(\Selector25~3_combout ),
	.cout());
// synopsys translate_off
defparam \Selector25~3 .lut_mask = 16'hFCF0;
defparam \Selector25~3 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X52_Y38_N16
cycloneive_lcell_comb \Add0~16 (
// Equation(s):
// \Add0~16_combout  = ((\porta~92_combout  $ (\portb~50_combout  $ (!\Add0~15 )))) # (GND)
// \Add0~17  = CARRY((\porta~92_combout  & ((\portb~50_combout ) # (!\Add0~15 ))) # (!\porta~92_combout  & (\portb~50_combout  & !\Add0~15 )))

	.dataa(porta8),
	.datab(portb23),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add0~15 ),
	.combout(\Add0~16_combout ),
	.cout(\Add0~17 ));
// synopsys translate_off
defparam \Add0~16 .lut_mask = 16'h698E;
defparam \Add0~16 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X52_Y38_N18
cycloneive_lcell_comb \Add0~18 (
// Equation(s):
// \Add0~18_combout  = (\porta~103_combout  & ((\portb~48_combout  & (\Add0~17  & VCC)) # (!\portb~48_combout  & (!\Add0~17 )))) # (!\porta~103_combout  & ((\portb~48_combout  & (!\Add0~17 )) # (!\portb~48_combout  & ((\Add0~17 ) # (GND)))))
// \Add0~19  = CARRY((\porta~103_combout  & (!\portb~48_combout  & !\Add0~17 )) # (!\porta~103_combout  & ((!\Add0~17 ) # (!\portb~48_combout ))))

	.dataa(porta19),
	.datab(portb22),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add0~17 ),
	.combout(\Add0~18_combout ),
	.cout(\Add0~19 ));
// synopsys translate_off
defparam \Add0~18 .lut_mask = 16'h9617;
defparam \Add0~18 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X54_Y38_N2
cycloneive_lcell_comb \Selector1~2 (
// Equation(s):
// \Selector1~2_combout  = (plif_idexaluop_l_3) # ((!\ShiftRight0~72_combout  & ((\portb~64_combout ) # (\portb~66_combout ))))

	.dataa(plif_idexaluop_l_3),
	.datab(portb30),
	.datac(portb31),
	.datad(\ShiftRight0~72_combout ),
	.cin(gnd),
	.combout(\Selector1~2_combout ),
	.cout());
// synopsys translate_off
defparam \Selector1~2 .lut_mask = 16'hAAFE;
defparam \Selector1~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y38_N8
cycloneive_lcell_comb \Selector16~1 (
// Equation(s):
// \Selector16~1_combout  = (plif_idexaluop_l_0 & (\Selector0~15_combout  & !\Selector1~2_combout ))

	.dataa(gnd),
	.datab(plif_idexaluop_l_0),
	.datac(\Selector0~15_combout ),
	.datad(\Selector1~2_combout ),
	.cin(gnd),
	.combout(\Selector16~1_combout ),
	.cout());
// synopsys translate_off
defparam \Selector16~1 .lut_mask = 16'h00C0;
defparam \Selector16~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y38_N18
cycloneive_lcell_comb \Selector1~3 (
// Equation(s):
// \Selector1~3_combout  = (!plif_idexaluop_l_1 & (!plif_idexaluop_l_2 & (!plif_idexaluop_l_3 & !\ShiftRight0~72_combout )))

	.dataa(plif_idexaluop_l_1),
	.datab(plif_idexaluop_l_2),
	.datac(plif_idexaluop_l_3),
	.datad(\ShiftRight0~72_combout ),
	.cin(gnd),
	.combout(\Selector1~3_combout ),
	.cout());
// synopsys translate_off
defparam \Selector1~3 .lut_mask = 16'h0001;
defparam \Selector1~3 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y37_N20
cycloneive_lcell_comb \Selector20~1 (
// Equation(s):
// \Selector20~1_combout  = (plif_idexaluop_l_0 & (!\portb~64_combout  & (\portb~66_combout  & \Selector1~3_combout )))

	.dataa(plif_idexaluop_l_0),
	.datab(portb30),
	.datac(portb31),
	.datad(\Selector1~3_combout ),
	.cin(gnd),
	.combout(\Selector20~1_combout ),
	.cout());
// synopsys translate_off
defparam \Selector20~1 .lut_mask = 16'h2000;
defparam \Selector20~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y41_N4
cycloneive_lcell_comb \Selector22~1 (
// Equation(s):
// \Selector22~1_combout  = (\Selector16~1_combout  & ((\ShiftRight0~25_combout ) # ((\ShiftRight0~32_combout  & \Selector20~1_combout )))) # (!\Selector16~1_combout  & (\ShiftRight0~32_combout  & (\Selector20~1_combout )))

	.dataa(\Selector16~1_combout ),
	.datab(\ShiftRight0~32_combout ),
	.datac(\Selector20~1_combout ),
	.datad(\ShiftRight0~25_combout ),
	.cin(gnd),
	.combout(\Selector22~1_combout ),
	.cout());
// synopsys translate_off
defparam \Selector22~1 .lut_mask = 16'hEAC0;
defparam \Selector22~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y40_N16
cycloneive_lcell_comb \Add1~16 (
// Equation(s):
// \Add1~16_combout  = ((\porta~92_combout  $ (\portb~50_combout  $ (\Add1~15 )))) # (GND)
// \Add1~17  = CARRY((\porta~92_combout  & ((!\Add1~15 ) # (!\portb~50_combout ))) # (!\porta~92_combout  & (!\portb~50_combout  & !\Add1~15 )))

	.dataa(porta8),
	.datab(portb23),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add1~15 ),
	.combout(\Add1~16_combout ),
	.cout(\Add1~17 ));
// synopsys translate_off
defparam \Add1~16 .lut_mask = 16'h962B;
defparam \Add1~16 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X57_Y40_N18
cycloneive_lcell_comb \Add1~18 (
// Equation(s):
// \Add1~18_combout  = (\porta~103_combout  & ((\portb~48_combout  & (!\Add1~17 )) # (!\portb~48_combout  & (\Add1~17  & VCC)))) # (!\porta~103_combout  & ((\portb~48_combout  & ((\Add1~17 ) # (GND))) # (!\portb~48_combout  & (!\Add1~17 ))))
// \Add1~19  = CARRY((\porta~103_combout  & (\portb~48_combout  & !\Add1~17 )) # (!\porta~103_combout  & ((\portb~48_combout ) # (!\Add1~17 ))))

	.dataa(porta19),
	.datab(portb22),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add1~17 ),
	.combout(\Add1~18_combout ),
	.cout(\Add1~19 ));
// synopsys translate_off
defparam \Add1~18 .lut_mask = 16'h694D;
defparam \Add1~18 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X50_Y35_N10
cycloneive_lcell_comb \Selector0~8 (
// Equation(s):
// \Selector0~8_combout  = (!plif_idexaluop_l_2 & (!plif_idexaluop_l_3 & (plif_idexaluop_l_1 & plif_idexaluop_l_0)))

	.dataa(plif_idexaluop_l_2),
	.datab(plif_idexaluop_l_3),
	.datac(plif_idexaluop_l_1),
	.datad(plif_idexaluop_l_0),
	.cin(gnd),
	.combout(\Selector0~8_combout ),
	.cout());
// synopsys translate_off
defparam \Selector0~8 .lut_mask = 16'h1000;
defparam \Selector0~8 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X50_Y38_N14
cycloneive_lcell_comb \ShiftLeft0~22 (
// Equation(s):
// \ShiftLeft0~22_combout  = (!\portb~64_combout  & (\ShiftLeft0~8_combout  & \portb~62_combout ))

	.dataa(portb30),
	.datab(gnd),
	.datac(\ShiftLeft0~8_combout ),
	.datad(portb29),
	.cin(gnd),
	.combout(\ShiftLeft0~22_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftLeft0~22 .lut_mask = 16'h5000;
defparam \ShiftLeft0~22 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X50_Y38_N24
cycloneive_lcell_comb \ShiftLeft0~21 (
// Equation(s):
// \ShiftLeft0~21_combout  = (!\portb~62_combout  & (\portb~64_combout  & (!\portb~60_combout  & \ShiftLeft0~2_combout )))

	.dataa(portb29),
	.datab(portb30),
	.datac(portb28),
	.datad(\ShiftLeft0~2_combout ),
	.cin(gnd),
	.combout(\ShiftLeft0~21_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftLeft0~21 .lut_mask = 16'h0400;
defparam \ShiftLeft0~21 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X50_Y38_N12
cycloneive_lcell_comb \ShiftLeft0~25 (
// Equation(s):
// \ShiftLeft0~25_combout  = (\ShiftLeft0~22_combout ) # ((\ShiftLeft0~21_combout ) # ((\ShiftLeft0~24_combout  & \ShiftRight0~74_combout )))

	.dataa(\ShiftLeft0~24_combout ),
	.datab(\ShiftRight0~74_combout ),
	.datac(\ShiftLeft0~22_combout ),
	.datad(\ShiftLeft0~21_combout ),
	.cin(gnd),
	.combout(\ShiftLeft0~25_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftLeft0~25 .lut_mask = 16'hFFF8;
defparam \ShiftLeft0~25 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X50_Y38_N10
cycloneive_lcell_comb \Selector22~2 (
// Equation(s):
// \Selector22~2_combout  = (\Selector0~14_combout  & (!\portb~66_combout  & (!\ShiftRight0~72_combout  & \ShiftLeft0~25_combout )))

	.dataa(\Selector0~14_combout ),
	.datab(portb31),
	.datac(\ShiftRight0~72_combout ),
	.datad(\ShiftLeft0~25_combout ),
	.cin(gnd),
	.combout(\Selector22~2_combout ),
	.cout());
// synopsys translate_off
defparam \Selector22~2 .lut_mask = 16'h0200;
defparam \Selector22~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y41_N24
cycloneive_lcell_comb \Selector22~4 (
// Equation(s):
// \Selector22~4_combout  = (\porta~103_combout  & (((\Selector0~10_combout )))) # (!\porta~103_combout  & (\Selector0~12_combout  & ((!\portb~48_combout ))))

	.dataa(\Selector0~12_combout ),
	.datab(\Selector0~10_combout ),
	.datac(portb22),
	.datad(porta19),
	.cin(gnd),
	.combout(\Selector22~4_combout ),
	.cout());
// synopsys translate_off
defparam \Selector22~4 .lut_mask = 16'hCC0A;
defparam \Selector22~4 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y41_N2
cycloneive_lcell_comb \Selector22~5 (
// Equation(s):
// \Selector22~5_combout  = (\Selector22~4_combout ) # ((\Selector0~13_combout  & (\portb~48_combout  $ (\porta~103_combout ))))

	.dataa(portb22),
	.datab(porta19),
	.datac(\Selector0~13_combout ),
	.datad(\Selector22~4_combout ),
	.cin(gnd),
	.combout(\Selector22~5_combout ),
	.cout());
// synopsys translate_off
defparam \Selector22~5 .lut_mask = 16'hFF60;
defparam \Selector22~5 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y41_N14
cycloneive_lcell_comb \Selector22~3 (
// Equation(s):
// \Selector22~3_combout  = (\portb~48_combout  & ((\Selector0~10_combout ) # ((\Selector0~11_combout  & \porta~103_combout ))))

	.dataa(\Selector0~11_combout ),
	.datab(\Selector0~10_combout ),
	.datac(portb22),
	.datad(porta19),
	.cin(gnd),
	.combout(\Selector22~3_combout ),
	.cout());
// synopsys translate_off
defparam \Selector22~3 .lut_mask = 16'hE0C0;
defparam \Selector22~3 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y41_N28
cycloneive_lcell_comb \Selector22~6 (
// Equation(s):
// \Selector22~6_combout  = (\Selector22~5_combout ) # ((\Selector22~3_combout ) # ((\Selector0~17_combout  & \Selector22~0_combout )))

	.dataa(\Selector0~17_combout ),
	.datab(\Selector22~5_combout ),
	.datac(\Selector22~3_combout ),
	.datad(\Selector22~0_combout ),
	.cin(gnd),
	.combout(\Selector22~6_combout ),
	.cout());
// synopsys translate_off
defparam \Selector22~6 .lut_mask = 16'hFEFC;
defparam \Selector22~6 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y41_N10
cycloneive_lcell_comb \Selector22~7 (
// Equation(s):
// \Selector22~7_combout  = (\Selector22~2_combout ) # ((\Selector22~6_combout ) # ((\Add1~18_combout  & \Selector0~8_combout )))

	.dataa(\Add1~18_combout ),
	.datab(\Selector0~8_combout ),
	.datac(\Selector22~2_combout ),
	.datad(\Selector22~6_combout ),
	.cin(gnd),
	.combout(\Selector22~7_combout ),
	.cout());
// synopsys translate_off
defparam \Selector22~7 .lut_mask = 16'hFFF8;
defparam \Selector22~7 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y41_N14
cycloneive_lcell_comb \ShiftLeft0~27 (
// Equation(s):
// \ShiftLeft0~27_combout  = (\portb~58_combout  & ((\porta~93_combout ))) # (!\portb~58_combout  & (\porta~92_combout ))

	.dataa(gnd),
	.datab(portb27),
	.datac(porta8),
	.datad(porta9),
	.cin(gnd),
	.combout(\ShiftLeft0~27_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftLeft0~27 .lut_mask = 16'hFC30;
defparam \ShiftLeft0~27 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y41_N30
cycloneive_lcell_comb \ShiftLeft0~28 (
// Equation(s):
// \ShiftLeft0~28_combout  = (\portb~60_combout  & (\ShiftLeft0~18_combout )) # (!\portb~60_combout  & ((\ShiftLeft0~27_combout )))

	.dataa(\ShiftLeft0~18_combout ),
	.datab(gnd),
	.datac(\ShiftLeft0~27_combout ),
	.datad(portb28),
	.cin(gnd),
	.combout(\ShiftLeft0~28_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftLeft0~28 .lut_mask = 16'hAAF0;
defparam \ShiftLeft0~28 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y40_N0
cycloneive_lcell_comb \ShiftLeft0~26 (
// Equation(s):
// \ShiftLeft0~26_combout  = (\portb~64_combout  & (!\portb~62_combout  & (\ShiftLeft0~10_combout ))) # (!\portb~64_combout  & (\portb~62_combout  & ((\ShiftLeft0~13_combout ))))

	.dataa(portb30),
	.datab(portb29),
	.datac(\ShiftLeft0~10_combout ),
	.datad(\ShiftLeft0~13_combout ),
	.cin(gnd),
	.combout(\ShiftLeft0~26_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftLeft0~26 .lut_mask = 16'h6420;
defparam \ShiftLeft0~26 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y40_N22
cycloneive_lcell_comb \ShiftLeft0~80 (
// Equation(s):
// \ShiftLeft0~80_combout  = (\ShiftLeft0~26_combout ) # ((!\portb~64_combout  & (\ShiftLeft0~28_combout  & !\portb~62_combout )))

	.dataa(portb30),
	.datab(\ShiftLeft0~28_combout ),
	.datac(portb29),
	.datad(\ShiftLeft0~26_combout ),
	.cin(gnd),
	.combout(\ShiftLeft0~80_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftLeft0~80 .lut_mask = 16'hFF04;
defparam \ShiftLeft0~80 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y40_N8
cycloneive_lcell_comb \Selector23~6 (
// Equation(s):
// \Selector23~6_combout  = (\Selector0~8_combout  & \Add1~16_combout )

	.dataa(\Selector0~8_combout ),
	.datab(gnd),
	.datac(gnd),
	.datad(\Add1~16_combout ),
	.cin(gnd),
	.combout(\Selector23~6_combout ),
	.cout());
// synopsys translate_off
defparam \Selector23~6 .lut_mask = 16'hAA00;
defparam \Selector23~6 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X50_Y40_N4
cycloneive_lcell_comb \Selector23~2 (
// Equation(s):
// \Selector23~2_combout  = (\portb~50_combout  & ((\porta~92_combout  & ((\Selector0~11_combout ))) # (!\porta~92_combout  & (\Selector0~13_combout )))) # (!\portb~50_combout  & ((\Selector0~13_combout ) # ((!\porta~92_combout ))))

	.dataa(portb23),
	.datab(\Selector0~13_combout ),
	.datac(\Selector0~11_combout ),
	.datad(porta8),
	.cin(gnd),
	.combout(\Selector23~2_combout ),
	.cout());
// synopsys translate_off
defparam \Selector23~2 .lut_mask = 16'hE4DD;
defparam \Selector23~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X50_Y40_N2
cycloneive_lcell_comb \Selector23~3 (
// Equation(s):
// \Selector23~3_combout  = (\porta~92_combout ) # ((\Selector0~12_combout ) # (\portb~50_combout ))

	.dataa(porta8),
	.datab(gnd),
	.datac(\Selector0~12_combout ),
	.datad(portb23),
	.cin(gnd),
	.combout(\Selector23~3_combout ),
	.cout());
// synopsys translate_off
defparam \Selector23~3 .lut_mask = 16'hFFFA;
defparam \Selector23~3 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X50_Y40_N20
cycloneive_lcell_comb \Selector23~4 (
// Equation(s):
// \Selector23~4_combout  = (\Selector23~3_combout  & ((\Selector0~10_combout ) # (\Selector23~2_combout )))

	.dataa(gnd),
	.datab(\Selector0~10_combout ),
	.datac(\Selector23~2_combout ),
	.datad(\Selector23~3_combout ),
	.cin(gnd),
	.combout(\Selector23~4_combout ),
	.cout());
// synopsys translate_off
defparam \Selector23~4 .lut_mask = 16'hFC00;
defparam \Selector23~4 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y40_N10
cycloneive_lcell_comb \Selector23~5 (
// Equation(s):
// \Selector23~5_combout  = (\Selector23~4_combout ) # ((!\portb~64_combout  & (\Selector23~1_combout  & \ShiftRight0~63_combout )))

	.dataa(portb30),
	.datab(\Selector23~1_combout ),
	.datac(\Selector23~4_combout ),
	.datad(\ShiftRight0~63_combout ),
	.cin(gnd),
	.combout(\Selector23~5_combout ),
	.cout());
// synopsys translate_off
defparam \Selector23~5 .lut_mask = 16'hF4F0;
defparam \Selector23~5 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y40_N14
cycloneive_lcell_comb \Selector23~7 (
// Equation(s):
// \Selector23~7_combout  = (\Selector23~6_combout ) # ((\Selector23~5_combout ) # ((\Selector0~9_combout  & \Add0~16_combout )))

	.dataa(\Selector0~9_combout ),
	.datab(\Selector23~6_combout ),
	.datac(\Add0~16_combout ),
	.datad(\Selector23~5_combout ),
	.cin(gnd),
	.combout(\Selector23~7_combout ),
	.cout());
// synopsys translate_off
defparam \Selector23~7 .lut_mask = 16'hFFEC;
defparam \Selector23~7 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y42_N22
cycloneive_lcell_comb \Selector0~16 (
// Equation(s):
// \Selector0~16_combout  = (!\portb~66_combout  & \portb~64_combout )

	.dataa(gnd),
	.datab(gnd),
	.datac(portb31),
	.datad(portb30),
	.cin(gnd),
	.combout(\Selector0~16_combout ),
	.cout());
// synopsys translate_off
defparam \Selector0~16 .lut_mask = 16'h0F00;
defparam \Selector0~16 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y38_N16
cycloneive_lcell_comb \Selector0~17 (
// Equation(s):
// \Selector0~17_combout  = (!plif_idexaluop_l_3 & (plif_idexaluop_l_0 & (\Selector0~16_combout  & \Selector0~15_combout )))

	.dataa(plif_idexaluop_l_3),
	.datab(plif_idexaluop_l_0),
	.datac(\Selector0~16_combout ),
	.datad(\Selector0~15_combout ),
	.cin(gnd),
	.combout(\Selector0~17_combout ),
	.cout());
// synopsys translate_off
defparam \Selector0~17 .lut_mask = 16'h4000;
defparam \Selector0~17 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y40_N24
cycloneive_lcell_comb \Selector23~8 (
// Equation(s):
// \Selector23~8_combout  = (\Selector0~17_combout  & ((\Selector23~0_combout ) # ((\Selector16~1_combout  & \ShiftRight0~55_combout )))) # (!\Selector0~17_combout  & (\Selector16~1_combout  & (\ShiftRight0~55_combout )))

	.dataa(\Selector0~17_combout ),
	.datab(\Selector16~1_combout ),
	.datac(\ShiftRight0~55_combout ),
	.datad(\Selector23~0_combout ),
	.cin(gnd),
	.combout(\Selector23~8_combout ),
	.cout());
// synopsys translate_off
defparam \Selector23~8 .lut_mask = 16'hEAC0;
defparam \Selector23~8 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X52_Y41_N12
cycloneive_lcell_comb \ShiftLeft0~23 (
// Equation(s):
// \ShiftLeft0~23_combout  = (\portb~58_combout  & ((\porta~92_combout ))) # (!\portb~58_combout  & (\porta~103_combout ))

	.dataa(portb27),
	.datab(gnd),
	.datac(porta19),
	.datad(porta8),
	.cin(gnd),
	.combout(\ShiftLeft0~23_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftLeft0~23 .lut_mask = 16'hFA50;
defparam \ShiftLeft0~23 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y34_N22
cycloneive_lcell_comb \ShiftLeft0~29 (
// Equation(s):
// \ShiftLeft0~29_combout  = (\portb~58_combout  & (\porta~102_combout )) # (!\portb~58_combout  & ((\porta~101_combout )))

	.dataa(gnd),
	.datab(porta18),
	.datac(portb27),
	.datad(porta17),
	.cin(gnd),
	.combout(\ShiftLeft0~29_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftLeft0~29 .lut_mask = 16'hCFC0;
defparam \ShiftLeft0~29 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y37_N10
cycloneive_lcell_comb \ShiftLeft0~30 (
// Equation(s):
// \ShiftLeft0~30_combout  = (\portb~60_combout  & (\ShiftLeft0~23_combout )) # (!\portb~60_combout  & ((\ShiftLeft0~29_combout )))

	.dataa(portb28),
	.datab(gnd),
	.datac(\ShiftLeft0~23_combout ),
	.datad(\ShiftLeft0~29_combout ),
	.cin(gnd),
	.combout(\ShiftLeft0~30_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftLeft0~30 .lut_mask = 16'hF5A0;
defparam \ShiftLeft0~30 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y37_N20
cycloneive_lcell_comb \ShiftLeft0~31 (
// Equation(s):
// \ShiftLeft0~31_combout  = (!\portb~64_combout  & ((\portb~62_combout  & (\ShiftLeft0~16_combout )) # (!\portb~62_combout  & ((\ShiftLeft0~30_combout )))))

	.dataa(portb29),
	.datab(\ShiftLeft0~16_combout ),
	.datac(portb30),
	.datad(\ShiftLeft0~30_combout ),
	.cin(gnd),
	.combout(\ShiftLeft0~31_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftLeft0~31 .lut_mask = 16'h0D08;
defparam \ShiftLeft0~31 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y36_N24
cycloneive_lcell_comb \ShiftLeft0~32 (
// Equation(s):
// \ShiftLeft0~32_combout  = (\ShiftLeft0~31_combout ) # ((\portb~64_combout  & (!\portb~62_combout  & \ShiftLeft0~4_combout )))

	.dataa(portb30),
	.datab(portb29),
	.datac(\ShiftLeft0~4_combout ),
	.datad(\ShiftLeft0~31_combout ),
	.cin(gnd),
	.combout(\ShiftLeft0~32_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftLeft0~32 .lut_mask = 16'hFF20;
defparam \ShiftLeft0~32 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y37_N26
cycloneive_lcell_comb \Selector20~8 (
// Equation(s):
// \Selector20~8_combout  = (\Selector20~0_combout  & ((\Selector0~17_combout ) # ((\Selector20~1_combout  & \ShiftRight0~81_combout )))) # (!\Selector20~0_combout  & (\Selector20~1_combout  & ((\ShiftRight0~81_combout ))))

	.dataa(\Selector20~0_combout ),
	.datab(\Selector20~1_combout ),
	.datac(\Selector0~17_combout ),
	.datad(\ShiftRight0~81_combout ),
	.cin(gnd),
	.combout(\Selector20~8_combout ),
	.cout());
// synopsys translate_off
defparam \Selector20~8 .lut_mask = 16'hECA0;
defparam \Selector20~8 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y40_N20
cycloneive_lcell_comb \Add1~20 (
// Equation(s):
// \Add1~20_combout  = ((\porta~102_combout  $ (\portb~46_combout  $ (\Add1~19 )))) # (GND)
// \Add1~21  = CARRY((\porta~102_combout  & ((!\Add1~19 ) # (!\portb~46_combout ))) # (!\porta~102_combout  & (!\portb~46_combout  & !\Add1~19 )))

	.dataa(porta18),
	.datab(portb21),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add1~19 ),
	.combout(\Add1~20_combout ),
	.cout(\Add1~21 ));
// synopsys translate_off
defparam \Add1~20 .lut_mask = 16'h962B;
defparam \Add1~20 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X57_Y40_N22
cycloneive_lcell_comb \Add1~22 (
// Equation(s):
// \Add1~22_combout  = (\porta~101_combout  & ((\portb~44_combout  & (!\Add1~21 )) # (!\portb~44_combout  & (\Add1~21  & VCC)))) # (!\porta~101_combout  & ((\portb~44_combout  & ((\Add1~21 ) # (GND))) # (!\portb~44_combout  & (!\Add1~21 ))))
// \Add1~23  = CARRY((\porta~101_combout  & (\portb~44_combout  & !\Add1~21 )) # (!\porta~101_combout  & ((\portb~44_combout ) # (!\Add1~21 ))))

	.dataa(porta17),
	.datab(portb20),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add1~21 ),
	.combout(\Add1~22_combout ),
	.cout(\Add1~23 ));
// synopsys translate_off
defparam \Add1~22 .lut_mask = 16'h694D;
defparam \Add1~22 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X52_Y38_N20
cycloneive_lcell_comb \Add0~20 (
// Equation(s):
// \Add0~20_combout  = ((\portb~46_combout  $ (\porta~102_combout  $ (!\Add0~19 )))) # (GND)
// \Add0~21  = CARRY((\portb~46_combout  & ((\porta~102_combout ) # (!\Add0~19 ))) # (!\portb~46_combout  & (\porta~102_combout  & !\Add0~19 )))

	.dataa(portb21),
	.datab(porta18),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add0~19 ),
	.combout(\Add0~20_combout ),
	.cout(\Add0~21 ));
// synopsys translate_off
defparam \Add0~20 .lut_mask = 16'h698E;
defparam \Add0~20 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X52_Y38_N22
cycloneive_lcell_comb \Add0~22 (
// Equation(s):
// \Add0~22_combout  = (\portb~44_combout  & ((\porta~101_combout  & (\Add0~21  & VCC)) # (!\porta~101_combout  & (!\Add0~21 )))) # (!\portb~44_combout  & ((\porta~101_combout  & (!\Add0~21 )) # (!\porta~101_combout  & ((\Add0~21 ) # (GND)))))
// \Add0~23  = CARRY((\portb~44_combout  & (!\porta~101_combout  & !\Add0~21 )) # (!\portb~44_combout  & ((!\Add0~21 ) # (!\porta~101_combout ))))

	.dataa(portb20),
	.datab(porta17),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add0~21 ),
	.combout(\Add0~22_combout ),
	.cout(\Add0~23 ));
// synopsys translate_off
defparam \Add0~22 .lut_mask = 16'h9617;
defparam \Add0~22 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X54_Y37_N30
cycloneive_lcell_comb \Selector20~6 (
// Equation(s):
// \Selector20~6_combout  = (\Selector0~9_combout  & \Add0~22_combout )

	.dataa(gnd),
	.datab(gnd),
	.datac(\Selector0~9_combout ),
	.datad(\Add0~22_combout ),
	.cin(gnd),
	.combout(\Selector20~6_combout ),
	.cout());
// synopsys translate_off
defparam \Selector20~6 .lut_mask = 16'hF000;
defparam \Selector20~6 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y38_N22
cycloneive_lcell_comb \Selector20~3 (
// Equation(s):
// \Selector20~3_combout  = (\portb~44_combout ) # ((\porta~101_combout ) # (\Selector0~12_combout ))

	.dataa(portb20),
	.datab(porta17),
	.datac(gnd),
	.datad(\Selector0~12_combout ),
	.cin(gnd),
	.combout(\Selector20~3_combout ),
	.cout());
// synopsys translate_off
defparam \Selector20~3 .lut_mask = 16'hFFEE;
defparam \Selector20~3 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y38_N12
cycloneive_lcell_comb \Selector0~18 (
// Equation(s):
// \Selector0~18_combout  = (!plif_idexaluop_l_1 & (!\ShiftRight0~72_combout  & (!plif_idexaluop_l_2 & !\Selector1~2_combout )))

	.dataa(plif_idexaluop_l_1),
	.datab(\ShiftRight0~72_combout ),
	.datac(plif_idexaluop_l_2),
	.datad(\Selector1~2_combout ),
	.cin(gnd),
	.combout(\Selector0~18_combout ),
	.cout());
// synopsys translate_off
defparam \Selector0~18 .lut_mask = 16'h0001;
defparam \Selector0~18 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y38_N10
cycloneive_lcell_comb \Selector20~4 (
// Equation(s):
// \Selector20~4_combout  = (plif_idexaluop_l_0 & (\ShiftRight0~77_combout  & \Selector0~18_combout ))

	.dataa(gnd),
	.datab(plif_idexaluop_l_0),
	.datac(\ShiftRight0~77_combout ),
	.datad(\Selector0~18_combout ),
	.cin(gnd),
	.combout(\Selector20~4_combout ),
	.cout());
// synopsys translate_off
defparam \Selector20~4 .lut_mask = 16'hC000;
defparam \Selector20~4 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y38_N28
cycloneive_lcell_comb \Selector20~5 (
// Equation(s):
// \Selector20~5_combout  = (\Selector20~4_combout ) # ((\Selector20~3_combout  & ((\Selector20~2_combout ) # (\Selector0~10_combout ))))

	.dataa(\Selector20~2_combout ),
	.datab(\Selector20~3_combout ),
	.datac(\Selector0~10_combout ),
	.datad(\Selector20~4_combout ),
	.cin(gnd),
	.combout(\Selector20~5_combout ),
	.cout());
// synopsys translate_off
defparam \Selector20~5 .lut_mask = 16'hFFC8;
defparam \Selector20~5 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y37_N24
cycloneive_lcell_comb \Selector20~7 (
// Equation(s):
// \Selector20~7_combout  = (\Selector20~6_combout ) # ((\Selector20~5_combout ) # ((\Add1~22_combout  & \Selector0~8_combout )))

	.dataa(\Add1~22_combout ),
	.datab(\Selector0~8_combout ),
	.datac(\Selector20~6_combout ),
	.datad(\Selector20~5_combout ),
	.cin(gnd),
	.combout(\Selector20~7_combout ),
	.cout());
// synopsys translate_off
defparam \Selector20~7 .lut_mask = 16'hFFF8;
defparam \Selector20~7 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y41_N28
cycloneive_lcell_comb \ShiftLeft0~33 (
// Equation(s):
// \ShiftLeft0~33_combout  = (\portb~58_combout  & ((\porta~103_combout ))) # (!\portb~58_combout  & (\porta~102_combout ))

	.dataa(gnd),
	.datab(portb27),
	.datac(porta18),
	.datad(porta19),
	.cin(gnd),
	.combout(\ShiftLeft0~33_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftLeft0~33 .lut_mask = 16'hFC30;
defparam \ShiftLeft0~33 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y41_N26
cycloneive_lcell_comb \ShiftLeft0~34 (
// Equation(s):
// \ShiftLeft0~34_combout  = (\portb~60_combout  & (\ShiftLeft0~27_combout )) # (!\portb~60_combout  & ((\ShiftLeft0~33_combout )))

	.dataa(portb28),
	.datab(gnd),
	.datac(\ShiftLeft0~27_combout ),
	.datad(\ShiftLeft0~33_combout ),
	.cin(gnd),
	.combout(\ShiftLeft0~34_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftLeft0~34 .lut_mask = 16'hF5A0;
defparam \ShiftLeft0~34 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y41_N0
cycloneive_lcell_comb \ShiftLeft0~35 (
// Equation(s):
// \ShiftLeft0~35_combout  = (!\portb~62_combout  & ((\portb~64_combout  & ((\ShiftLeft0~6_combout ))) # (!\portb~64_combout  & (\ShiftLeft0~34_combout ))))

	.dataa(portb29),
	.datab(portb30),
	.datac(\ShiftLeft0~34_combout ),
	.datad(\ShiftLeft0~6_combout ),
	.cin(gnd),
	.combout(\ShiftLeft0~35_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftLeft0~35 .lut_mask = 16'h5410;
defparam \ShiftLeft0~35 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y41_N30
cycloneive_lcell_comb \ShiftLeft0~36 (
// Equation(s):
// \ShiftLeft0~36_combout  = (\ShiftLeft0~35_combout ) # ((\portb~62_combout  & (!\portb~64_combout  & \ShiftLeft0~19_combout )))

	.dataa(portb29),
	.datab(portb30),
	.datac(\ShiftLeft0~19_combout ),
	.datad(\ShiftLeft0~35_combout ),
	.cin(gnd),
	.combout(\ShiftLeft0~36_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftLeft0~36 .lut_mask = 16'hFF20;
defparam \ShiftLeft0~36 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y37_N8
cycloneive_lcell_comb \Selector21~7 (
// Equation(s):
// \Selector21~7_combout  = (\Selector21~0_combout  & ((\Selector0~17_combout ) # ((\ShiftRight0~90_combout  & \Selector20~1_combout )))) # (!\Selector21~0_combout  & (\ShiftRight0~90_combout  & ((\Selector20~1_combout ))))

	.dataa(\Selector21~0_combout ),
	.datab(\ShiftRight0~90_combout ),
	.datac(\Selector0~17_combout ),
	.datad(\Selector20~1_combout ),
	.cin(gnd),
	.combout(\Selector21~7_combout ),
	.cout());
// synopsys translate_off
defparam \Selector21~7 .lut_mask = 16'hECA0;
defparam \Selector21~7 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X50_Y39_N16
cycloneive_lcell_comb \Selector21~4 (
// Equation(s):
// \Selector21~4_combout  = (\porta~102_combout  & (((\Selector0~10_combout )))) # (!\porta~102_combout  & (!\portb~46_combout  & ((\Selector0~12_combout ))))

	.dataa(portb21),
	.datab(\Selector0~10_combout ),
	.datac(porta18),
	.datad(\Selector0~12_combout ),
	.cin(gnd),
	.combout(\Selector21~4_combout ),
	.cout());
// synopsys translate_off
defparam \Selector21~4 .lut_mask = 16'hC5C0;
defparam \Selector21~4 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X50_Y39_N14
cycloneive_lcell_comb \Selector21~2 (
// Equation(s):
// \Selector21~2_combout  = (\portb~46_combout  & ((\Selector0~10_combout ) # ((\Selector0~11_combout  & \porta~102_combout ))))

	.dataa(portb21),
	.datab(\Selector0~11_combout ),
	.datac(porta18),
	.datad(\Selector0~10_combout ),
	.cin(gnd),
	.combout(\Selector21~2_combout ),
	.cout());
// synopsys translate_off
defparam \Selector21~2 .lut_mask = 16'hAA80;
defparam \Selector21~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X50_Y39_N28
cycloneive_lcell_comb \Selector21~1 (
// Equation(s):
// \Selector21~1_combout  = (\Selector0~8_combout  & ((\Add1~20_combout ) # ((\Selector0~9_combout  & \Add0~20_combout )))) # (!\Selector0~8_combout  & (\Selector0~9_combout  & (\Add0~20_combout )))

	.dataa(\Selector0~8_combout ),
	.datab(\Selector0~9_combout ),
	.datac(\Add0~20_combout ),
	.datad(\Add1~20_combout ),
	.cin(gnd),
	.combout(\Selector21~1_combout ),
	.cout());
// synopsys translate_off
defparam \Selector21~1 .lut_mask = 16'hEAC0;
defparam \Selector21~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X50_Y39_N6
cycloneive_lcell_comb \Selector21~5 (
// Equation(s):
// \Selector21~5_combout  = (\Selector21~3_combout ) # ((\Selector21~4_combout ) # ((\Selector21~2_combout ) # (\Selector21~1_combout )))

	.dataa(\Selector21~3_combout ),
	.datab(\Selector21~4_combout ),
	.datac(\Selector21~2_combout ),
	.datad(\Selector21~1_combout ),
	.cin(gnd),
	.combout(\Selector21~5_combout ),
	.cout());
// synopsys translate_off
defparam \Selector21~5 .lut_mask = 16'hFFFE;
defparam \Selector21~5 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y37_N2
cycloneive_lcell_comb \Selector21~6 (
// Equation(s):
// \Selector21~6_combout  = (\Selector21~5_combout ) # ((plif_idexaluop_l_0 & (\ShiftRight0~88_combout  & \Selector0~18_combout )))

	.dataa(plif_idexaluop_l_0),
	.datab(\ShiftRight0~88_combout ),
	.datac(\Selector0~18_combout ),
	.datad(\Selector21~5_combout ),
	.cin(gnd),
	.combout(\Selector21~6_combout ),
	.cout());
// synopsys translate_off
defparam \Selector21~6 .lut_mask = 16'hFF80;
defparam \Selector21~6 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y38_N24
cycloneive_lcell_comb \Selector18~7 (
// Equation(s):
// \Selector18~7_combout  = (plif_idexaluop_l_0 & (\Selector0~15_combout  & (!\Selector1~2_combout  & \ShiftRight0~94_combout )))

	.dataa(plif_idexaluop_l_0),
	.datab(\Selector0~15_combout ),
	.datac(\Selector1~2_combout ),
	.datad(\ShiftRight0~94_combout ),
	.cin(gnd),
	.combout(\Selector18~7_combout ),
	.cout());
// synopsys translate_off
defparam \Selector18~7 .lut_mask = 16'h0800;
defparam \Selector18~7 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y38_N22
cycloneive_lcell_comb \Selector18~6 (
// Equation(s):
// \Selector18~6_combout  = (\Selector0~17_combout  & ((\portb~62_combout  & ((\ShiftRight0~31_combout ))) # (!\portb~62_combout  & (\ShiftRight0~35_combout ))))

	.dataa(portb29),
	.datab(\ShiftRight0~35_combout ),
	.datac(\Selector0~17_combout ),
	.datad(\ShiftRight0~31_combout ),
	.cin(gnd),
	.combout(\Selector18~6_combout ),
	.cout());
// synopsys translate_off
defparam \Selector18~6 .lut_mask = 16'hE040;
defparam \Selector18~6 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y40_N24
cycloneive_lcell_comb \Add1~24 (
// Equation(s):
// \Add1~24_combout  = ((\portb~42_combout  $ (\porta~100_combout  $ (\Add1~23 )))) # (GND)
// \Add1~25  = CARRY((\portb~42_combout  & (\porta~100_combout  & !\Add1~23 )) # (!\portb~42_combout  & ((\porta~100_combout ) # (!\Add1~23 ))))

	.dataa(portb19),
	.datab(porta16),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add1~23 ),
	.combout(\Add1~24_combout ),
	.cout(\Add1~25 ));
// synopsys translate_off
defparam \Add1~24 .lut_mask = 16'h964D;
defparam \Add1~24 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X57_Y40_N26
cycloneive_lcell_comb \Add1~26 (
// Equation(s):
// \Add1~26_combout  = (\portb~40_combout  & ((\porta~99_combout  & (!\Add1~25 )) # (!\porta~99_combout  & ((\Add1~25 ) # (GND))))) # (!\portb~40_combout  & ((\porta~99_combout  & (\Add1~25  & VCC)) # (!\porta~99_combout  & (!\Add1~25 ))))
// \Add1~27  = CARRY((\portb~40_combout  & ((!\Add1~25 ) # (!\porta~99_combout ))) # (!\portb~40_combout  & (!\porta~99_combout  & !\Add1~25 )))

	.dataa(portb18),
	.datab(porta15),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add1~25 ),
	.combout(\Add1~26_combout ),
	.cout(\Add1~27 ));
// synopsys translate_off
defparam \Add1~26 .lut_mask = 16'h692B;
defparam \Add1~26 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X53_Y38_N18
cycloneive_lcell_comb \Selector18~8 (
// Equation(s):
// \Selector18~8_combout  = (\Selector18~7_combout ) # ((\Selector18~6_combout ) # ((\Selector0~8_combout  & \Add1~26_combout )))

	.dataa(\Selector0~8_combout ),
	.datab(\Selector18~7_combout ),
	.datac(\Selector18~6_combout ),
	.datad(\Add1~26_combout ),
	.cin(gnd),
	.combout(\Selector18~8_combout ),
	.cout());
// synopsys translate_off
defparam \Selector18~8 .lut_mask = 16'hFEFC;
defparam \Selector18~8 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X52_Y38_N24
cycloneive_lcell_comb \Add0~24 (
// Equation(s):
// \Add0~24_combout  = ((\portb~42_combout  $ (\porta~100_combout  $ (!\Add0~23 )))) # (GND)
// \Add0~25  = CARRY((\portb~42_combout  & ((\porta~100_combout ) # (!\Add0~23 ))) # (!\portb~42_combout  & (\porta~100_combout  & !\Add0~23 )))

	.dataa(portb19),
	.datab(porta16),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add0~23 ),
	.combout(\Add0~24_combout ),
	.cout(\Add0~25 ));
// synopsys translate_off
defparam \Add0~24 .lut_mask = 16'h698E;
defparam \Add0~24 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X52_Y38_N26
cycloneive_lcell_comb \Add0~26 (
// Equation(s):
// \Add0~26_combout  = (\portb~40_combout  & ((\porta~99_combout  & (\Add0~25  & VCC)) # (!\porta~99_combout  & (!\Add0~25 )))) # (!\portb~40_combout  & ((\porta~99_combout  & (!\Add0~25 )) # (!\porta~99_combout  & ((\Add0~25 ) # (GND)))))
// \Add0~27  = CARRY((\portb~40_combout  & (!\porta~99_combout  & !\Add0~25 )) # (!\portb~40_combout  & ((!\Add0~25 ) # (!\porta~99_combout ))))

	.dataa(portb18),
	.datab(porta15),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add0~25 ),
	.combout(\Add0~26_combout ),
	.cout(\Add0~27 ));
// synopsys translate_off
defparam \Add0~26 .lut_mask = 16'h9617;
defparam \Add0~26 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X53_Y41_N26
cycloneive_lcell_comb \Selector18~0 (
// Equation(s):
// \Selector18~0_combout  = (\porta~99_combout  & (((\Selector0~10_combout )))) # (!\porta~99_combout  & (\Selector0~12_combout  & ((!\portb~40_combout ))))

	.dataa(\Selector0~12_combout ),
	.datab(porta15),
	.datac(\Selector0~10_combout ),
	.datad(portb18),
	.cin(gnd),
	.combout(\Selector18~0_combout ),
	.cout());
// synopsys translate_off
defparam \Selector18~0 .lut_mask = 16'hC0E2;
defparam \Selector18~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y41_N8
cycloneive_lcell_comb \Selector18~1 (
// Equation(s):
// \Selector18~1_combout  = (\Selector18~0_combout ) # ((\Selector0~13_combout  & (\portb~40_combout  $ (\porta~99_combout ))))

	.dataa(portb18),
	.datab(\Selector0~13_combout ),
	.datac(\Selector18~0_combout ),
	.datad(porta15),
	.cin(gnd),
	.combout(\Selector18~1_combout ),
	.cout());
// synopsys translate_off
defparam \Selector18~1 .lut_mask = 16'hF4F8;
defparam \Selector18~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y36_N18
cycloneive_lcell_comb \ShiftLeft0~37 (
// Equation(s):
// \ShiftLeft0~37_combout  = (\portb~58_combout  & (\porta~100_combout )) # (!\portb~58_combout  & ((\porta~99_combout )))

	.dataa(gnd),
	.datab(porta16),
	.datac(portb27),
	.datad(porta15),
	.cin(gnd),
	.combout(\ShiftLeft0~37_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftLeft0~37 .lut_mask = 16'hCFC0;
defparam \ShiftLeft0~37 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y38_N14
cycloneive_lcell_comb \ShiftLeft0~38 (
// Equation(s):
// \ShiftLeft0~38_combout  = (\portb~60_combout  & ((\ShiftLeft0~29_combout ))) # (!\portb~60_combout  & (\ShiftLeft0~37_combout ))

	.dataa(portb28),
	.datab(gnd),
	.datac(\ShiftLeft0~37_combout ),
	.datad(\ShiftLeft0~29_combout ),
	.cin(gnd),
	.combout(\ShiftLeft0~38_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftLeft0~38 .lut_mask = 16'hFA50;
defparam \ShiftLeft0~38 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X52_Y41_N0
cycloneive_lcell_comb \ShiftLeft0~15 (
// Equation(s):
// \ShiftLeft0~15_combout  = (\portb~58_combout  & ((\porta~94_combout ))) # (!\portb~58_combout  & (\porta~93_combout ))

	.dataa(porta9),
	.datab(gnd),
	.datac(porta10),
	.datad(portb27),
	.cin(gnd),
	.combout(\ShiftLeft0~15_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftLeft0~15 .lut_mask = 16'hF0AA;
defparam \ShiftLeft0~15 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X52_Y41_N26
cycloneive_lcell_comb \ShiftLeft0~24 (
// Equation(s):
// \ShiftLeft0~24_combout  = (\portb~60_combout  & (\ShiftLeft0~15_combout )) # (!\portb~60_combout  & ((\ShiftLeft0~23_combout )))

	.dataa(gnd),
	.datab(\ShiftLeft0~15_combout ),
	.datac(portb28),
	.datad(\ShiftLeft0~23_combout ),
	.cin(gnd),
	.combout(\ShiftLeft0~24_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftLeft0~24 .lut_mask = 16'hCFC0;
defparam \ShiftLeft0~24 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y38_N8
cycloneive_lcell_comb \Selector10~0 (
// Equation(s):
// \Selector10~0_combout  = (\portb~62_combout  & ((\ShiftLeft0~24_combout ))) # (!\portb~62_combout  & (\ShiftLeft0~38_combout ))

	.dataa(portb29),
	.datab(gnd),
	.datac(\ShiftLeft0~38_combout ),
	.datad(\ShiftLeft0~24_combout ),
	.cin(gnd),
	.combout(\Selector10~0_combout ),
	.cout());
// synopsys translate_off
defparam \Selector10~0 .lut_mask = 16'hFA50;
defparam \Selector10~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y38_N6
cycloneive_lcell_comb \ShiftLeft0~39 (
// Equation(s):
// \ShiftLeft0~39_combout  = (\portb~64_combout  & ((\ShiftLeft0~9_combout ))) # (!\portb~64_combout  & (\Selector10~0_combout ))

	.dataa(gnd),
	.datab(portb30),
	.datac(\Selector10~0_combout ),
	.datad(\ShiftLeft0~9_combout ),
	.cin(gnd),
	.combout(\ShiftLeft0~39_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftLeft0~39 .lut_mask = 16'hFC30;
defparam \ShiftLeft0~39 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y38_N26
cycloneive_lcell_comb \Selector18~4 (
// Equation(s):
// \Selector18~4_combout  = (\Selector18~3_combout  & ((\ShiftRight0~28_combout ) # ((\Selector16~0_combout  & \ShiftLeft0~39_combout )))) # (!\Selector18~3_combout  & (\Selector16~0_combout  & ((\ShiftLeft0~39_combout ))))

	.dataa(\Selector18~3_combout ),
	.datab(\Selector16~0_combout ),
	.datac(\ShiftRight0~28_combout ),
	.datad(\ShiftLeft0~39_combout ),
	.cin(gnd),
	.combout(\Selector18~4_combout ),
	.cout());
// synopsys translate_off
defparam \Selector18~4 .lut_mask = 16'hECA0;
defparam \Selector18~4 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X52_Y35_N22
cycloneive_lcell_comb \Selector18~2 (
// Equation(s):
// \Selector18~2_combout  = (\Selector0~10_combout ) # ((\porta~99_combout  & \Selector0~11_combout ))

	.dataa(\Selector0~10_combout ),
	.datab(porta15),
	.datac(\Selector0~11_combout ),
	.datad(gnd),
	.cin(gnd),
	.combout(\Selector18~2_combout ),
	.cout());
// synopsys translate_off
defparam \Selector18~2 .lut_mask = 16'hEAEA;
defparam \Selector18~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y38_N20
cycloneive_lcell_comb \Selector18~5 (
// Equation(s):
// \Selector18~5_combout  = (\Selector18~1_combout ) # ((\Selector18~4_combout ) # ((\portb~40_combout  & \Selector18~2_combout )))

	.dataa(\Selector18~1_combout ),
	.datab(portb18),
	.datac(\Selector18~4_combout ),
	.datad(\Selector18~2_combout ),
	.cin(gnd),
	.combout(\Selector18~5_combout ),
	.cout());
// synopsys translate_off
defparam \Selector18~5 .lut_mask = 16'hFEFA;
defparam \Selector18~5 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y40_N22
cycloneive_lcell_comb \Selector19~6 (
// Equation(s):
// \Selector19~6_combout  = (\Selector0~17_combout  & ((\portb~62_combout  & ((\ShiftRight0~62_combout ))) # (!\portb~62_combout  & (\ShiftRight0~66_combout ))))

	.dataa(portb29),
	.datab(\ShiftRight0~66_combout ),
	.datac(\ShiftRight0~62_combout ),
	.datad(\Selector0~17_combout ),
	.cin(gnd),
	.combout(\Selector19~6_combout ),
	.cout());
// synopsys translate_off
defparam \Selector19~6 .lut_mask = 16'hE400;
defparam \Selector19~6 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y38_N24
cycloneive_lcell_comb \ShiftLeft0~40 (
// Equation(s):
// \ShiftLeft0~40_combout  = (\portb~58_combout  & (\porta~101_combout )) # (!\portb~58_combout  & ((\porta~100_combout )))

	.dataa(porta17),
	.datab(gnd),
	.datac(porta16),
	.datad(portb27),
	.cin(gnd),
	.combout(\ShiftLeft0~40_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftLeft0~40 .lut_mask = 16'hAAF0;
defparam \ShiftLeft0~40 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y40_N10
cycloneive_lcell_comb \ShiftLeft0~41 (
// Equation(s):
// \ShiftLeft0~41_combout  = (\portb~60_combout  & ((\ShiftLeft0~33_combout ))) # (!\portb~60_combout  & (\ShiftLeft0~40_combout ))

	.dataa(portb28),
	.datab(gnd),
	.datac(\ShiftLeft0~40_combout ),
	.datad(\ShiftLeft0~33_combout ),
	.cin(gnd),
	.combout(\ShiftLeft0~41_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftLeft0~41 .lut_mask = 16'hFA50;
defparam \ShiftLeft0~41 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y40_N16
cycloneive_lcell_comb \Selector11~0 (
// Equation(s):
// \Selector11~0_combout  = (\portb~62_combout  & (\ShiftLeft0~28_combout )) # (!\portb~62_combout  & ((\ShiftLeft0~41_combout )))

	.dataa(gnd),
	.datab(portb29),
	.datac(\ShiftLeft0~28_combout ),
	.datad(\ShiftLeft0~41_combout ),
	.cin(gnd),
	.combout(\Selector11~0_combout ),
	.cout());
// synopsys translate_off
defparam \Selector11~0 .lut_mask = 16'hF3C0;
defparam \Selector11~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y40_N0
cycloneive_lcell_comb \Selector19~0 (
// Equation(s):
// \Selector19~0_combout  = (\Selector16~0_combout  & ((\portb~64_combout  & (\ShiftLeft0~14_combout )) # (!\portb~64_combout  & ((\Selector11~0_combout )))))

	.dataa(portb30),
	.datab(\ShiftLeft0~14_combout ),
	.datac(\Selector16~0_combout ),
	.datad(\Selector11~0_combout ),
	.cin(gnd),
	.combout(\Selector19~0_combout ),
	.cout());
// synopsys translate_off
defparam \Selector19~0 .lut_mask = 16'hD080;
defparam \Selector19~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X50_Y40_N28
cycloneive_lcell_comb \Selector19~3 (
// Equation(s):
// \Selector19~3_combout  = (\porta~100_combout  & ((\Selector0~10_combout ) # (!\portb~42_combout ))) # (!\porta~100_combout  & ((\portb~42_combout )))

	.dataa(gnd),
	.datab(\Selector0~10_combout ),
	.datac(porta16),
	.datad(portb19),
	.cin(gnd),
	.combout(\Selector19~3_combout ),
	.cout());
// synopsys translate_off
defparam \Selector19~3 .lut_mask = 16'hCFF0;
defparam \Selector19~3 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X50_Y40_N10
cycloneive_lcell_comb \Selector19~4 (
// Equation(s):
// \Selector19~4_combout  = (\Selector19~3_combout  & (((\Selector0~10_combout ) # (\Selector0~13_combout )))) # (!\Selector19~3_combout  & (\Selector19~2_combout ))

	.dataa(\Selector19~2_combout ),
	.datab(\Selector0~10_combout ),
	.datac(\Selector0~13_combout ),
	.datad(\Selector19~3_combout ),
	.cin(gnd),
	.combout(\Selector19~4_combout ),
	.cout());
// synopsys translate_off
defparam \Selector19~4 .lut_mask = 16'hFCAA;
defparam \Selector19~4 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y40_N18
cycloneive_lcell_comb \Selector19~1 (
// Equation(s):
// \Selector19~1_combout  = (!\portb~64_combout  & (!\portb~62_combout  & (\ShiftRight0~59_combout  & \Selector23~1_combout )))

	.dataa(portb30),
	.datab(portb29),
	.datac(\ShiftRight0~59_combout ),
	.datad(\Selector23~1_combout ),
	.cin(gnd),
	.combout(\Selector19~1_combout ),
	.cout());
// synopsys translate_off
defparam \Selector19~1 .lut_mask = 16'h1000;
defparam \Selector19~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y40_N4
cycloneive_lcell_comb \Selector19~5 (
// Equation(s):
// \Selector19~5_combout  = (\Selector19~4_combout ) # ((\Selector19~1_combout ) # ((\ShiftRight0~97_combout  & \Selector16~1_combout )))

	.dataa(\ShiftRight0~97_combout ),
	.datab(\Selector16~1_combout ),
	.datac(\Selector19~4_combout ),
	.datad(\Selector19~1_combout ),
	.cin(gnd),
	.combout(\Selector19~5_combout ),
	.cout());
// synopsys translate_off
defparam \Selector19~5 .lut_mask = 16'hFFF8;
defparam \Selector19~5 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y40_N16
cycloneive_lcell_comb \Selector19~7 (
// Equation(s):
// \Selector19~7_combout  = (\Selector0~8_combout  & ((\Add1~24_combout ) # ((\Selector0~9_combout  & \Add0~24_combout )))) # (!\Selector0~8_combout  & (\Selector0~9_combout  & ((\Add0~24_combout ))))

	.dataa(\Selector0~8_combout ),
	.datab(\Selector0~9_combout ),
	.datac(\Add1~24_combout ),
	.datad(\Add0~24_combout ),
	.cin(gnd),
	.combout(\Selector19~7_combout ),
	.cout());
// synopsys translate_off
defparam \Selector19~7 .lut_mask = 16'hECA0;
defparam \Selector19~7 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y40_N28
cycloneive_lcell_comb \Add1~28 (
// Equation(s):
// \Add1~28_combout  = ((\porta~98_combout  $ (\portb~38_combout  $ (\Add1~27 )))) # (GND)
// \Add1~29  = CARRY((\porta~98_combout  & ((!\Add1~27 ) # (!\portb~38_combout ))) # (!\porta~98_combout  & (!\portb~38_combout  & !\Add1~27 )))

	.dataa(porta14),
	.datab(portb17),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add1~27 ),
	.combout(\Add1~28_combout ),
	.cout(\Add1~29 ));
// synopsys translate_off
defparam \Add1~28 .lut_mask = 16'h962B;
defparam \Add1~28 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X57_Y40_N30
cycloneive_lcell_comb \Add1~30 (
// Equation(s):
// \Add1~30_combout  = (\porta~97_combout  & ((\portb~36_combout  & (!\Add1~29 )) # (!\portb~36_combout  & (\Add1~29  & VCC)))) # (!\porta~97_combout  & ((\portb~36_combout  & ((\Add1~29 ) # (GND))) # (!\portb~36_combout  & (!\Add1~29 ))))
// \Add1~31  = CARRY((\porta~97_combout  & (\portb~36_combout  & !\Add1~29 )) # (!\porta~97_combout  & ((\portb~36_combout ) # (!\Add1~29 ))))

	.dataa(porta13),
	.datab(portb16),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add1~29 ),
	.combout(\Add1~30_combout ),
	.cout(\Add1~31 ));
// synopsys translate_off
defparam \Add1~30 .lut_mask = 16'h694D;
defparam \Add1~30 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X50_Y36_N16
cycloneive_lcell_comb \Selector16~3 (
// Equation(s):
// \Selector16~3_combout  = (\portb~36_combout  & ((\Selector0~10_combout ) # ((\porta~97_combout  & \Selector0~11_combout ))))

	.dataa(\Selector0~10_combout ),
	.datab(porta13),
	.datac(\Selector0~11_combout ),
	.datad(portb16),
	.cin(gnd),
	.combout(\Selector16~3_combout ),
	.cout());
// synopsys translate_off
defparam \Selector16~3 .lut_mask = 16'hEA00;
defparam \Selector16~3 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X50_Y36_N14
cycloneive_lcell_comb \Selector16~2 (
// Equation(s):
// \Selector16~2_combout  = (\porta~97_combout  & (\Selector0~10_combout )) # (!\porta~97_combout  & (((\Selector0~12_combout  & !\portb~36_combout ))))

	.dataa(\Selector0~10_combout ),
	.datab(\Selector0~12_combout ),
	.datac(porta13),
	.datad(portb16),
	.cin(gnd),
	.combout(\Selector16~2_combout ),
	.cout());
// synopsys translate_off
defparam \Selector16~2 .lut_mask = 16'hA0AC;
defparam \Selector16~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X52_Y38_N28
cycloneive_lcell_comb \Add0~28 (
// Equation(s):
// \Add0~28_combout  = ((\portb~38_combout  $ (\porta~98_combout  $ (!\Add0~27 )))) # (GND)
// \Add0~29  = CARRY((\portb~38_combout  & ((\porta~98_combout ) # (!\Add0~27 ))) # (!\portb~38_combout  & (\porta~98_combout  & !\Add0~27 )))

	.dataa(portb17),
	.datab(porta14),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add0~27 ),
	.combout(\Add0~28_combout ),
	.cout(\Add0~29 ));
// synopsys translate_off
defparam \Add0~28 .lut_mask = 16'h698E;
defparam \Add0~28 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X52_Y38_N30
cycloneive_lcell_comb \Add0~30 (
// Equation(s):
// \Add0~30_combout  = (\porta~97_combout  & ((\portb~36_combout  & (\Add0~29  & VCC)) # (!\portb~36_combout  & (!\Add0~29 )))) # (!\porta~97_combout  & ((\portb~36_combout  & (!\Add0~29 )) # (!\portb~36_combout  & ((\Add0~29 ) # (GND)))))
// \Add0~31  = CARRY((\porta~97_combout  & (!\portb~36_combout  & !\Add0~29 )) # (!\porta~97_combout  & ((!\Add0~29 ) # (!\portb~36_combout ))))

	.dataa(porta13),
	.datab(portb16),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add0~29 ),
	.combout(\Add0~30_combout ),
	.cout(\Add0~31 ));
// synopsys translate_off
defparam \Add0~30 .lut_mask = 16'h9617;
defparam \Add0~30 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X50_Y36_N6
cycloneive_lcell_comb \Selector16~4 (
// Equation(s):
// \Selector16~4_combout  = (\Selector16~3_combout ) # ((\Selector16~2_combout ) # ((\Selector0~9_combout  & \Add0~30_combout )))

	.dataa(\Selector0~9_combout ),
	.datab(\Selector16~3_combout ),
	.datac(\Selector16~2_combout ),
	.datad(\Add0~30_combout ),
	.cin(gnd),
	.combout(\Selector16~4_combout ),
	.cout());
// synopsys translate_off
defparam \Selector16~4 .lut_mask = 16'hFEFC;
defparam \Selector16~4 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X52_Y35_N0
cycloneive_lcell_comb \Selector16~5 (
// Equation(s):
// \Selector16~5_combout  = (plif_idexaluop_l_0 & (!\ShiftRight0~71_combout  & (\portb~66_combout  & \Selector1~3_combout )))

	.dataa(plif_idexaluop_l_0),
	.datab(\ShiftRight0~71_combout ),
	.datac(portb31),
	.datad(\Selector1~3_combout ),
	.cin(gnd),
	.combout(\Selector16~5_combout ),
	.cout());
// synopsys translate_off
defparam \Selector16~5 .lut_mask = 16'h2000;
defparam \Selector16~5 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X52_Y36_N20
cycloneive_lcell_comb \Selector16~7 (
// Equation(s):
// \Selector16~7_combout  = (\Selector0~17_combout  & ((\portb~62_combout  & ((\ShiftRight0~80_combout ))) # (!\portb~62_combout  & (\ShiftRight0~82_combout ))))

	.dataa(portb29),
	.datab(\ShiftRight0~82_combout ),
	.datac(\ShiftRight0~80_combout ),
	.datad(\Selector0~17_combout ),
	.cin(gnd),
	.combout(\Selector16~7_combout ),
	.cout());
// synopsys translate_off
defparam \Selector16~7 .lut_mask = 16'hE400;
defparam \Selector16~7 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X52_Y36_N30
cycloneive_lcell_comb \Selector16~8 (
// Equation(s):
// \Selector16~8_combout  = (\Selector16~7_combout ) # ((\Selector0~13_combout  & (\porta~97_combout  $ (\portb~36_combout ))))

	.dataa(porta13),
	.datab(portb16),
	.datac(\Selector0~13_combout ),
	.datad(\Selector16~7_combout ),
	.cin(gnd),
	.combout(\Selector16~8_combout ),
	.cout());
// synopsys translate_off
defparam \Selector16~8 .lut_mask = 16'hFF60;
defparam \Selector16~8 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y36_N28
cycloneive_lcell_comb \ShiftLeft0~42 (
// Equation(s):
// \ShiftLeft0~42_combout  = (\portb~58_combout  & ((\porta~98_combout ))) # (!\portb~58_combout  & (\porta~97_combout ))

	.dataa(portb27),
	.datab(gnd),
	.datac(porta13),
	.datad(porta14),
	.cin(gnd),
	.combout(\ShiftLeft0~42_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftLeft0~42 .lut_mask = 16'hFA50;
defparam \ShiftLeft0~42 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X52_Y36_N4
cycloneive_lcell_comb \ShiftLeft0~43 (
// Equation(s):
// \ShiftLeft0~43_combout  = (\portb~60_combout  & (\ShiftLeft0~37_combout )) # (!\portb~60_combout  & ((\ShiftLeft0~42_combout )))

	.dataa(portb28),
	.datab(gnd),
	.datac(\ShiftLeft0~37_combout ),
	.datad(\ShiftLeft0~42_combout ),
	.cin(gnd),
	.combout(\ShiftLeft0~43_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftLeft0~43 .lut_mask = 16'hF5A0;
defparam \ShiftLeft0~43 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X52_Y36_N6
cycloneive_lcell_comb \Selector8~0 (
// Equation(s):
// \Selector8~0_combout  = (\portb~62_combout  & ((\ShiftLeft0~30_combout ))) # (!\portb~62_combout  & (\ShiftLeft0~43_combout ))

	.dataa(portb29),
	.datab(gnd),
	.datac(\ShiftLeft0~43_combout ),
	.datad(\ShiftLeft0~30_combout ),
	.cin(gnd),
	.combout(\Selector8~0_combout ),
	.cout());
// synopsys translate_off
defparam \Selector8~0 .lut_mask = 16'hFA50;
defparam \Selector8~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X52_Y36_N12
cycloneive_lcell_comb \ShiftLeft0~44 (
// Equation(s):
// \ShiftLeft0~44_combout  = (\portb~64_combout  & (\ShiftLeft0~17_combout )) # (!\portb~64_combout  & ((\Selector8~0_combout )))

	.dataa(gnd),
	.datab(portb30),
	.datac(\ShiftLeft0~17_combout ),
	.datad(\Selector8~0_combout ),
	.cin(gnd),
	.combout(\ShiftLeft0~44_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftLeft0~44 .lut_mask = 16'hF3C0;
defparam \ShiftLeft0~44 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X52_Y36_N18
cycloneive_lcell_comb \Selector16~6 (
// Equation(s):
// \Selector16~6_combout  = (\ShiftRight0~100_combout  & ((\Selector16~1_combout ) # ((\Selector16~0_combout  & \ShiftLeft0~44_combout )))) # (!\ShiftRight0~100_combout  & (\Selector16~0_combout  & ((\ShiftLeft0~44_combout ))))

	.dataa(\ShiftRight0~100_combout ),
	.datab(\Selector16~0_combout ),
	.datac(\Selector16~1_combout ),
	.datad(\ShiftLeft0~44_combout ),
	.cin(gnd),
	.combout(\Selector16~6_combout ),
	.cout());
// synopsys translate_off
defparam \Selector16~6 .lut_mask = 16'hECA0;
defparam \Selector16~6 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X52_Y36_N16
cycloneive_lcell_comb \Selector16~9 (
// Equation(s):
// \Selector16~9_combout  = (\Selector16~8_combout ) # ((\Selector16~6_combout ) # ((\porta~104_combout  & \Selector16~5_combout )))

	.dataa(porta20),
	.datab(\Selector16~5_combout ),
	.datac(\Selector16~8_combout ),
	.datad(\Selector16~6_combout ),
	.cin(gnd),
	.combout(\Selector16~9_combout ),
	.cout());
// synopsys translate_off
defparam \Selector16~9 .lut_mask = 16'hFFF8;
defparam \Selector16~9 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y39_N12
cycloneive_lcell_comb \Selector17~4 (
// Equation(s):
// \Selector17~4_combout  = (\Selector0~17_combout  & ((\portb~62_combout  & (\ShiftRight0~89_combout )) # (!\portb~62_combout  & ((\ShiftRight0~91_combout )))))

	.dataa(\ShiftRight0~89_combout ),
	.datab(\ShiftRight0~91_combout ),
	.datac(portb29),
	.datad(\Selector0~17_combout ),
	.cin(gnd),
	.combout(\Selector17~4_combout ),
	.cout());
// synopsys translate_off
defparam \Selector17~4 .lut_mask = 16'hAC00;
defparam \Selector17~4 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y39_N10
cycloneive_lcell_comb \Selector17~5 (
// Equation(s):
// \Selector17~5_combout  = (\portb~38_combout  & ((\Selector0~10_combout ) # ((\Selector0~11_combout  & \porta~98_combout ))))

	.dataa(\Selector0~11_combout ),
	.datab(portb17),
	.datac(\Selector0~10_combout ),
	.datad(porta14),
	.cin(gnd),
	.combout(\Selector17~5_combout ),
	.cout());
// synopsys translate_off
defparam \Selector17~5 .lut_mask = 16'hC8C0;
defparam \Selector17~5 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y39_N18
cycloneive_lcell_comb \Selector17~6 (
// Equation(s):
// \Selector17~6_combout  = (\Selector17~4_combout ) # ((\Selector17~5_combout ) # ((\Selector0~8_combout  & \Add1~28_combout )))

	.dataa(\Selector17~4_combout ),
	.datab(\Selector0~8_combout ),
	.datac(\Selector17~5_combout ),
	.datad(\Add1~28_combout ),
	.cin(gnd),
	.combout(\Selector17~6_combout ),
	.cout());
// synopsys translate_off
defparam \Selector17~6 .lut_mask = 16'hFEFA;
defparam \Selector17~6 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X50_Y40_N8
cycloneive_lcell_comb \Selector17~2 (
// Equation(s):
// \Selector17~2_combout  = (\portb~38_combout  & (\Selector0~13_combout  & ((!\porta~98_combout )))) # (!\portb~38_combout  & ((\porta~98_combout  & (\Selector0~13_combout )) # (!\porta~98_combout  & ((\Selector0~12_combout )))))

	.dataa(portb17),
	.datab(\Selector0~13_combout ),
	.datac(\Selector0~12_combout ),
	.datad(porta14),
	.cin(gnd),
	.combout(\Selector17~2_combout ),
	.cout());
// synopsys translate_off
defparam \Selector17~2 .lut_mask = 16'h44D8;
defparam \Selector17~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y41_N24
cycloneive_lcell_comb \ShiftLeft0~46 (
// Equation(s):
// \ShiftLeft0~46_combout  = (\portb~60_combout  & ((\ShiftLeft0~40_combout ))) # (!\portb~60_combout  & (\ShiftLeft0~45_combout ))

	.dataa(\ShiftLeft0~45_combout ),
	.datab(gnd),
	.datac(\ShiftLeft0~40_combout ),
	.datad(portb28),
	.cin(gnd),
	.combout(\ShiftLeft0~46_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftLeft0~46 .lut_mask = 16'hF0AA;
defparam \ShiftLeft0~46 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y41_N2
cycloneive_lcell_comb \Selector9~0 (
// Equation(s):
// \Selector9~0_combout  = (\portb~62_combout  & (\ShiftLeft0~34_combout )) # (!\portb~62_combout  & ((\ShiftLeft0~46_combout )))

	.dataa(portb29),
	.datab(gnd),
	.datac(\ShiftLeft0~34_combout ),
	.datad(\ShiftLeft0~46_combout ),
	.cin(gnd),
	.combout(\Selector9~0_combout ),
	.cout());
// synopsys translate_off
defparam \Selector9~0 .lut_mask = 16'hF5A0;
defparam \Selector9~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y41_N12
cycloneive_lcell_comb \ShiftLeft0~47 (
// Equation(s):
// \ShiftLeft0~47_combout  = (\portb~64_combout  & (\ShiftLeft0~20_combout )) # (!\portb~64_combout  & ((\Selector9~0_combout )))

	.dataa(portb30),
	.datab(gnd),
	.datac(\ShiftLeft0~20_combout ),
	.datad(\Selector9~0_combout ),
	.cin(gnd),
	.combout(\ShiftLeft0~47_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftLeft0~47 .lut_mask = 16'hF5A0;
defparam \ShiftLeft0~47 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y39_N2
cycloneive_lcell_comb \Selector17~0 (
// Equation(s):
// \Selector17~0_combout  = (\Selector16~0_combout  & ((\ShiftLeft0~47_combout ) # ((\Selector16~1_combout  & \ShiftRight0~102_combout )))) # (!\Selector16~0_combout  & (\Selector16~1_combout  & (\ShiftRight0~102_combout )))

	.dataa(\Selector16~0_combout ),
	.datab(\Selector16~1_combout ),
	.datac(\ShiftRight0~102_combout ),
	.datad(\ShiftLeft0~47_combout ),
	.cin(gnd),
	.combout(\Selector17~0_combout ),
	.cout());
// synopsys translate_off
defparam \Selector17~0 .lut_mask = 16'hEAC0;
defparam \Selector17~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y39_N28
cycloneive_lcell_comb \Selector17~1 (
// Equation(s):
// \Selector17~1_combout  = (\Selector17~0_combout ) # ((\ShiftRight0~57_combout  & (!\Selector1~0_combout  & \Selector20~1_combout )))

	.dataa(\ShiftRight0~57_combout ),
	.datab(\Selector1~0_combout ),
	.datac(\Selector20~1_combout ),
	.datad(\Selector17~0_combout ),
	.cin(gnd),
	.combout(\Selector17~1_combout ),
	.cout());
// synopsys translate_off
defparam \Selector17~1 .lut_mask = 16'hFF20;
defparam \Selector17~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y39_N18
cycloneive_lcell_comb \Selector17~3 (
// Equation(s):
// \Selector17~3_combout  = (\Selector17~2_combout ) # ((\Selector17~1_combout ) # ((\Selector0~10_combout  & \porta~98_combout )))

	.dataa(\Selector0~10_combout ),
	.datab(porta14),
	.datac(\Selector17~2_combout ),
	.datad(\Selector17~1_combout ),
	.cin(gnd),
	.combout(\Selector17~3_combout ),
	.cout());
// synopsys translate_off
defparam \Selector17~3 .lut_mask = 16'hFFF8;
defparam \Selector17~3 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y39_N0
cycloneive_lcell_comb \Add1~32 (
// Equation(s):
// \Add1~32_combout  = ((\portb~34_combout  $ (\porta~96_combout  $ (\Add1~31 )))) # (GND)
// \Add1~33  = CARRY((\portb~34_combout  & (\porta~96_combout  & !\Add1~31 )) # (!\portb~34_combout  & ((\porta~96_combout ) # (!\Add1~31 ))))

	.dataa(portb15),
	.datab(porta12),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add1~31 ),
	.combout(\Add1~32_combout ),
	.cout(\Add1~33 ));
// synopsys translate_off
defparam \Add1~32 .lut_mask = 16'h964D;
defparam \Add1~32 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X57_Y39_N2
cycloneive_lcell_comb \Add1~34 (
// Equation(s):
// \Add1~34_combout  = (\porta~118_combout  & ((\portb~32_combout  & (!\Add1~33 )) # (!\portb~32_combout  & (\Add1~33  & VCC)))) # (!\porta~118_combout  & ((\portb~32_combout  & ((\Add1~33 ) # (GND))) # (!\portb~32_combout  & (!\Add1~33 ))))
// \Add1~35  = CARRY((\porta~118_combout  & (\portb~32_combout  & !\Add1~33 )) # (!\porta~118_combout  & ((\portb~32_combout ) # (!\Add1~33 ))))

	.dataa(porta34),
	.datab(portb14),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add1~33 ),
	.combout(\Add1~34_combout ),
	.cout(\Add1~35 ));
// synopsys translate_off
defparam \Add1~34 .lut_mask = 16'h694D;
defparam \Add1~34 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X53_Y37_N18
cycloneive_lcell_comb \Selector1~4 (
// Equation(s):
// \Selector1~4_combout  = (\portb~66_combout  & (!plif_idexaluop_l_0 & (!plif_idexaluop_l_3 & \Selector0~15_combout )))

	.dataa(portb31),
	.datab(plif_idexaluop_l_0),
	.datac(plif_idexaluop_l_3),
	.datad(\Selector0~15_combout ),
	.cin(gnd),
	.combout(\Selector1~4_combout ),
	.cout());
// synopsys translate_off
defparam \Selector1~4 .lut_mask = 16'h0200;
defparam \Selector1~4 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y41_N2
cycloneive_lcell_comb \Selector14~6 (
// Equation(s):
// \Selector14~6_combout  = (!\portb~64_combout  & (\ShiftLeft0~2_combout  & (!\Selector1~0_combout  & \Selector1~4_combout )))

	.dataa(portb30),
	.datab(\ShiftLeft0~2_combout ),
	.datac(\Selector1~0_combout ),
	.datad(\Selector1~4_combout ),
	.cin(gnd),
	.combout(\Selector14~6_combout ),
	.cout());
// synopsys translate_off
defparam \Selector14~6 .lut_mask = 16'h0400;
defparam \Selector14~6 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y41_N12
cycloneive_lcell_comb \Selector14~7 (
// Equation(s):
// \Selector14~7_combout  = (\Selector14~6_combout ) # ((\Selector0~8_combout  & \Add1~34_combout ))

	.dataa(\Selector0~8_combout ),
	.datab(gnd),
	.datac(\Add1~34_combout ),
	.datad(\Selector14~6_combout ),
	.cin(gnd),
	.combout(\Selector14~7_combout ),
	.cout());
// synopsys translate_off
defparam \Selector14~7 .lut_mask = 16'hFFA0;
defparam \Selector14~7 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X52_Y37_N0
cycloneive_lcell_comb \Add0~32 (
// Equation(s):
// \Add0~32_combout  = ((\porta~96_combout  $ (\portb~34_combout  $ (!\Add0~31 )))) # (GND)
// \Add0~33  = CARRY((\porta~96_combout  & ((\portb~34_combout ) # (!\Add0~31 ))) # (!\porta~96_combout  & (\portb~34_combout  & !\Add0~31 )))

	.dataa(porta12),
	.datab(portb15),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add0~31 ),
	.combout(\Add0~32_combout ),
	.cout(\Add0~33 ));
// synopsys translate_off
defparam \Add0~32 .lut_mask = 16'h698E;
defparam \Add0~32 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X52_Y37_N2
cycloneive_lcell_comb \Add0~34 (
// Equation(s):
// \Add0~34_combout  = (\porta~118_combout  & ((\portb~32_combout  & (\Add0~33  & VCC)) # (!\portb~32_combout  & (!\Add0~33 )))) # (!\porta~118_combout  & ((\portb~32_combout  & (!\Add0~33 )) # (!\portb~32_combout  & ((\Add0~33 ) # (GND)))))
// \Add0~35  = CARRY((\porta~118_combout  & (!\portb~32_combout  & !\Add0~33 )) # (!\porta~118_combout  & ((!\Add0~33 ) # (!\portb~32_combout ))))

	.dataa(porta34),
	.datab(portb14),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add0~33 ),
	.combout(\Add0~34_combout ),
	.cout(\Add0~35 ));
// synopsys translate_off
defparam \Add0~34 .lut_mask = 16'h9617;
defparam \Add0~34 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X50_Y35_N8
cycloneive_lcell_comb \Selector14~2 (
// Equation(s):
// \Selector14~2_combout  = (\Selector14~1_combout ) # ((\Selector0~13_combout  & (\porta~118_combout  $ (\portb~32_combout ))))

	.dataa(\Selector14~1_combout ),
	.datab(\Selector0~13_combout ),
	.datac(porta34),
	.datad(portb14),
	.cin(gnd),
	.combout(\Selector14~2_combout ),
	.cout());
// synopsys translate_off
defparam \Selector14~2 .lut_mask = 16'hAEEA;
defparam \Selector14~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X52_Y35_N2
cycloneive_lcell_comb \Selector14~0 (
// Equation(s):
// \Selector14~0_combout  = (\portb~32_combout  & ((\Selector0~10_combout ) # ((\porta~118_combout  & \Selector0~11_combout ))))

	.dataa(\Selector0~10_combout ),
	.datab(porta34),
	.datac(\Selector0~11_combout ),
	.datad(portb14),
	.cin(gnd),
	.combout(\Selector14~0_combout ),
	.cout());
// synopsys translate_off
defparam \Selector14~0 .lut_mask = 16'hEA00;
defparam \Selector14~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y42_N8
cycloneive_lcell_comb \Selector0~19 (
// Equation(s):
// \Selector0~19_combout  = (\Selector0~16_combout  & (!plif_idexaluop_l_3 & (\Selector0~15_combout  & !plif_idexaluop_l_0)))

	.dataa(\Selector0~16_combout ),
	.datab(plif_idexaluop_l_3),
	.datac(\Selector0~15_combout ),
	.datad(plif_idexaluop_l_0),
	.cin(gnd),
	.combout(\Selector0~19_combout ),
	.cout());
// synopsys translate_off
defparam \Selector0~19 .lut_mask = 16'h0020;
defparam \Selector0~19 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y41_N22
cycloneive_lcell_comb \Selector14~3 (
// Equation(s):
// \Selector14~3_combout  = (\Selector0~19_combout  & ((\portb~62_combout  & (\ShiftLeft0~8_combout )) # (!\portb~62_combout  & ((\ShiftLeft0~24_combout )))))

	.dataa(\ShiftLeft0~8_combout ),
	.datab(portb29),
	.datac(\Selector0~19_combout ),
	.datad(\ShiftLeft0~24_combout ),
	.cin(gnd),
	.combout(\Selector14~3_combout ),
	.cout());
// synopsys translate_off
defparam \Selector14~3 .lut_mask = 16'hB080;
defparam \Selector14~3 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X52_Y42_N30
cycloneive_lcell_comb \Selector0~21 (
// Equation(s):
// \Selector0~21_combout  = (\Selector0~15_combout  & (!plif_idexaluop_l_0 & !\Selector1~2_combout ))

	.dataa(\Selector0~15_combout ),
	.datab(plif_idexaluop_l_0),
	.datac(\Selector1~2_combout ),
	.datad(gnd),
	.cin(gnd),
	.combout(\Selector0~21_combout ),
	.cout());
// synopsys translate_off
defparam \Selector0~21 .lut_mask = 16'h0202;
defparam \Selector0~21 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y40_N4
cycloneive_lcell_comb \ShiftLeft0~48 (
// Equation(s):
// \ShiftLeft0~48_combout  = (\portb~58_combout  & ((\porta~96_combout ))) # (!\portb~58_combout  & (\porta~118_combout ))

	.dataa(gnd),
	.datab(portb27),
	.datac(porta34),
	.datad(porta12),
	.cin(gnd),
	.combout(\ShiftLeft0~48_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftLeft0~48 .lut_mask = 16'hFC30;
defparam \ShiftLeft0~48 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y36_N26
cycloneive_lcell_comb \ShiftLeft0~49 (
// Equation(s):
// \ShiftLeft0~49_combout  = (\portb~60_combout  & ((\ShiftLeft0~42_combout ))) # (!\portb~60_combout  & (\ShiftLeft0~48_combout ))

	.dataa(portb28),
	.datab(gnd),
	.datac(\ShiftLeft0~48_combout ),
	.datad(\ShiftLeft0~42_combout ),
	.cin(gnd),
	.combout(\ShiftLeft0~49_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftLeft0~49 .lut_mask = 16'hFA50;
defparam \ShiftLeft0~49 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X50_Y38_N20
cycloneive_lcell_comb \ShiftLeft0~50 (
// Equation(s):
// \ShiftLeft0~50_combout  = (\portb~62_combout  & (\ShiftLeft0~38_combout )) # (!\portb~62_combout  & ((\ShiftLeft0~49_combout )))

	.dataa(portb29),
	.datab(gnd),
	.datac(\ShiftLeft0~38_combout ),
	.datad(\ShiftLeft0~49_combout ),
	.cin(gnd),
	.combout(\ShiftLeft0~50_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftLeft0~50 .lut_mask = 16'hF5A0;
defparam \ShiftLeft0~50 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y41_N18
cycloneive_lcell_comb \Selector14~4 (
// Equation(s):
// \Selector14~4_combout  = (\Selector8~1_combout  & ((\ShiftRight0~39_combout ) # ((\Selector0~21_combout  & \ShiftLeft0~50_combout )))) # (!\Selector8~1_combout  & (((\Selector0~21_combout  & \ShiftLeft0~50_combout ))))

	.dataa(\Selector8~1_combout ),
	.datab(\ShiftRight0~39_combout ),
	.datac(\Selector0~21_combout ),
	.datad(\ShiftLeft0~50_combout ),
	.cin(gnd),
	.combout(\Selector14~4_combout ),
	.cout());
// synopsys translate_off
defparam \Selector14~4 .lut_mask = 16'hF888;
defparam \Selector14~4 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y41_N16
cycloneive_lcell_comb \Selector14~5 (
// Equation(s):
// \Selector14~5_combout  = (\Selector14~2_combout ) # ((\Selector14~0_combout ) # ((\Selector14~3_combout ) # (\Selector14~4_combout )))

	.dataa(\Selector14~2_combout ),
	.datab(\Selector14~0_combout ),
	.datac(\Selector14~3_combout ),
	.datad(\Selector14~4_combout ),
	.cin(gnd),
	.combout(\Selector14~5_combout ),
	.cout());
// synopsys translate_off
defparam \Selector14~5 .lut_mask = 16'hFFFE;
defparam \Selector14~5 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X50_Y35_N14
cycloneive_lcell_comb \Selector0~20 (
// Equation(s):
// \Selector0~20_combout  = (!plif_idexaluop_l_2 & (!plif_idexaluop_l_3 & (!plif_idexaluop_l_1 & plif_idexaluop_l_0)))

	.dataa(plif_idexaluop_l_2),
	.datab(plif_idexaluop_l_3),
	.datac(plif_idexaluop_l_1),
	.datad(plif_idexaluop_l_0),
	.cin(gnd),
	.combout(\Selector0~20_combout ),
	.cout());
// synopsys translate_off
defparam \Selector0~20 .lut_mask = 16'h0100;
defparam \Selector0~20 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y38_N30
cycloneive_lcell_comb \Selector8~1 (
// Equation(s):
// \Selector8~1_combout  = (\Selector0~20_combout  & (!\portb~66_combout  & (!\ShiftRight0~41_combout  & !\ShiftRight0~8_combout )))

	.dataa(\Selector0~20_combout ),
	.datab(portb31),
	.datac(\ShiftRight0~41_combout ),
	.datad(\ShiftRight0~8_combout ),
	.cin(gnd),
	.combout(\Selector8~1_combout ),
	.cout());
// synopsys translate_off
defparam \Selector8~1 .lut_mask = 16'h0002;
defparam \Selector8~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X52_Y35_N8
cycloneive_lcell_comb \Selector15~0 (
// Equation(s):
// \Selector15~0_combout  = (\Selector0~19_combout  & ((\portb~62_combout  & ((\ShiftLeft0~13_combout ))) # (!\portb~62_combout  & (\ShiftLeft0~28_combout ))))

	.dataa(\ShiftLeft0~28_combout ),
	.datab(portb29),
	.datac(\ShiftLeft0~13_combout ),
	.datad(\Selector0~19_combout ),
	.cin(gnd),
	.combout(\Selector15~0_combout ),
	.cout());
// synopsys translate_off
defparam \Selector15~0 .lut_mask = 16'hE200;
defparam \Selector15~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y35_N4
cycloneive_lcell_comb \Selector15~3 (
// Equation(s):
// \Selector15~3_combout  = (\porta~96_combout  & (\Selector0~13_combout  & ((!\portb~34_combout )))) # (!\porta~96_combout  & ((\portb~34_combout  & (\Selector0~13_combout )) # (!\portb~34_combout  & ((\Selector0~12_combout )))))

	.dataa(porta12),
	.datab(\Selector0~13_combout ),
	.datac(\Selector0~12_combout ),
	.datad(portb15),
	.cin(gnd),
	.combout(\Selector15~3_combout ),
	.cout());
// synopsys translate_off
defparam \Selector15~3 .lut_mask = 16'h44D8;
defparam \Selector15~3 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y41_N30
cycloneive_lcell_comb \ShiftLeft0~45 (
// Equation(s):
// \ShiftLeft0~45_combout  = (\portb~58_combout  & (\porta~99_combout )) # (!\portb~58_combout  & ((\porta~98_combout )))

	.dataa(porta15),
	.datab(porta14),
	.datac(portb27),
	.datad(gnd),
	.cin(gnd),
	.combout(\ShiftLeft0~45_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftLeft0~45 .lut_mask = 16'hACAC;
defparam \ShiftLeft0~45 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y40_N16
cycloneive_lcell_comb \ShiftLeft0~51 (
// Equation(s):
// \ShiftLeft0~51_combout  = (\portb~58_combout  & (\porta~97_combout )) # (!\portb~58_combout  & ((\porta~96_combout )))

	.dataa(porta13),
	.datab(gnd),
	.datac(portb27),
	.datad(porta12),
	.cin(gnd),
	.combout(\ShiftLeft0~51_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftLeft0~51 .lut_mask = 16'hAFA0;
defparam \ShiftLeft0~51 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y40_N26
cycloneive_lcell_comb \ShiftLeft0~52 (
// Equation(s):
// \ShiftLeft0~52_combout  = (\portb~60_combout  & (\ShiftLeft0~45_combout )) # (!\portb~60_combout  & ((\ShiftLeft0~51_combout )))

	.dataa(portb28),
	.datab(gnd),
	.datac(\ShiftLeft0~45_combout ),
	.datad(\ShiftLeft0~51_combout ),
	.cin(gnd),
	.combout(\ShiftLeft0~52_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftLeft0~52 .lut_mask = 16'hF5A0;
defparam \ShiftLeft0~52 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y40_N18
cycloneive_lcell_comb \ShiftLeft0~53 (
// Equation(s):
// \ShiftLeft0~53_combout  = (\portb~62_combout  & ((\ShiftLeft0~41_combout ))) # (!\portb~62_combout  & (\ShiftLeft0~52_combout ))

	.dataa(gnd),
	.datab(portb29),
	.datac(\ShiftLeft0~52_combout ),
	.datad(\ShiftLeft0~41_combout ),
	.cin(gnd),
	.combout(\ShiftLeft0~53_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftLeft0~53 .lut_mask = 16'hFC30;
defparam \ShiftLeft0~53 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y37_N16
cycloneive_lcell_comb \Selector15~1 (
// Equation(s):
// \Selector15~1_combout  = (!plif_idexaluop_l_0 & (\Selector0~15_combout  & (\ShiftLeft0~53_combout  & !\Selector1~2_combout )))

	.dataa(plif_idexaluop_l_0),
	.datab(\Selector0~15_combout ),
	.datac(\ShiftLeft0~53_combout ),
	.datad(\Selector1~2_combout ),
	.cin(gnd),
	.combout(\Selector15~1_combout ),
	.cout());
// synopsys translate_off
defparam \Selector15~1 .lut_mask = 16'h0040;
defparam \Selector15~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y37_N6
cycloneive_lcell_comb \Selector15~2 (
// Equation(s):
// \Selector15~2_combout  = (\Selector15~1_combout ) # ((\porta~91_combout  & (\Selector1~4_combout  & !\ShiftRight0~71_combout )))

	.dataa(porta7),
	.datab(\Selector1~4_combout ),
	.datac(\ShiftRight0~71_combout ),
	.datad(\Selector15~1_combout ),
	.cin(gnd),
	.combout(\Selector15~2_combout ),
	.cout());
// synopsys translate_off
defparam \Selector15~2 .lut_mask = 16'hFF08;
defparam \Selector15~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y37_N4
cycloneive_lcell_comb \Selector15~4 (
// Equation(s):
// \Selector15~4_combout  = (\Selector15~3_combout ) # ((\Selector15~2_combout ) # ((\porta~96_combout  & \Selector0~10_combout )))

	.dataa(porta12),
	.datab(\Selector0~10_combout ),
	.datac(\Selector15~3_combout ),
	.datad(\Selector15~2_combout ),
	.cin(gnd),
	.combout(\Selector15~4_combout ),
	.cout());
// synopsys translate_off
defparam \Selector15~4 .lut_mask = 16'hFFF8;
defparam \Selector15~4 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X50_Y36_N12
cycloneive_lcell_comb \Selector15~5 (
// Equation(s):
// \Selector15~5_combout  = (\portb~34_combout  & ((\Selector0~10_combout ) # ((\porta~96_combout  & \Selector0~11_combout ))))

	.dataa(\Selector0~10_combout ),
	.datab(porta12),
	.datac(\Selector0~11_combout ),
	.datad(portb15),
	.cin(gnd),
	.combout(\Selector15~5_combout ),
	.cout());
// synopsys translate_off
defparam \Selector15~5 .lut_mask = 16'hEA00;
defparam \Selector15~5 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X50_Y37_N26
cycloneive_lcell_comb \Selector15~6 (
// Equation(s):
// \Selector15~6_combout  = (\Selector15~5_combout ) # ((\Selector0~9_combout  & \Add0~32_combout ))

	.dataa(gnd),
	.datab(\Selector0~9_combout ),
	.datac(\Add0~32_combout ),
	.datad(\Selector15~5_combout ),
	.cin(gnd),
	.combout(\Selector15~6_combout ),
	.cout());
// synopsys translate_off
defparam \Selector15~6 .lut_mask = 16'hFFC0;
defparam \Selector15~6 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y37_N2
cycloneive_lcell_comb \Selector15~7 (
// Equation(s):
// \Selector15~7_combout  = (\Selector15~4_combout ) # ((\Selector15~6_combout ) # ((\Selector0~8_combout  & \Add1~32_combout )))

	.dataa(\Selector0~8_combout ),
	.datab(\Add1~32_combout ),
	.datac(\Selector15~4_combout ),
	.datad(\Selector15~6_combout ),
	.cin(gnd),
	.combout(\Selector15~7_combout ),
	.cout());
// synopsys translate_off
defparam \Selector15~7 .lut_mask = 16'hFFF8;
defparam \Selector15~7 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X52_Y37_N4
cycloneive_lcell_comb \Add0~36 (
// Equation(s):
// \Add0~36_combout  = ((\porta~117_combout  $ (\portb~30_combout  $ (!\Add0~35 )))) # (GND)
// \Add0~37  = CARRY((\porta~117_combout  & ((\portb~30_combout ) # (!\Add0~35 ))) # (!\porta~117_combout  & (\portb~30_combout  & !\Add0~35 )))

	.dataa(porta33),
	.datab(portb13),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add0~35 ),
	.combout(\Add0~36_combout ),
	.cout(\Add0~37 ));
// synopsys translate_off
defparam \Add0~36 .lut_mask = 16'h698E;
defparam \Add0~36 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X52_Y37_N6
cycloneive_lcell_comb \Add0~38 (
// Equation(s):
// \Add0~38_combout  = (\porta~116_combout  & ((\portb~28_combout  & (\Add0~37  & VCC)) # (!\portb~28_combout  & (!\Add0~37 )))) # (!\porta~116_combout  & ((\portb~28_combout  & (!\Add0~37 )) # (!\portb~28_combout  & ((\Add0~37 ) # (GND)))))
// \Add0~39  = CARRY((\porta~116_combout  & (!\portb~28_combout  & !\Add0~37 )) # (!\porta~116_combout  & ((!\Add0~37 ) # (!\portb~28_combout ))))

	.dataa(porta32),
	.datab(portb12),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add0~37 ),
	.combout(\Add0~38_combout ),
	.cout(\Add0~39 ));
// synopsys translate_off
defparam \Add0~38 .lut_mask = 16'h9617;
defparam \Add0~38 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X57_Y39_N4
cycloneive_lcell_comb \Add1~36 (
// Equation(s):
// \Add1~36_combout  = ((\portb~30_combout  $ (\porta~117_combout  $ (\Add1~35 )))) # (GND)
// \Add1~37  = CARRY((\portb~30_combout  & (\porta~117_combout  & !\Add1~35 )) # (!\portb~30_combout  & ((\porta~117_combout ) # (!\Add1~35 ))))

	.dataa(portb13),
	.datab(porta33),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add1~35 ),
	.combout(\Add1~36_combout ),
	.cout(\Add1~37 ));
// synopsys translate_off
defparam \Add1~36 .lut_mask = 16'h964D;
defparam \Add1~36 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X57_Y39_N6
cycloneive_lcell_comb \Add1~38 (
// Equation(s):
// \Add1~38_combout  = (\porta~116_combout  & ((\portb~28_combout  & (!\Add1~37 )) # (!\portb~28_combout  & (\Add1~37  & VCC)))) # (!\porta~116_combout  & ((\portb~28_combout  & ((\Add1~37 ) # (GND))) # (!\portb~28_combout  & (!\Add1~37 ))))
// \Add1~39  = CARRY((\porta~116_combout  & (\portb~28_combout  & !\Add1~37 )) # (!\porta~116_combout  & ((\portb~28_combout ) # (!\Add1~37 ))))

	.dataa(porta32),
	.datab(portb12),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add1~37 ),
	.combout(\Add1~38_combout ),
	.cout(\Add1~39 ));
// synopsys translate_off
defparam \Add1~38 .lut_mask = 16'h694D;
defparam \Add1~38 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X53_Y37_N30
cycloneive_lcell_comb \Selector12~9 (
// Equation(s):
// \Selector12~9_combout  = (\Selector0~9_combout  & ((\Add0~38_combout ) # ((\Selector0~8_combout  & \Add1~38_combout )))) # (!\Selector0~9_combout  & (\Selector0~8_combout  & ((\Add1~38_combout ))))

	.dataa(\Selector0~9_combout ),
	.datab(\Selector0~8_combout ),
	.datac(\Add0~38_combout ),
	.datad(\Add1~38_combout ),
	.cin(gnd),
	.combout(\Selector12~9_combout ),
	.cout());
// synopsys translate_off
defparam \Selector12~9 .lut_mask = 16'hECA0;
defparam \Selector12~9 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y37_N18
cycloneive_lcell_comb \Selector12~2 (
// Equation(s):
// \Selector12~2_combout  = (\Selector8~1_combout  & ((\portb~64_combout  & ((\ShiftRight0~81_combout ))) # (!\portb~64_combout  & (\Selector20~0_combout ))))

	.dataa(\Selector8~1_combout ),
	.datab(portb30),
	.datac(\Selector20~0_combout ),
	.datad(\ShiftRight0~81_combout ),
	.cin(gnd),
	.combout(\Selector12~2_combout ),
	.cout());
// synopsys translate_off
defparam \Selector12~2 .lut_mask = 16'hA820;
defparam \Selector12~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X50_Y40_N18
cycloneive_lcell_comb \Selector12~5 (
// Equation(s):
// \Selector12~5_combout  = (\porta~116_combout  & (((\Selector0~10_combout )))) # (!\porta~116_combout  & (!\portb~28_combout  & (\Selector0~12_combout )))

	.dataa(portb12),
	.datab(\Selector0~12_combout ),
	.datac(porta32),
	.datad(\Selector0~10_combout ),
	.cin(gnd),
	.combout(\Selector12~5_combout ),
	.cout());
// synopsys translate_off
defparam \Selector12~5 .lut_mask = 16'hF404;
defparam \Selector12~5 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X50_Y40_N12
cycloneive_lcell_comb \Selector12~6 (
// Equation(s):
// \Selector12~6_combout  = (\Selector12~5_combout ) # ((\Selector0~13_combout  & (\portb~28_combout  $ (\porta~116_combout ))))

	.dataa(portb12),
	.datab(\Selector0~13_combout ),
	.datac(porta32),
	.datad(\Selector12~5_combout ),
	.cin(gnd),
	.combout(\Selector12~6_combout ),
	.cout());
// synopsys translate_off
defparam \Selector12~6 .lut_mask = 16'hFF48;
defparam \Selector12~6 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X50_Y36_N30
cycloneive_lcell_comb \Selector12~4 (
// Equation(s):
// \Selector12~4_combout  = (\portb~28_combout  & ((\Selector0~10_combout ) # ((\Selector0~11_combout  & \porta~116_combout ))))

	.dataa(\Selector0~11_combout ),
	.datab(porta32),
	.datac(portb12),
	.datad(\Selector0~10_combout ),
	.cin(gnd),
	.combout(\Selector12~4_combout ),
	.cout());
// synopsys translate_off
defparam \Selector12~4 .lut_mask = 16'hF080;
defparam \Selector12~4 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y37_N26
cycloneive_lcell_comb \Selector12~12 (
// Equation(s):
// \Selector12~12_combout  = (!\portb~62_combout  & (\Selector1~4_combout  & (!\portb~64_combout  & \ShiftLeft0~4_combout )))

	.dataa(portb29),
	.datab(\Selector1~4_combout ),
	.datac(portb30),
	.datad(\ShiftLeft0~4_combout ),
	.cin(gnd),
	.combout(\Selector12~12_combout ),
	.cout());
// synopsys translate_off
defparam \Selector12~12 .lut_mask = 16'h0400;
defparam \Selector12~12 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y36_N4
cycloneive_lcell_comb \ShiftLeft0~54 (
// Equation(s):
// \ShiftLeft0~54_combout  = (\portb~58_combout  & ((\porta~117_combout ))) # (!\portb~58_combout  & (\porta~116_combout ))

	.dataa(porta32),
	.datab(gnd),
	.datac(porta33),
	.datad(portb27),
	.cin(gnd),
	.combout(\ShiftLeft0~54_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftLeft0~54 .lut_mask = 16'hF0AA;
defparam \ShiftLeft0~54 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X52_Y36_N28
cycloneive_lcell_comb \ShiftLeft0~55 (
// Equation(s):
// \ShiftLeft0~55_combout  = (\portb~60_combout  & ((\ShiftLeft0~48_combout ))) # (!\portb~60_combout  & (\ShiftLeft0~54_combout ))

	.dataa(gnd),
	.datab(\ShiftLeft0~54_combout ),
	.datac(portb28),
	.datad(\ShiftLeft0~48_combout ),
	.cin(gnd),
	.combout(\ShiftLeft0~55_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftLeft0~55 .lut_mask = 16'hFC0C;
defparam \ShiftLeft0~55 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X52_Y36_N10
cycloneive_lcell_comb \ShiftLeft0~56 (
// Equation(s):
// \ShiftLeft0~56_combout  = (\portb~62_combout  & (\ShiftLeft0~43_combout )) # (!\portb~62_combout  & ((\ShiftLeft0~55_combout )))

	.dataa(portb29),
	.datab(gnd),
	.datac(\ShiftLeft0~43_combout ),
	.datad(\ShiftLeft0~55_combout ),
	.cin(gnd),
	.combout(\ShiftLeft0~56_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftLeft0~56 .lut_mask = 16'hF5A0;
defparam \ShiftLeft0~56 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y37_N24
cycloneive_lcell_comb \Selector12~3 (
// Equation(s):
// \Selector12~3_combout  = (!plif_idexaluop_l_0 & (\Selector0~15_combout  & (\ShiftLeft0~56_combout  & !\Selector1~2_combout )))

	.dataa(plif_idexaluop_l_0),
	.datab(\Selector0~15_combout ),
	.datac(\ShiftLeft0~56_combout ),
	.datad(\Selector1~2_combout ),
	.cin(gnd),
	.combout(\Selector12~3_combout ),
	.cout());
// synopsys translate_off
defparam \Selector12~3 .lut_mask = 16'h0040;
defparam \Selector12~3 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y37_N14
cycloneive_lcell_comb \Selector12~7 (
// Equation(s):
// \Selector12~7_combout  = (\Selector12~6_combout ) # ((\Selector12~4_combout ) # ((\Selector12~12_combout ) # (\Selector12~3_combout )))

	.dataa(\Selector12~6_combout ),
	.datab(\Selector12~4_combout ),
	.datac(\Selector12~12_combout ),
	.datad(\Selector12~3_combout ),
	.cin(gnd),
	.combout(\Selector12~7_combout ),
	.cout());
// synopsys translate_off
defparam \Selector12~7 .lut_mask = 16'hFFFE;
defparam \Selector12~7 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y37_N12
cycloneive_lcell_comb \Selector12~8 (
// Equation(s):
// \Selector12~8_combout  = (\Selector0~19_combout  & ((\portb~62_combout  & ((\ShiftLeft0~16_combout ))) # (!\portb~62_combout  & (\ShiftLeft0~30_combout ))))

	.dataa(\ShiftLeft0~30_combout ),
	.datab(\ShiftLeft0~16_combout ),
	.datac(portb29),
	.datad(\Selector0~19_combout ),
	.cin(gnd),
	.combout(\Selector12~8_combout ),
	.cout());
// synopsys translate_off
defparam \Selector12~8 .lut_mask = 16'hCA00;
defparam \Selector12~8 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y37_N4
cycloneive_lcell_comb \Selector13~1 (
// Equation(s):
// \Selector13~1_combout  = (\ShiftLeft0~59_combout  & (\Selector0~15_combout  & (!plif_idexaluop_l_0 & !\Selector1~2_combout )))

	.dataa(\ShiftLeft0~59_combout ),
	.datab(\Selector0~15_combout ),
	.datac(plif_idexaluop_l_0),
	.datad(\Selector1~2_combout ),
	.cin(gnd),
	.combout(\Selector13~1_combout ),
	.cout());
// synopsys translate_off
defparam \Selector13~1 .lut_mask = 16'h0008;
defparam \Selector13~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y37_N24
cycloneive_lcell_comb \Selector13~2 (
// Equation(s):
// \Selector13~2_combout  = (\porta~117_combout  & (((\Selector0~10_combout )))) # (!\porta~117_combout  & (\Selector0~12_combout  & ((!\portb~30_combout ))))

	.dataa(\Selector0~12_combout ),
	.datab(\Selector0~10_combout ),
	.datac(porta33),
	.datad(portb13),
	.cin(gnd),
	.combout(\Selector13~2_combout ),
	.cout());
// synopsys translate_off
defparam \Selector13~2 .lut_mask = 16'hC0CA;
defparam \Selector13~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y37_N26
cycloneive_lcell_comb \Selector13~3 (
// Equation(s):
// \Selector13~3_combout  = (\Selector13~2_combout ) # ((\Selector0~13_combout  & (\portb~30_combout  $ (\porta~117_combout ))))

	.dataa(\Selector0~13_combout ),
	.datab(portb13),
	.datac(porta33),
	.datad(\Selector13~2_combout ),
	.cin(gnd),
	.combout(\Selector13~3_combout ),
	.cout());
// synopsys translate_off
defparam \Selector13~3 .lut_mask = 16'hFF28;
defparam \Selector13~3 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y38_N30
cycloneive_lcell_comb \Selector12~11 (
// Equation(s):
// \Selector12~11_combout  = (\ShiftRight0~74_combout  & (\portb~66_combout  & (!plif_idexaluop_l_0 & \Selector1~3_combout )))

	.dataa(\ShiftRight0~74_combout ),
	.datab(portb31),
	.datac(plif_idexaluop_l_0),
	.datad(\Selector1~3_combout ),
	.cin(gnd),
	.combout(\Selector12~11_combout ),
	.cout());
// synopsys translate_off
defparam \Selector12~11 .lut_mask = 16'h0800;
defparam \Selector12~11 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y37_N0
cycloneive_lcell_comb \Selector13~5 (
// Equation(s):
// \Selector13~5_combout  = (\Selector8~1_combout  & ((\ShiftRight0~93_combout ) # ((\ShiftLeft0~6_combout  & \Selector12~11_combout )))) # (!\Selector8~1_combout  & (\ShiftLeft0~6_combout  & (\Selector12~11_combout )))

	.dataa(\Selector8~1_combout ),
	.datab(\ShiftLeft0~6_combout ),
	.datac(\Selector12~11_combout ),
	.datad(\ShiftRight0~93_combout ),
	.cin(gnd),
	.combout(\Selector13~5_combout ),
	.cout());
// synopsys translate_off
defparam \Selector13~5 .lut_mask = 16'hEAC0;
defparam \Selector13~5 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y37_N16
cycloneive_lcell_comb \Selector13~6 (
// Equation(s):
// \Selector13~6_combout  = (\Selector13~3_combout ) # ((\Selector13~5_combout ) # ((\Selector13~4_combout  & \portb~30_combout )))

	.dataa(\Selector13~4_combout ),
	.datab(portb13),
	.datac(\Selector13~3_combout ),
	.datad(\Selector13~5_combout ),
	.cin(gnd),
	.combout(\Selector13~6_combout ),
	.cout());
// synopsys translate_off
defparam \Selector13~6 .lut_mask = 16'hFFF8;
defparam \Selector13~6 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y37_N30
cycloneive_lcell_comb \Selector13~7 (
// Equation(s):
// \Selector13~7_combout  = (\Selector13~1_combout ) # ((\Selector13~6_combout ) # ((\Add0~36_combout  & \Selector0~9_combout )))

	.dataa(\Add0~36_combout ),
	.datab(\Selector0~9_combout ),
	.datac(\Selector13~1_combout ),
	.datad(\Selector13~6_combout ),
	.cin(gnd),
	.combout(\Selector13~7_combout ),
	.cout());
// synopsys translate_off
defparam \Selector13~7 .lut_mask = 16'hFFF8;
defparam \Selector13~7 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y41_N6
cycloneive_lcell_comb \Selector13~0 (
// Equation(s):
// \Selector13~0_combout  = (\Selector0~19_combout  & ((\portb~62_combout  & (\ShiftLeft0~19_combout )) # (!\portb~62_combout  & ((\ShiftLeft0~34_combout )))))

	.dataa(\ShiftLeft0~19_combout ),
	.datab(\Selector0~19_combout ),
	.datac(\ShiftLeft0~34_combout ),
	.datad(portb29),
	.cin(gnd),
	.combout(\Selector13~0_combout ),
	.cout());
// synopsys translate_off
defparam \Selector13~0 .lut_mask = 16'h88C0;
defparam \Selector13~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y38_N14
cycloneive_lcell_comb \Selector10~1 (
// Equation(s):
// \Selector10~1_combout  = (\portb~24_combout  & ((\Selector0~10_combout ) # ((\porta~114_combout  & \Selector0~11_combout ))))

	.dataa(porta30),
	.datab(portb10),
	.datac(\Selector0~10_combout ),
	.datad(\Selector0~11_combout ),
	.cin(gnd),
	.combout(\Selector10~1_combout ),
	.cout());
// synopsys translate_off
defparam \Selector10~1 .lut_mask = 16'hC8C0;
defparam \Selector10~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X52_Y37_N8
cycloneive_lcell_comb \Add0~40 (
// Equation(s):
// \Add0~40_combout  = ((\portb~26_combout  $ (\porta~115_combout  $ (!\Add0~39 )))) # (GND)
// \Add0~41  = CARRY((\portb~26_combout  & ((\porta~115_combout ) # (!\Add0~39 ))) # (!\portb~26_combout  & (\porta~115_combout  & !\Add0~39 )))

	.dataa(portb11),
	.datab(porta31),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add0~39 ),
	.combout(\Add0~40_combout ),
	.cout(\Add0~41 ));
// synopsys translate_off
defparam \Add0~40 .lut_mask = 16'h698E;
defparam \Add0~40 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X52_Y37_N10
cycloneive_lcell_comb \Add0~42 (
// Equation(s):
// \Add0~42_combout  = (\porta~114_combout  & ((\portb~24_combout  & (\Add0~41  & VCC)) # (!\portb~24_combout  & (!\Add0~41 )))) # (!\porta~114_combout  & ((\portb~24_combout  & (!\Add0~41 )) # (!\portb~24_combout  & ((\Add0~41 ) # (GND)))))
// \Add0~43  = CARRY((\porta~114_combout  & (!\portb~24_combout  & !\Add0~41 )) # (!\porta~114_combout  & ((!\Add0~41 ) # (!\portb~24_combout ))))

	.dataa(porta30),
	.datab(portb10),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add0~41 ),
	.combout(\Add0~42_combout ),
	.cout(\Add0~43 ));
// synopsys translate_off
defparam \Add0~42 .lut_mask = 16'h9617;
defparam \Add0~42 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X59_Y38_N4
cycloneive_lcell_comb \Selector10~5 (
// Equation(s):
// \Selector10~5_combout  = (\porta~114_combout  & (((\Selector0~10_combout )))) # (!\porta~114_combout  & (!\portb~24_combout  & ((\Selector0~12_combout ))))

	.dataa(porta30),
	.datab(portb10),
	.datac(\Selector0~10_combout ),
	.datad(\Selector0~12_combout ),
	.cin(gnd),
	.combout(\Selector10~5_combout ),
	.cout());
// synopsys translate_off
defparam \Selector10~5 .lut_mask = 16'hB1A0;
defparam \Selector10~5 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y38_N26
cycloneive_lcell_comb \Selector10~6 (
// Equation(s):
// \Selector10~6_combout  = (\Selector10~5_combout ) # ((\Selector0~13_combout  & (\porta~114_combout  $ (\portb~24_combout ))))

	.dataa(porta30),
	.datab(portb10),
	.datac(\Selector10~5_combout ),
	.datad(\Selector0~13_combout ),
	.cin(gnd),
	.combout(\Selector10~6_combout ),
	.cout());
// synopsys translate_off
defparam \Selector10~6 .lut_mask = 16'hF6F0;
defparam \Selector10~6 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y39_N8
cycloneive_lcell_comb \Add1~40 (
// Equation(s):
// \Add1~40_combout  = ((\porta~115_combout  $ (\portb~26_combout  $ (\Add1~39 )))) # (GND)
// \Add1~41  = CARRY((\porta~115_combout  & ((!\Add1~39 ) # (!\portb~26_combout ))) # (!\porta~115_combout  & (!\portb~26_combout  & !\Add1~39 )))

	.dataa(porta31),
	.datab(portb11),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add1~39 ),
	.combout(\Add1~40_combout ),
	.cout(\Add1~41 ));
// synopsys translate_off
defparam \Add1~40 .lut_mask = 16'h962B;
defparam \Add1~40 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X57_Y39_N10
cycloneive_lcell_comb \Add1~42 (
// Equation(s):
// \Add1~42_combout  = (\porta~114_combout  & ((\portb~24_combout  & (!\Add1~41 )) # (!\portb~24_combout  & (\Add1~41  & VCC)))) # (!\porta~114_combout  & ((\portb~24_combout  & ((\Add1~41 ) # (GND))) # (!\portb~24_combout  & (!\Add1~41 ))))
// \Add1~43  = CARRY((\porta~114_combout  & (\portb~24_combout  & !\Add1~41 )) # (!\porta~114_combout  & ((\portb~24_combout ) # (!\Add1~41 ))))

	.dataa(porta30),
	.datab(portb10),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add1~41 ),
	.combout(\Add1~42_combout ),
	.cout(\Add1~43 ));
// synopsys translate_off
defparam \Add1~42 .lut_mask = 16'h694D;
defparam \Add1~42 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X54_Y42_N18
cycloneive_lcell_comb \Selector8~2 (
// Equation(s):
// \Selector8~2_combout  = (!\portb~64_combout  & (\portb~66_combout  & (!plif_idexaluop_l_0 & \Selector1~3_combout )))

	.dataa(portb30),
	.datab(portb31),
	.datac(plif_idexaluop_l_0),
	.datad(\Selector1~3_combout ),
	.cin(gnd),
	.combout(\Selector8~2_combout ),
	.cout());
// synopsys translate_off
defparam \Selector8~2 .lut_mask = 16'h0400;
defparam \Selector8~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y42_N14
cycloneive_lcell_comb \Selector10~3 (
// Equation(s):
// \Selector10~3_combout  = (\Selector8~1_combout  & ((\ShiftRight0~96_combout ) # ((\Selector0~19_combout  & \Selector10~0_combout )))) # (!\Selector8~1_combout  & (\Selector0~19_combout  & (\Selector10~0_combout )))

	.dataa(\Selector8~1_combout ),
	.datab(\Selector0~19_combout ),
	.datac(\Selector10~0_combout ),
	.datad(\ShiftRight0~96_combout ),
	.cin(gnd),
	.combout(\Selector10~3_combout ),
	.cout());
// synopsys translate_off
defparam \Selector10~3 .lut_mask = 16'hEAC0;
defparam \Selector10~3 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y36_N16
cycloneive_lcell_comb \ShiftLeft0~62 (
// Equation(s):
// \ShiftLeft0~62_combout  = (\portb~62_combout  & ((\ShiftLeft0~49_combout ))) # (!\portb~62_combout  & (\ShiftLeft0~61_combout ))

	.dataa(\ShiftLeft0~61_combout ),
	.datab(gnd),
	.datac(\ShiftLeft0~49_combout ),
	.datad(portb29),
	.cin(gnd),
	.combout(\ShiftLeft0~62_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftLeft0~62 .lut_mask = 16'hF0AA;
defparam \ShiftLeft0~62 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y42_N12
cycloneive_lcell_comb \Selector10~2 (
// Equation(s):
// \Selector10~2_combout  = (!plif_idexaluop_l_0 & (\ShiftLeft0~62_combout  & \Selector0~18_combout ))

	.dataa(gnd),
	.datab(plif_idexaluop_l_0),
	.datac(\ShiftLeft0~62_combout ),
	.datad(\Selector0~18_combout ),
	.cin(gnd),
	.combout(\Selector10~2_combout ),
	.cout());
// synopsys translate_off
defparam \Selector10~2 .lut_mask = 16'h3000;
defparam \Selector10~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y42_N24
cycloneive_lcell_comb \Selector10~4 (
// Equation(s):
// \Selector10~4_combout  = (\Selector10~3_combout ) # ((\Selector10~2_combout ) # ((\ShiftLeft0~9_combout  & \Selector8~2_combout )))

	.dataa(\ShiftLeft0~9_combout ),
	.datab(\Selector8~2_combout ),
	.datac(\Selector10~3_combout ),
	.datad(\Selector10~2_combout ),
	.cin(gnd),
	.combout(\Selector10~4_combout ),
	.cout());
// synopsys translate_off
defparam \Selector10~4 .lut_mask = 16'hFFF8;
defparam \Selector10~4 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y42_N2
cycloneive_lcell_comb \Selector10~7 (
// Equation(s):
// \Selector10~7_combout  = (\Selector10~6_combout ) # ((\Selector10~4_combout ) # ((\Selector0~8_combout  & \Add1~42_combout )))

	.dataa(\Selector0~8_combout ),
	.datab(\Selector10~6_combout ),
	.datac(\Add1~42_combout ),
	.datad(\Selector10~4_combout ),
	.cin(gnd),
	.combout(\Selector10~7_combout ),
	.cout());
// synopsys translate_off
defparam \Selector10~7 .lut_mask = 16'hFFEC;
defparam \Selector10~7 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y39_N0
cycloneive_lcell_comb \Selector11~4 (
// Equation(s):
// \Selector11~4_combout  = (\Selector0~13_combout  & (\portb~26_combout  $ (\porta~115_combout )))

	.dataa(gnd),
	.datab(\Selector0~13_combout ),
	.datac(portb11),
	.datad(porta31),
	.cin(gnd),
	.combout(\Selector11~4_combout ),
	.cout());
// synopsys translate_off
defparam \Selector11~4 .lut_mask = 16'h0CC0;
defparam \Selector11~4 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X50_Y41_N18
cycloneive_lcell_comb \Selector11~1 (
// Equation(s):
// \Selector11~1_combout  = (\porta~115_combout  & (((\Selector0~10_combout )))) # (!\porta~115_combout  & (\Selector0~12_combout  & ((!\portb~26_combout ))))

	.dataa(\Selector0~12_combout ),
	.datab(\Selector0~10_combout ),
	.datac(porta31),
	.datad(portb11),
	.cin(gnd),
	.combout(\Selector11~1_combout ),
	.cout());
// synopsys translate_off
defparam \Selector11~1 .lut_mask = 16'hC0CA;
defparam \Selector11~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y39_N18
cycloneive_lcell_comb \Selector11~3 (
// Equation(s):
// \Selector11~3_combout  = (\Selector11~2_combout ) # ((\Selector11~1_combout ) # ((\ShiftRight0~99_combout  & \Selector8~1_combout )))

	.dataa(\Selector11~2_combout ),
	.datab(\Selector11~1_combout ),
	.datac(\ShiftRight0~99_combout ),
	.datad(\Selector8~1_combout ),
	.cin(gnd),
	.combout(\Selector11~3_combout ),
	.cout());
// synopsys translate_off
defparam \Selector11~3 .lut_mask = 16'hFEEE;
defparam \Selector11~3 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y39_N26
cycloneive_lcell_comb \Selector11~5 (
// Equation(s):
// \Selector11~5_combout  = (\Selector11~4_combout ) # ((\Selector11~3_combout ) # ((\Add1~40_combout  & \Selector0~8_combout )))

	.dataa(\Add1~40_combout ),
	.datab(\Selector11~4_combout ),
	.datac(\Selector0~8_combout ),
	.datad(\Selector11~3_combout ),
	.cin(gnd),
	.combout(\Selector11~5_combout ),
	.cout());
// synopsys translate_off
defparam \Selector11~5 .lut_mask = 16'hFFEC;
defparam \Selector11~5 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y42_N4
cycloneive_lcell_comb \Selector11~7 (
// Equation(s):
// \Selector11~7_combout  = (\portb~26_combout  & ((\Selector0~10_combout ) # ((\Selector0~11_combout  & \porta~115_combout ))))

	.dataa(\Selector0~10_combout ),
	.datab(portb11),
	.datac(\Selector0~11_combout ),
	.datad(porta31),
	.cin(gnd),
	.combout(\Selector11~7_combout ),
	.cout());
// synopsys translate_off
defparam \Selector11~7 .lut_mask = 16'hC888;
defparam \Selector11~7 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y42_N6
cycloneive_lcell_comb \Selector11~6 (
// Equation(s):
// \Selector11~6_combout  = (\ShiftLeft0~14_combout  & ((\Selector8~2_combout ) # ((\Selector0~19_combout  & \Selector11~0_combout )))) # (!\ShiftLeft0~14_combout  & (\Selector0~19_combout  & (\Selector11~0_combout )))

	.dataa(\ShiftLeft0~14_combout ),
	.datab(\Selector0~19_combout ),
	.datac(\Selector11~0_combout ),
	.datad(\Selector8~2_combout ),
	.cin(gnd),
	.combout(\Selector11~6_combout ),
	.cout());
// synopsys translate_off
defparam \Selector11~6 .lut_mask = 16'hEAC0;
defparam \Selector11~6 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y42_N30
cycloneive_lcell_comb \Selector11~8 (
// Equation(s):
// \Selector11~8_combout  = (\Selector11~7_combout ) # (\Selector11~6_combout )

	.dataa(gnd),
	.datab(gnd),
	.datac(\Selector11~7_combout ),
	.datad(\Selector11~6_combout ),
	.cin(gnd),
	.combout(\Selector11~8_combout ),
	.cout());
// synopsys translate_off
defparam \Selector11~8 .lut_mask = 16'hFFF0;
defparam \Selector11~8 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X50_Y40_N0
cycloneive_lcell_comb \Selector8~7 (
// Equation(s):
// \Selector8~7_combout  = (\porta~112_combout  & ((\Selector0~10_combout ) # (!\portb~20_combout ))) # (!\porta~112_combout  & ((\portb~20_combout )))

	.dataa(gnd),
	.datab(porta28),
	.datac(\Selector0~10_combout ),
	.datad(portb8),
	.cin(gnd),
	.combout(\Selector8~7_combout ),
	.cout());
// synopsys translate_off
defparam \Selector8~7 .lut_mask = 16'hF3CC;
defparam \Selector8~7 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X50_Y40_N6
cycloneive_lcell_comb \Selector8~8 (
// Equation(s):
// \Selector8~8_combout  = (\Selector8~7_combout  & (((\Selector0~10_combout ) # (\Selector0~13_combout )))) # (!\Selector8~7_combout  & (\Selector8~6_combout ))

	.dataa(\Selector8~6_combout ),
	.datab(\Selector0~10_combout ),
	.datac(\Selector0~13_combout ),
	.datad(\Selector8~7_combout ),
	.cin(gnd),
	.combout(\Selector8~8_combout ),
	.cout());
// synopsys translate_off
defparam \Selector8~8 .lut_mask = 16'hFCAA;
defparam \Selector8~8 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X52_Y37_N12
cycloneive_lcell_comb \Add0~44 (
// Equation(s):
// \Add0~44_combout  = ((\portb~22_combout  $ (\porta~113_combout  $ (!\Add0~43 )))) # (GND)
// \Add0~45  = CARRY((\portb~22_combout  & ((\porta~113_combout ) # (!\Add0~43 ))) # (!\portb~22_combout  & (\porta~113_combout  & !\Add0~43 )))

	.dataa(portb9),
	.datab(porta29),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add0~43 ),
	.combout(\Add0~44_combout ),
	.cout(\Add0~45 ));
// synopsys translate_off
defparam \Add0~44 .lut_mask = 16'h698E;
defparam \Add0~44 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X52_Y37_N14
cycloneive_lcell_comb \Add0~46 (
// Equation(s):
// \Add0~46_combout  = (\portb~20_combout  & ((\porta~112_combout  & (\Add0~45  & VCC)) # (!\porta~112_combout  & (!\Add0~45 )))) # (!\portb~20_combout  & ((\porta~112_combout  & (!\Add0~45 )) # (!\porta~112_combout  & ((\Add0~45 ) # (GND)))))
// \Add0~47  = CARRY((\portb~20_combout  & (!\porta~112_combout  & !\Add0~45 )) # (!\portb~20_combout  & ((!\Add0~45 ) # (!\porta~112_combout ))))

	.dataa(portb8),
	.datab(porta28),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add0~45 ),
	.combout(\Add0~46_combout ),
	.cout(\Add0~47 ));
// synopsys translate_off
defparam \Add0~46 .lut_mask = 16'h9617;
defparam \Add0~46 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X52_Y39_N10
cycloneive_lcell_comb \Selector8~9 (
// Equation(s):
// \Selector8~9_combout  = (\Selector8~8_combout ) # ((\Selector0~9_combout  & \Add0~46_combout ))

	.dataa(\Selector0~9_combout ),
	.datab(\Selector8~8_combout ),
	.datac(gnd),
	.datad(\Add0~46_combout ),
	.cin(gnd),
	.combout(\Selector8~9_combout ),
	.cout());
// synopsys translate_off
defparam \Selector8~9 .lut_mask = 16'hEECC;
defparam \Selector8~9 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y39_N12
cycloneive_lcell_comb \Add1~44 (
// Equation(s):
// \Add1~44_combout  = ((\portb~22_combout  $ (\porta~113_combout  $ (\Add1~43 )))) # (GND)
// \Add1~45  = CARRY((\portb~22_combout  & (\porta~113_combout  & !\Add1~43 )) # (!\portb~22_combout  & ((\porta~113_combout ) # (!\Add1~43 ))))

	.dataa(portb9),
	.datab(porta29),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add1~43 ),
	.combout(\Add1~44_combout ),
	.cout(\Add1~45 ));
// synopsys translate_off
defparam \Add1~44 .lut_mask = 16'h964D;
defparam \Add1~44 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X57_Y39_N14
cycloneive_lcell_comb \Add1~46 (
// Equation(s):
// \Add1~46_combout  = (\portb~20_combout  & ((\porta~112_combout  & (!\Add1~45 )) # (!\porta~112_combout  & ((\Add1~45 ) # (GND))))) # (!\portb~20_combout  & ((\porta~112_combout  & (\Add1~45  & VCC)) # (!\porta~112_combout  & (!\Add1~45 ))))
// \Add1~47  = CARRY((\portb~20_combout  & ((!\Add1~45 ) # (!\porta~112_combout ))) # (!\portb~20_combout  & (!\porta~112_combout  & !\Add1~45 )))

	.dataa(portb8),
	.datab(porta28),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add1~45 ),
	.combout(\Add1~46_combout ),
	.cout(\Add1~47 ));
// synopsys translate_off
defparam \Add1~46 .lut_mask = 16'h692B;
defparam \Add1~46 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X53_Y36_N20
cycloneive_lcell_comb \ShiftLeft0~60 (
// Equation(s):
// \ShiftLeft0~60_combout  = (\portb~58_combout  & ((\porta~115_combout ))) # (!\portb~58_combout  & (\porta~114_combout ))

	.dataa(porta30),
	.datab(porta31),
	.datac(portb27),
	.datad(gnd),
	.cin(gnd),
	.combout(\ShiftLeft0~60_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftLeft0~60 .lut_mask = 16'hCACA;
defparam \ShiftLeft0~60 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y36_N10
cycloneive_lcell_comb \ShiftLeft0~66 (
// Equation(s):
// \ShiftLeft0~66_combout  = (\portb~58_combout  & (\porta~113_combout )) # (!\portb~58_combout  & ((\porta~112_combout )))

	.dataa(portb27),
	.datab(gnd),
	.datac(porta29),
	.datad(porta28),
	.cin(gnd),
	.combout(\ShiftLeft0~66_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftLeft0~66 .lut_mask = 16'hF5A0;
defparam \ShiftLeft0~66 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y36_N0
cycloneive_lcell_comb \ShiftLeft0~67 (
// Equation(s):
// \ShiftLeft0~67_combout  = (\portb~60_combout  & (\ShiftLeft0~60_combout )) # (!\portb~60_combout  & ((\ShiftLeft0~66_combout )))

	.dataa(gnd),
	.datab(\ShiftLeft0~60_combout ),
	.datac(portb28),
	.datad(\ShiftLeft0~66_combout ),
	.cin(gnd),
	.combout(\ShiftLeft0~67_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftLeft0~67 .lut_mask = 16'hCFC0;
defparam \ShiftLeft0~67 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X52_Y42_N0
cycloneive_lcell_comb \Selector8~3 (
// Equation(s):
// \Selector8~3_combout  = (\Selector0~21_combout  & ((\portb~62_combout  & ((\ShiftLeft0~55_combout ))) # (!\portb~62_combout  & (\ShiftLeft0~67_combout ))))

	.dataa(\Selector0~21_combout ),
	.datab(portb29),
	.datac(\ShiftLeft0~67_combout ),
	.datad(\ShiftLeft0~55_combout ),
	.cin(gnd),
	.combout(\Selector8~3_combout ),
	.cout());
// synopsys translate_off
defparam \Selector8~3 .lut_mask = 16'hA820;
defparam \Selector8~3 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y42_N6
cycloneive_lcell_comb \Selector8~4 (
// Equation(s):
// \Selector8~4_combout  = (\Selector8~1_combout  & ((\ShiftRight0~105_combout ) # ((\Selector8~2_combout  & \ShiftLeft0~17_combout )))) # (!\Selector8~1_combout  & (\Selector8~2_combout  & ((\ShiftLeft0~17_combout ))))

	.dataa(\Selector8~1_combout ),
	.datab(\Selector8~2_combout ),
	.datac(\ShiftRight0~105_combout ),
	.datad(\ShiftLeft0~17_combout ),
	.cin(gnd),
	.combout(\Selector8~4_combout ),
	.cout());
// synopsys translate_off
defparam \Selector8~4 .lut_mask = 16'hECA0;
defparam \Selector8~4 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y42_N16
cycloneive_lcell_comb \Selector8~5 (
// Equation(s):
// \Selector8~5_combout  = (\Selector8~3_combout ) # ((\Selector8~4_combout ) # ((\Selector0~19_combout  & \Selector8~0_combout )))

	.dataa(\Selector8~3_combout ),
	.datab(\Selector0~19_combout ),
	.datac(\Selector8~0_combout ),
	.datad(\Selector8~4_combout ),
	.cin(gnd),
	.combout(\Selector8~5_combout ),
	.cout());
// synopsys translate_off
defparam \Selector8~5 .lut_mask = 16'hFFEA;
defparam \Selector8~5 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y39_N24
cycloneive_lcell_comb \Selector9~1 (
// Equation(s):
// \Selector9~1_combout  = (\Selector8~1_combout  & ((\ShiftRight0~104_combout ) # ((\ShiftRight0~74_combout  & \ShiftRight0~91_combout ))))

	.dataa(\ShiftRight0~74_combout ),
	.datab(\ShiftRight0~91_combout ),
	.datac(\ShiftRight0~104_combout ),
	.datad(\Selector8~1_combout ),
	.cin(gnd),
	.combout(\Selector9~1_combout ),
	.cout());
// synopsys translate_off
defparam \Selector9~1 .lut_mask = 16'hF800;
defparam \Selector9~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y39_N26
cycloneive_lcell_comb \Selector9~2 (
// Equation(s):
// \Selector9~2_combout  = (\portb~22_combout  & ((\Selector0~10_combout ) # ((\Selector0~11_combout  & \porta~113_combout ))))

	.dataa(\Selector0~10_combout ),
	.datab(\Selector0~11_combout ),
	.datac(portb9),
	.datad(porta29),
	.cin(gnd),
	.combout(\Selector9~2_combout ),
	.cout());
// synopsys translate_off
defparam \Selector9~2 .lut_mask = 16'hE0A0;
defparam \Selector9~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y40_N10
cycloneive_lcell_comb \ShiftLeft0~57 (
// Equation(s):
// \ShiftLeft0~57_combout  = (\portb~58_combout  & (\porta~118_combout )) # (!\portb~58_combout  & ((\porta~117_combout )))

	.dataa(gnd),
	.datab(portb27),
	.datac(porta34),
	.datad(porta33),
	.cin(gnd),
	.combout(\ShiftLeft0~57_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftLeft0~57 .lut_mask = 16'hF3C0;
defparam \ShiftLeft0~57 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y40_N2
cycloneive_lcell_comb \ShiftLeft0~58 (
// Equation(s):
// \ShiftLeft0~58_combout  = (\portb~60_combout  & ((\ShiftLeft0~51_combout ))) # (!\portb~60_combout  & (\ShiftLeft0~57_combout ))

	.dataa(portb28),
	.datab(gnd),
	.datac(\ShiftLeft0~57_combout ),
	.datad(\ShiftLeft0~51_combout ),
	.cin(gnd),
	.combout(\ShiftLeft0~58_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftLeft0~58 .lut_mask = 16'hFA50;
defparam \ShiftLeft0~58 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X52_Y36_N24
cycloneive_lcell_comb \ShiftLeft0~68 (
// Equation(s):
// \ShiftLeft0~68_combout  = (\portb~58_combout  & (\porta~114_combout )) # (!\portb~58_combout  & ((\porta~113_combout )))

	.dataa(portb27),
	.datab(gnd),
	.datac(porta30),
	.datad(porta29),
	.cin(gnd),
	.combout(\ShiftLeft0~68_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftLeft0~68 .lut_mask = 16'hF5A0;
defparam \ShiftLeft0~68 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y40_N26
cycloneive_lcell_comb \ShiftLeft0~69 (
// Equation(s):
// \ShiftLeft0~69_combout  = (\portb~60_combout  & (\ShiftLeft0~63_combout )) # (!\portb~60_combout  & ((\ShiftLeft0~68_combout )))

	.dataa(\ShiftLeft0~63_combout ),
	.datab(portb28),
	.datac(gnd),
	.datad(\ShiftLeft0~68_combout ),
	.cin(gnd),
	.combout(\ShiftLeft0~69_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftLeft0~69 .lut_mask = 16'hBB88;
defparam \ShiftLeft0~69 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y42_N16
cycloneive_lcell_comb \Selector1~5 (
// Equation(s):
// \Selector1~5_combout  = (\portb~62_combout  & (\ShiftLeft0~58_combout )) # (!\portb~62_combout  & ((\ShiftLeft0~69_combout )))

	.dataa(gnd),
	.datab(portb29),
	.datac(\ShiftLeft0~58_combout ),
	.datad(\ShiftLeft0~69_combout ),
	.cin(gnd),
	.combout(\Selector1~5_combout ),
	.cout());
// synopsys translate_off
defparam \Selector1~5 .lut_mask = 16'hF3C0;
defparam \Selector1~5 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X52_Y42_N10
cycloneive_lcell_comb \Selector9~5 (
// Equation(s):
// \Selector9~5_combout  = (\Selector0~19_combout  & ((\Selector9~0_combout ) # ((\Selector0~21_combout  & \Selector1~5_combout )))) # (!\Selector0~19_combout  & (((\Selector0~21_combout  & \Selector1~5_combout ))))

	.dataa(\Selector0~19_combout ),
	.datab(\Selector9~0_combout ),
	.datac(\Selector0~21_combout ),
	.datad(\Selector1~5_combout ),
	.cin(gnd),
	.combout(\Selector9~5_combout ),
	.cout());
// synopsys translate_off
defparam \Selector9~5 .lut_mask = 16'hF888;
defparam \Selector9~5 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X52_Y39_N12
cycloneive_lcell_comb \Selector9~6 (
// Equation(s):
// \Selector9~6_combout  = (\Selector9~4_combout ) # ((\Selector9~5_combout ) # ((\ShiftLeft0~20_combout  & \Selector8~2_combout )))

	.dataa(\Selector9~4_combout ),
	.datab(\ShiftLeft0~20_combout ),
	.datac(\Selector8~2_combout ),
	.datad(\Selector9~5_combout ),
	.cin(gnd),
	.combout(\Selector9~6_combout ),
	.cout());
// synopsys translate_off
defparam \Selector9~6 .lut_mask = 16'hFFEA;
defparam \Selector9~6 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X52_Y39_N6
cycloneive_lcell_comb \Selector9~7 (
// Equation(s):
// \Selector9~7_combout  = (\Selector9~2_combout ) # ((\Selector9~6_combout ) # ((\Selector0~9_combout  & \Add0~44_combout )))

	.dataa(\Selector0~9_combout ),
	.datab(\Selector9~2_combout ),
	.datac(\Add0~44_combout ),
	.datad(\Selector9~6_combout ),
	.cin(gnd),
	.combout(\Selector9~7_combout ),
	.cout());
// synopsys translate_off
defparam \Selector9~7 .lut_mask = 16'hFFEC;
defparam \Selector9~7 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y39_N16
cycloneive_lcell_comb \Add1~48 (
// Equation(s):
// \Add1~48_combout  = ((\portb~18_combout  $ (\porta~111_combout  $ (\Add1~47 )))) # (GND)
// \Add1~49  = CARRY((\portb~18_combout  & (\porta~111_combout  & !\Add1~47 )) # (!\portb~18_combout  & ((\porta~111_combout ) # (!\Add1~47 ))))

	.dataa(portb7),
	.datab(porta27),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add1~47 ),
	.combout(\Add1~48_combout ),
	.cout(\Add1~49 ));
// synopsys translate_off
defparam \Add1~48 .lut_mask = 16'h964D;
defparam \Add1~48 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X57_Y39_N18
cycloneive_lcell_comb \Add1~50 (
// Equation(s):
// \Add1~50_combout  = (\porta~110_combout  & ((\portb~16_combout  & (!\Add1~49 )) # (!\portb~16_combout  & (\Add1~49  & VCC)))) # (!\porta~110_combout  & ((\portb~16_combout  & ((\Add1~49 ) # (GND))) # (!\portb~16_combout  & (!\Add1~49 ))))
// \Add1~51  = CARRY((\porta~110_combout  & (\portb~16_combout  & !\Add1~49 )) # (!\porta~110_combout  & ((\portb~16_combout ) # (!\Add1~49 ))))

	.dataa(porta26),
	.datab(portb6),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add1~49 ),
	.combout(\Add1~50_combout ),
	.cout(\Add1~51 ));
// synopsys translate_off
defparam \Add1~50 .lut_mask = 16'h694D;
defparam \Add1~50 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X52_Y37_N16
cycloneive_lcell_comb \Add0~48 (
// Equation(s):
// \Add0~48_combout  = ((\portb~18_combout  $ (\porta~111_combout  $ (!\Add0~47 )))) # (GND)
// \Add0~49  = CARRY((\portb~18_combout  & ((\porta~111_combout ) # (!\Add0~47 ))) # (!\portb~18_combout  & (\porta~111_combout  & !\Add0~47 )))

	.dataa(portb7),
	.datab(porta27),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add0~47 ),
	.combout(\Add0~48_combout ),
	.cout(\Add0~49 ));
// synopsys translate_off
defparam \Add0~48 .lut_mask = 16'h698E;
defparam \Add0~48 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X52_Y37_N18
cycloneive_lcell_comb \Add0~50 (
// Equation(s):
// \Add0~50_combout  = (\portb~16_combout  & ((\porta~110_combout  & (\Add0~49  & VCC)) # (!\porta~110_combout  & (!\Add0~49 )))) # (!\portb~16_combout  & ((\porta~110_combout  & (!\Add0~49 )) # (!\porta~110_combout  & ((\Add0~49 ) # (GND)))))
// \Add0~51  = CARRY((\portb~16_combout  & (!\porta~110_combout  & !\Add0~49 )) # (!\portb~16_combout  & ((!\Add0~49 ) # (!\porta~110_combout ))))

	.dataa(portb6),
	.datab(porta26),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add0~49 ),
	.combout(\Add0~50_combout ),
	.cout(\Add0~51 ));
// synopsys translate_off
defparam \Add0~50 .lut_mask = 16'h9617;
defparam \Add0~50 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X54_Y36_N14
cycloneive_lcell_comb \Selector6~7 (
// Equation(s):
// \Selector6~7_combout  = (\Add0~50_combout  & \Selector0~5_combout )

	.dataa(\Add0~50_combout ),
	.datab(gnd),
	.datac(gnd),
	.datad(\Selector0~5_combout ),
	.cin(gnd),
	.combout(\Selector6~7_combout ),
	.cout());
// synopsys translate_off
defparam \Selector6~7 .lut_mask = 16'hAA00;
defparam \Selector6~7 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y38_N16
cycloneive_lcell_comb \Selector4~0 (
// Equation(s):
// \Selector4~0_combout  = (!\ShiftRight0~72_combout  & (\Selector0~0_combout  & (!\portb~66_combout  & !\portb~64_combout )))

	.dataa(\ShiftRight0~72_combout ),
	.datab(\Selector0~0_combout ),
	.datac(portb31),
	.datad(portb30),
	.cin(gnd),
	.combout(\Selector4~0_combout ),
	.cout());
// synopsys translate_off
defparam \Selector4~0 .lut_mask = 16'h0004;
defparam \Selector4~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y36_N28
cycloneive_lcell_comb \Selector6~0 (
// Equation(s):
// \Selector6~0_combout  = (\portb~16_combout  & ((\Selector0~3_combout ) # ((\porta~110_combout  & \Selector0~4_combout ))))

	.dataa(porta26),
	.datab(\Selector0~3_combout ),
	.datac(portb6),
	.datad(\Selector0~4_combout ),
	.cin(gnd),
	.combout(\Selector6~0_combout ),
	.cout());
// synopsys translate_off
defparam \Selector6~0 .lut_mask = 16'hE0C0;
defparam \Selector6~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y36_N8
cycloneive_lcell_comb \porto~0 (
// Equation(s):
// \porto~0_combout  = \portb~16_combout  $ (((\porta~81_combout ) # ((plif_idexrdat1_l_25 & !\porta~63_combout ))))

	.dataa(portb6),
	.datab(porta6),
	.datac(plif_idexrdat1_l_25),
	.datad(porta4),
	.cin(gnd),
	.combout(\porto~0_combout ),
	.cout());
// synopsys translate_off
defparam \porto~0 .lut_mask = 16'h6656;
defparam \porto~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y36_N2
cycloneive_lcell_comb \Selector6~1 (
// Equation(s):
// \Selector6~1_combout  = (\porta~110_combout  & (((\Selector0~3_combout )))) # (!\porta~110_combout  & (!\portb~16_combout  & ((\Selector0~7_combout ))))

	.dataa(portb6),
	.datab(\Selector0~3_combout ),
	.datac(\Selector0~7_combout ),
	.datad(porta26),
	.cin(gnd),
	.combout(\Selector6~1_combout ),
	.cout());
// synopsys translate_off
defparam \Selector6~1 .lut_mask = 16'hCC50;
defparam \Selector6~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y36_N14
cycloneive_lcell_comb \Selector6~2 (
// Equation(s):
// \Selector6~2_combout  = (\Selector6~0_combout ) # ((\Selector6~1_combout ) # ((\Selector0~2_combout  & \porto~0_combout )))

	.dataa(\Selector0~2_combout ),
	.datab(\Selector6~0_combout ),
	.datac(\porto~0_combout ),
	.datad(\Selector6~1_combout ),
	.cin(gnd),
	.combout(\Selector6~2_combout ),
	.cout());
// synopsys translate_off
defparam \Selector6~2 .lut_mask = 16'hFFEC;
defparam \Selector6~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y36_N30
cycloneive_lcell_comb \ShiftLeft0~70 (
// Equation(s):
// \ShiftLeft0~70_combout  = (\portb~58_combout  & ((\porta~111_combout ))) # (!\portb~58_combout  & (\porta~110_combout ))

	.dataa(portb27),
	.datab(gnd),
	.datac(porta26),
	.datad(porta27),
	.cin(gnd),
	.combout(\ShiftLeft0~70_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftLeft0~70 .lut_mask = 16'hFA50;
defparam \ShiftLeft0~70 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y36_N8
cycloneive_lcell_comb \ShiftLeft0~71 (
// Equation(s):
// \ShiftLeft0~71_combout  = (\portb~60_combout  & ((\ShiftLeft0~66_combout ))) # (!\portb~60_combout  & (\ShiftLeft0~70_combout ))

	.dataa(portb28),
	.datab(gnd),
	.datac(\ShiftLeft0~70_combout ),
	.datad(\ShiftLeft0~66_combout ),
	.cin(gnd),
	.combout(\ShiftLeft0~71_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftLeft0~71 .lut_mask = 16'hFA50;
defparam \ShiftLeft0~71 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y36_N22
cycloneive_lcell_comb \ShiftLeft0~61 (
// Equation(s):
// \ShiftLeft0~61_combout  = (\portb~60_combout  & (\ShiftLeft0~54_combout )) # (!\portb~60_combout  & ((\ShiftLeft0~60_combout )))

	.dataa(portb28),
	.datab(gnd),
	.datac(\ShiftLeft0~54_combout ),
	.datad(\ShiftLeft0~60_combout ),
	.cin(gnd),
	.combout(\ShiftLeft0~61_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftLeft0~61 .lut_mask = 16'hF5A0;
defparam \ShiftLeft0~61 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X50_Y38_N22
cycloneive_lcell_comb \Selector6~3 (
// Equation(s):
// \Selector6~3_combout  = (\Selector7~0_combout  & (((!\Selector7~1_combout )))) # (!\Selector7~0_combout  & ((\Selector7~1_combout  & ((\ShiftLeft0~61_combout ))) # (!\Selector7~1_combout  & (\ShiftLeft0~71_combout ))))

	.dataa(\Selector7~0_combout ),
	.datab(\ShiftLeft0~71_combout ),
	.datac(\ShiftLeft0~61_combout ),
	.datad(\Selector7~1_combout ),
	.cin(gnd),
	.combout(\Selector6~3_combout ),
	.cout());
// synopsys translate_off
defparam \Selector6~3 .lut_mask = 16'h50EE;
defparam \Selector6~3 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X50_Y38_N16
cycloneive_lcell_comb \Selector6~4 (
// Equation(s):
// \Selector6~4_combout  = (!\ShiftRight0~72_combout  & ((\Selector7~0_combout  & ((\ShiftLeft0~50_combout ) # (!\Selector6~3_combout ))) # (!\Selector7~0_combout  & (\Selector6~3_combout ))))

	.dataa(\Selector7~0_combout ),
	.datab(\ShiftRight0~72_combout ),
	.datac(\Selector6~3_combout ),
	.datad(\ShiftLeft0~50_combout ),
	.cin(gnd),
	.combout(\Selector6~4_combout ),
	.cout());
// synopsys translate_off
defparam \Selector6~4 .lut_mask = 16'h3212;
defparam \Selector6~4 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X50_Y38_N6
cycloneive_lcell_comb \Selector6~5 (
// Equation(s):
// \Selector6~5_combout  = (\Selector0~1_combout  & (\Selector6~4_combout  & ((\ShiftLeft0~25_combout ) # (\Selector6~3_combout ))))

	.dataa(\ShiftLeft0~25_combout ),
	.datab(\Selector0~1_combout ),
	.datac(\Selector6~3_combout ),
	.datad(\Selector6~4_combout ),
	.cin(gnd),
	.combout(\Selector6~5_combout ),
	.cout());
// synopsys translate_off
defparam \Selector6~5 .lut_mask = 16'hC800;
defparam \Selector6~5 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y36_N16
cycloneive_lcell_comb \Selector6~6 (
// Equation(s):
// \Selector6~6_combout  = (\Selector6~2_combout ) # ((\Selector6~5_combout ) # ((\Selector4~0_combout  & \ShiftRight0~32_combout )))

	.dataa(\Selector4~0_combout ),
	.datab(\Selector6~2_combout ),
	.datac(\ShiftRight0~32_combout ),
	.datad(\Selector6~5_combout ),
	.cin(gnd),
	.combout(\Selector6~6_combout ),
	.cout());
// synopsys translate_off
defparam \Selector6~6 .lut_mask = 16'hFFEC;
defparam \Selector6~6 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y38_N4
cycloneive_lcell_comb \Selector7~9 (
// Equation(s):
// \Selector7~9_combout  = (\portb~18_combout  & ((\Selector0~3_combout ) # ((\Selector0~4_combout  & \porta~111_combout ))))

	.dataa(\Selector0~3_combout ),
	.datab(\Selector0~4_combout ),
	.datac(portb7),
	.datad(porta27),
	.cin(gnd),
	.combout(\Selector7~9_combout ),
	.cout());
// synopsys translate_off
defparam \Selector7~9 .lut_mask = 16'hE0A0;
defparam \Selector7~9 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y38_N18
cycloneive_lcell_comb \Selector7~8 (
// Equation(s):
// \Selector7~8_combout  = (!\portb~64_combout  & (\Selector0~0_combout  & (\ShiftRight0~63_combout  & !\Selector1~1_combout )))

	.dataa(portb30),
	.datab(\Selector0~0_combout ),
	.datac(\ShiftRight0~63_combout ),
	.datad(\Selector1~1_combout ),
	.cin(gnd),
	.combout(\Selector7~8_combout ),
	.cout());
// synopsys translate_off
defparam \Selector7~8 .lut_mask = 16'h0040;
defparam \Selector7~8 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y38_N30
cycloneive_lcell_comb \Selector7~10 (
// Equation(s):
// \Selector7~10_combout  = (\Selector7~9_combout ) # (\Selector7~8_combout )

	.dataa(gnd),
	.datab(gnd),
	.datac(\Selector7~9_combout ),
	.datad(\Selector7~8_combout ),
	.cin(gnd),
	.combout(\Selector7~10_combout ),
	.cout());
// synopsys translate_off
defparam \Selector7~10 .lut_mask = 16'hFFF0;
defparam \Selector7~10 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y35_N0
cycloneive_lcell_comb \Selector7~2 (
// Equation(s):
// \Selector7~2_combout  = (\porta~111_combout  & (\Selector0~3_combout )) # (!\porta~111_combout  & (((\Selector0~7_combout  & !\portb~18_combout ))))

	.dataa(\Selector0~3_combout ),
	.datab(\Selector0~7_combout ),
	.datac(portb7),
	.datad(porta27),
	.cin(gnd),
	.combout(\Selector7~2_combout ),
	.cout());
// synopsys translate_off
defparam \Selector7~2 .lut_mask = 16'hAA0C;
defparam \Selector7~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y35_N30
cycloneive_lcell_comb \Selector7~3 (
// Equation(s):
// \Selector7~3_combout  = (\Selector7~2_combout ) # ((\Selector0~2_combout  & (\portb~18_combout  $ (\porta~111_combout ))))

	.dataa(portb7),
	.datab(\Selector7~2_combout ),
	.datac(\Selector0~2_combout ),
	.datad(porta27),
	.cin(gnd),
	.combout(\Selector7~3_combout ),
	.cout());
// synopsys translate_off
defparam \Selector7~3 .lut_mask = 16'hDCEC;
defparam \Selector7~3 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X52_Y36_N8
cycloneive_lcell_comb \ShiftLeft0~73 (
// Equation(s):
// \ShiftLeft0~73_combout  = (\portb~60_combout  & ((\ShiftLeft0~68_combout ))) # (!\portb~60_combout  & (\ShiftLeft0~72_combout ))

	.dataa(\ShiftLeft0~72_combout ),
	.datab(gnd),
	.datac(portb28),
	.datad(\ShiftLeft0~68_combout ),
	.cin(gnd),
	.combout(\ShiftLeft0~73_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftLeft0~73 .lut_mask = 16'hFA0A;
defparam \ShiftLeft0~73 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y40_N24
cycloneive_lcell_comb \Selector7~4 (
// Equation(s):
// \Selector7~4_combout  = (\Selector7~1_combout  & (\Selector7~0_combout )) # (!\Selector7~1_combout  & ((\Selector7~0_combout  & ((\ShiftLeft0~53_combout ))) # (!\Selector7~0_combout  & (\ShiftLeft0~73_combout ))))

	.dataa(\Selector7~1_combout ),
	.datab(\Selector7~0_combout ),
	.datac(\ShiftLeft0~73_combout ),
	.datad(\ShiftLeft0~53_combout ),
	.cin(gnd),
	.combout(\Selector7~4_combout ),
	.cout());
// synopsys translate_off
defparam \Selector7~4 .lut_mask = 16'hDC98;
defparam \Selector7~4 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y40_N10
cycloneive_lcell_comb \ShiftLeft0~63 (
// Equation(s):
// \ShiftLeft0~63_combout  = (\portb~58_combout  & ((\porta~116_combout ))) # (!\portb~58_combout  & (\porta~115_combout ))

	.dataa(gnd),
	.datab(portb27),
	.datac(porta31),
	.datad(porta32),
	.cin(gnd),
	.combout(\ShiftLeft0~63_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftLeft0~63 .lut_mask = 16'hFC30;
defparam \ShiftLeft0~63 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y40_N4
cycloneive_lcell_comb \ShiftLeft0~64 (
// Equation(s):
// \ShiftLeft0~64_combout  = (\portb~60_combout  & (\ShiftLeft0~57_combout )) # (!\portb~60_combout  & ((\ShiftLeft0~63_combout )))

	.dataa(portb28),
	.datab(gnd),
	.datac(\ShiftLeft0~57_combout ),
	.datad(\ShiftLeft0~63_combout ),
	.cin(gnd),
	.combout(\ShiftLeft0~64_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftLeft0~64 .lut_mask = 16'hF5A0;
defparam \ShiftLeft0~64 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y35_N16
cycloneive_lcell_comb \Selector7~5 (
// Equation(s):
// \Selector7~5_combout  = (!\ShiftRight0~72_combout  & ((\Selector7~1_combout  & ((\ShiftLeft0~80_combout ) # (!\Selector7~4_combout ))) # (!\Selector7~1_combout  & ((\Selector7~4_combout )))))

	.dataa(\Selector7~1_combout ),
	.datab(\ShiftRight0~72_combout ),
	.datac(\ShiftLeft0~80_combout ),
	.datad(\Selector7~4_combout ),
	.cin(gnd),
	.combout(\Selector7~5_combout ),
	.cout());
// synopsys translate_off
defparam \Selector7~5 .lut_mask = 16'h3122;
defparam \Selector7~5 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y35_N10
cycloneive_lcell_comb \Selector7~6 (
// Equation(s):
// \Selector7~6_combout  = (\Selector0~1_combout  & (\Selector7~5_combout  & ((\Selector7~4_combout ) # (\ShiftLeft0~64_combout ))))

	.dataa(\Selector0~1_combout ),
	.datab(\Selector7~4_combout ),
	.datac(\ShiftLeft0~64_combout ),
	.datad(\Selector7~5_combout ),
	.cin(gnd),
	.combout(\Selector7~6_combout ),
	.cout());
// synopsys translate_off
defparam \Selector7~6 .lut_mask = 16'hA800;
defparam \Selector7~6 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y35_N24
cycloneive_lcell_comb \Selector7~7 (
// Equation(s):
// \Selector7~7_combout  = (\Selector7~3_combout ) # ((\Selector7~6_combout ) # ((\Add1~48_combout  & \Selector0~6_combout )))

	.dataa(\Add1~48_combout ),
	.datab(\Selector0~6_combout ),
	.datac(\Selector7~3_combout ),
	.datad(\Selector7~6_combout ),
	.cin(gnd),
	.combout(\Selector7~7_combout ),
	.cout());
// synopsys translate_off
defparam \Selector7~7 .lut_mask = 16'hFFF8;
defparam \Selector7~7 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y42_N22
cycloneive_lcell_comb \Selector4~8 (
// Equation(s):
// \Selector4~8_combout  = (\portb~12_combout  & ((\Selector0~3_combout ) # ((\porta~108_combout  & \Selector0~4_combout ))))

	.dataa(\Selector0~3_combout ),
	.datab(portb4),
	.datac(porta24),
	.datad(\Selector0~4_combout ),
	.cin(gnd),
	.combout(\Selector4~8_combout ),
	.cout());
// synopsys translate_off
defparam \Selector4~8 .lut_mask = 16'hC888;
defparam \Selector4~8 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y38_N12
cycloneive_lcell_comb \Selector4~7 (
// Equation(s):
// \Selector4~7_combout  = (!\portb~64_combout  & (\Selector0~0_combout  & (\ShiftRight0~81_combout  & !\Selector1~1_combout )))

	.dataa(portb30),
	.datab(\Selector0~0_combout ),
	.datac(\ShiftRight0~81_combout ),
	.datad(\Selector1~1_combout ),
	.cin(gnd),
	.combout(\Selector4~7_combout ),
	.cout());
// synopsys translate_off
defparam \Selector4~7 .lut_mask = 16'h0040;
defparam \Selector4~7 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y38_N2
cycloneive_lcell_comb \Selector4~9 (
// Equation(s):
// \Selector4~9_combout  = (\Selector4~8_combout ) # (\Selector4~7_combout )

	.dataa(gnd),
	.datab(gnd),
	.datac(\Selector4~8_combout ),
	.datad(\Selector4~7_combout ),
	.cin(gnd),
	.combout(\Selector4~9_combout ),
	.cout());
// synopsys translate_off
defparam \Selector4~9 .lut_mask = 16'hFFF0;
defparam \Selector4~9 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y39_N20
cycloneive_lcell_comb \Add1~52 (
// Equation(s):
// \Add1~52_combout  = ((\porta~109_combout  $ (\portb~14_combout  $ (\Add1~51 )))) # (GND)
// \Add1~53  = CARRY((\porta~109_combout  & ((!\Add1~51 ) # (!\portb~14_combout ))) # (!\porta~109_combout  & (!\portb~14_combout  & !\Add1~51 )))

	.dataa(porta25),
	.datab(portb5),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add1~51 ),
	.combout(\Add1~52_combout ),
	.cout(\Add1~53 ));
// synopsys translate_off
defparam \Add1~52 .lut_mask = 16'h962B;
defparam \Add1~52 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X57_Y39_N22
cycloneive_lcell_comb \Add1~54 (
// Equation(s):
// \Add1~54_combout  = (\porta~108_combout  & ((\portb~12_combout  & (!\Add1~53 )) # (!\portb~12_combout  & (\Add1~53  & VCC)))) # (!\porta~108_combout  & ((\portb~12_combout  & ((\Add1~53 ) # (GND))) # (!\portb~12_combout  & (!\Add1~53 ))))
// \Add1~55  = CARRY((\porta~108_combout  & (\portb~12_combout  & !\Add1~53 )) # (!\porta~108_combout  & ((\portb~12_combout ) # (!\Add1~53 ))))

	.dataa(porta24),
	.datab(portb4),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add1~53 ),
	.combout(\Add1~54_combout ),
	.cout(\Add1~55 ));
// synopsys translate_off
defparam \Add1~54 .lut_mask = 16'h694D;
defparam \Add1~54 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X57_Y36_N20
cycloneive_lcell_comb \Selector4~4 (
// Equation(s):
// \Selector4~4_combout  = (\porta~108_combout  & (((\Selector0~3_combout )))) # (!\porta~108_combout  & (\Selector0~7_combout  & (!\portb~12_combout )))

	.dataa(\Selector0~7_combout ),
	.datab(portb4),
	.datac(porta24),
	.datad(\Selector0~3_combout ),
	.cin(gnd),
	.combout(\Selector4~4_combout ),
	.cout());
// synopsys translate_off
defparam \Selector4~4 .lut_mask = 16'hF202;
defparam \Selector4~4 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y36_N26
cycloneive_lcell_comb \Selector4~5 (
// Equation(s):
// \Selector4~5_combout  = (\Selector4~4_combout ) # ((\Selector0~2_combout  & (\portb~12_combout  $ (\porta~108_combout ))))

	.dataa(\Selector0~2_combout ),
	.datab(portb4),
	.datac(porta24),
	.datad(\Selector4~4_combout ),
	.cin(gnd),
	.combout(\Selector4~5_combout ),
	.cout());
// synopsys translate_off
defparam \Selector4~5 .lut_mask = 16'hFF28;
defparam \Selector4~5 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X52_Y37_N20
cycloneive_lcell_comb \Add0~52 (
// Equation(s):
// \Add0~52_combout  = ((\portb~14_combout  $ (\porta~109_combout  $ (!\Add0~51 )))) # (GND)
// \Add0~53  = CARRY((\portb~14_combout  & ((\porta~109_combout ) # (!\Add0~51 ))) # (!\portb~14_combout  & (\porta~109_combout  & !\Add0~51 )))

	.dataa(portb5),
	.datab(porta25),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add0~51 ),
	.combout(\Add0~52_combout ),
	.cout(\Add0~53 ));
// synopsys translate_off
defparam \Add0~52 .lut_mask = 16'h698E;
defparam \Add0~52 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X52_Y37_N22
cycloneive_lcell_comb \Add0~54 (
// Equation(s):
// \Add0~54_combout  = (\porta~108_combout  & ((\portb~12_combout  & (\Add0~53  & VCC)) # (!\portb~12_combout  & (!\Add0~53 )))) # (!\porta~108_combout  & ((\portb~12_combout  & (!\Add0~53 )) # (!\portb~12_combout  & ((\Add0~53 ) # (GND)))))
// \Add0~55  = CARRY((\porta~108_combout  & (!\portb~12_combout  & !\Add0~53 )) # (!\porta~108_combout  & ((!\Add0~53 ) # (!\portb~12_combout ))))

	.dataa(porta24),
	.datab(portb4),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add0~53 ),
	.combout(\Add0~54_combout ),
	.cout(\Add0~55 ));
// synopsys translate_off
defparam \Add0~54 .lut_mask = 16'h9617;
defparam \Add0~54 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X50_Y37_N20
cycloneive_lcell_comb \ShiftLeft0~74 (
// Equation(s):
// \ShiftLeft0~74_combout  = (\portb~58_combout  & (\porta~109_combout )) # (!\portb~58_combout  & ((\porta~108_combout )))

	.dataa(gnd),
	.datab(porta25),
	.datac(portb27),
	.datad(porta24),
	.cin(gnd),
	.combout(\ShiftLeft0~74_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftLeft0~74 .lut_mask = 16'hCFC0;
defparam \ShiftLeft0~74 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y36_N2
cycloneive_lcell_comb \ShiftLeft0~75 (
// Equation(s):
// \ShiftLeft0~75_combout  = (\portb~60_combout  & (\ShiftLeft0~70_combout )) # (!\portb~60_combout  & ((\ShiftLeft0~74_combout )))

	.dataa(\ShiftLeft0~70_combout ),
	.datab(gnd),
	.datac(portb28),
	.datad(\ShiftLeft0~74_combout ),
	.cin(gnd),
	.combout(\ShiftLeft0~75_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftLeft0~75 .lut_mask = 16'hAFA0;
defparam \ShiftLeft0~75 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y36_N4
cycloneive_lcell_comb \Selector4~1 (
// Equation(s):
// \Selector4~1_combout  = (\Selector7~0_combout  & (((\Selector7~1_combout )))) # (!\Selector7~0_combout  & ((\Selector7~1_combout  & (\ShiftLeft0~67_combout )) # (!\Selector7~1_combout  & ((\ShiftLeft0~75_combout )))))

	.dataa(\Selector7~0_combout ),
	.datab(\ShiftLeft0~67_combout ),
	.datac(\Selector7~1_combout ),
	.datad(\ShiftLeft0~75_combout ),
	.cin(gnd),
	.combout(\Selector4~1_combout ),
	.cout());
// synopsys translate_off
defparam \Selector4~1 .lut_mask = 16'hE5E0;
defparam \Selector4~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y36_N6
cycloneive_lcell_comb \Selector4~2 (
// Equation(s):
// \Selector4~2_combout  = (!\ShiftRight0~72_combout  & ((\Selector7~0_combout  & ((\ShiftLeft0~32_combout ) # (!\Selector4~1_combout ))) # (!\Selector7~0_combout  & (\Selector4~1_combout ))))

	.dataa(\Selector7~0_combout ),
	.datab(\Selector4~1_combout ),
	.datac(\ShiftRight0~72_combout ),
	.datad(\ShiftLeft0~32_combout ),
	.cin(gnd),
	.combout(\Selector4~2_combout ),
	.cout());
// synopsys translate_off
defparam \Selector4~2 .lut_mask = 16'h0E06;
defparam \Selector4~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y36_N12
cycloneive_lcell_comb \Selector4~3 (
// Equation(s):
// \Selector4~3_combout  = (\Selector0~1_combout  & (\Selector4~2_combout  & ((\ShiftLeft0~56_combout ) # (\Selector4~1_combout ))))

	.dataa(\ShiftLeft0~56_combout ),
	.datab(\Selector0~1_combout ),
	.datac(\Selector4~1_combout ),
	.datad(\Selector4~2_combout ),
	.cin(gnd),
	.combout(\Selector4~3_combout ),
	.cout());
// synopsys translate_off
defparam \Selector4~3 .lut_mask = 16'hC800;
defparam \Selector4~3 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y36_N14
cycloneive_lcell_comb \Selector4~6 (
// Equation(s):
// \Selector4~6_combout  = (\Selector4~5_combout ) # ((\Selector4~3_combout ) # ((\Selector0~5_combout  & \Add0~54_combout )))

	.dataa(\Selector0~5_combout ),
	.datab(\Selector4~5_combout ),
	.datac(\Add0~54_combout ),
	.datad(\Selector4~3_combout ),
	.cin(gnd),
	.combout(\Selector4~6_combout ),
	.cout());
// synopsys translate_off
defparam \Selector4~6 .lut_mask = 16'hFFEC;
defparam \Selector4~6 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y42_N4
cycloneive_lcell_comb \Selector5~0 (
// Equation(s):
// \Selector5~0_combout  = (\porta~109_combout  & ((\Selector0~4_combout ))) # (!\porta~109_combout  & (\Selector0~7_combout ))

	.dataa(\Selector0~7_combout ),
	.datab(gnd),
	.datac(\Selector0~4_combout ),
	.datad(porta25),
	.cin(gnd),
	.combout(\Selector5~0_combout ),
	.cout());
// synopsys translate_off
defparam \Selector5~0 .lut_mask = 16'hF0AA;
defparam \Selector5~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y42_N10
cycloneive_lcell_comb \Selector5~1 (
// Equation(s):
// \Selector5~1_combout  = (\portb~14_combout  & ((\Selector0~3_combout ) # (!\porta~109_combout ))) # (!\portb~14_combout  & ((\porta~109_combout )))

	.dataa(\Selector0~3_combout ),
	.datab(gnd),
	.datac(portb5),
	.datad(porta25),
	.cin(gnd),
	.combout(\Selector5~1_combout ),
	.cout());
// synopsys translate_off
defparam \Selector5~1 .lut_mask = 16'hAFF0;
defparam \Selector5~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y42_N0
cycloneive_lcell_comb \Selector5~2 (
// Equation(s):
// \Selector5~2_combout  = (\Selector5~1_combout  & ((\Selector0~3_combout ) # ((\Selector0~2_combout )))) # (!\Selector5~1_combout  & (((\Selector5~0_combout ))))

	.dataa(\Selector0~3_combout ),
	.datab(\Selector0~2_combout ),
	.datac(\Selector5~0_combout ),
	.datad(\Selector5~1_combout ),
	.cin(gnd),
	.combout(\Selector5~2_combout ),
	.cout());
// synopsys translate_off
defparam \Selector5~2 .lut_mask = 16'hEEF0;
defparam \Selector5~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X52_Y36_N0
cycloneive_lcell_comb \ShiftLeft0~76 (
// Equation(s):
// \ShiftLeft0~76_combout  = (\portb~58_combout  & (\porta~110_combout )) # (!\portb~58_combout  & ((\porta~109_combout )))

	.dataa(porta26),
	.datab(porta25),
	.datac(gnd),
	.datad(portb27),
	.cin(gnd),
	.combout(\ShiftLeft0~76_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftLeft0~76 .lut_mask = 16'hAACC;
defparam \ShiftLeft0~76 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X52_Y36_N2
cycloneive_lcell_comb \ShiftLeft0~77 (
// Equation(s):
// \ShiftLeft0~77_combout  = (\portb~60_combout  & (\ShiftLeft0~72_combout )) # (!\portb~60_combout  & ((\ShiftLeft0~76_combout )))

	.dataa(\ShiftLeft0~72_combout ),
	.datab(gnd),
	.datac(portb28),
	.datad(\ShiftLeft0~76_combout ),
	.cin(gnd),
	.combout(\ShiftLeft0~77_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftLeft0~77 .lut_mask = 16'hAFA0;
defparam \ShiftLeft0~77 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y40_N0
cycloneive_lcell_comb \ShiftLeft0~59 (
// Equation(s):
// \ShiftLeft0~59_combout  = (\portb~62_combout  & ((\ShiftLeft0~46_combout ))) # (!\portb~62_combout  & (\ShiftLeft0~58_combout ))

	.dataa(gnd),
	.datab(\ShiftLeft0~58_combout ),
	.datac(portb29),
	.datad(\ShiftLeft0~46_combout ),
	.cin(gnd),
	.combout(\ShiftLeft0~59_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftLeft0~59 .lut_mask = 16'hFC0C;
defparam \ShiftLeft0~59 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y40_N24
cycloneive_lcell_comb \Selector5~3 (
// Equation(s):
// \Selector5~3_combout  = (\Selector7~1_combout  & (!\Selector7~0_combout )) # (!\Selector7~1_combout  & ((\Selector7~0_combout  & ((\ShiftLeft0~59_combout ))) # (!\Selector7~0_combout  & (\ShiftLeft0~77_combout ))))

	.dataa(\Selector7~1_combout ),
	.datab(\Selector7~0_combout ),
	.datac(\ShiftLeft0~77_combout ),
	.datad(\ShiftLeft0~59_combout ),
	.cin(gnd),
	.combout(\Selector5~3_combout ),
	.cout());
// synopsys translate_off
defparam \Selector5~3 .lut_mask = 16'h7632;
defparam \Selector5~3 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y40_N6
cycloneive_lcell_comb \Selector5~4 (
// Equation(s):
// \Selector5~4_combout  = (!\ShiftRight0~72_combout  & ((\Selector7~1_combout  & ((\ShiftLeft0~69_combout ) # (!\Selector5~3_combout ))) # (!\Selector7~1_combout  & ((\Selector5~3_combout )))))

	.dataa(\ShiftLeft0~69_combout ),
	.datab(\ShiftRight0~72_combout ),
	.datac(\Selector7~1_combout ),
	.datad(\Selector5~3_combout ),
	.cin(gnd),
	.combout(\Selector5~4_combout ),
	.cout());
// synopsys translate_off
defparam \Selector5~4 .lut_mask = 16'h2330;
defparam \Selector5~4 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y40_N12
cycloneive_lcell_comb \Selector5~5 (
// Equation(s):
// \Selector5~5_combout  = (\Selector0~1_combout  & (\Selector5~4_combout  & ((\Selector5~3_combout ) # (\ShiftLeft0~36_combout ))))

	.dataa(\Selector0~1_combout ),
	.datab(\Selector5~3_combout ),
	.datac(\ShiftLeft0~36_combout ),
	.datad(\Selector5~4_combout ),
	.cin(gnd),
	.combout(\Selector5~5_combout ),
	.cout());
// synopsys translate_off
defparam \Selector5~5 .lut_mask = 16'hA800;
defparam \Selector5~5 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y40_N14
cycloneive_lcell_comb \Selector5~6 (
// Equation(s):
// \Selector5~6_combout  = (\Selector5~2_combout ) # ((\Selector5~5_combout ) # ((\Selector4~0_combout  & \ShiftRight0~90_combout )))

	.dataa(\Selector4~0_combout ),
	.datab(\ShiftRight0~90_combout ),
	.datac(\Selector5~2_combout ),
	.datad(\Selector5~5_combout ),
	.cin(gnd),
	.combout(\Selector5~6_combout ),
	.cout());
// synopsys translate_off
defparam \Selector5~6 .lut_mask = 16'hFFF8;
defparam \Selector5~6 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y36_N24
cycloneive_lcell_comb \Selector5~7 (
// Equation(s):
// \Selector5~7_combout  = (\Selector0~6_combout  & \Add1~52_combout )

	.dataa(\Selector0~6_combout ),
	.datab(gnd),
	.datac(gnd),
	.datad(\Add1~52_combout ),
	.cin(gnd),
	.combout(\Selector5~7_combout ),
	.cout());
// synopsys translate_off
defparam \Selector5~7 .lut_mask = 16'hAA00;
defparam \Selector5~7 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y39_N24
cycloneive_lcell_comb \Add1~56 (
// Equation(s):
// \Add1~56_combout  = ((\portb~10_combout  $ (\porta~107_combout  $ (\Add1~55 )))) # (GND)
// \Add1~57  = CARRY((\portb~10_combout  & (\porta~107_combout  & !\Add1~55 )) # (!\portb~10_combout  & ((\porta~107_combout ) # (!\Add1~55 ))))

	.dataa(portb3),
	.datab(porta23),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add1~55 ),
	.combout(\Add1~56_combout ),
	.cout(\Add1~57 ));
// synopsys translate_off
defparam \Add1~56 .lut_mask = 16'h964D;
defparam \Add1~56 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X57_Y39_N26
cycloneive_lcell_comb \Add1~58 (
// Equation(s):
// \Add1~58_combout  = (\portb~8_combout  & ((\porta~105_combout  & (!\Add1~57 )) # (!\porta~105_combout  & ((\Add1~57 ) # (GND))))) # (!\portb~8_combout  & ((\porta~105_combout  & (\Add1~57  & VCC)) # (!\porta~105_combout  & (!\Add1~57 ))))
// \Add1~59  = CARRY((\portb~8_combout  & ((!\Add1~57 ) # (!\porta~105_combout ))) # (!\portb~8_combout  & (!\porta~105_combout  & !\Add1~57 )))

	.dataa(portb2),
	.datab(porta21),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add1~57 ),
	.combout(\Add1~58_combout ),
	.cout(\Add1~59 ));
// synopsys translate_off
defparam \Add1~58 .lut_mask = 16'h692B;
defparam \Add1~58 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X52_Y37_N24
cycloneive_lcell_comb \Add0~56 (
// Equation(s):
// \Add0~56_combout  = ((\portb~10_combout  $ (\porta~107_combout  $ (!\Add0~55 )))) # (GND)
// \Add0~57  = CARRY((\portb~10_combout  & ((\porta~107_combout ) # (!\Add0~55 ))) # (!\portb~10_combout  & (\porta~107_combout  & !\Add0~55 )))

	.dataa(portb3),
	.datab(porta23),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add0~55 ),
	.combout(\Add0~56_combout ),
	.cout(\Add0~57 ));
// synopsys translate_off
defparam \Add0~56 .lut_mask = 16'h698E;
defparam \Add0~56 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X52_Y37_N26
cycloneive_lcell_comb \Add0~58 (
// Equation(s):
// \Add0~58_combout  = (\portb~8_combout  & ((\porta~105_combout  & (\Add0~57  & VCC)) # (!\porta~105_combout  & (!\Add0~57 )))) # (!\portb~8_combout  & ((\porta~105_combout  & (!\Add0~57 )) # (!\porta~105_combout  & ((\Add0~57 ) # (GND)))))
// \Add0~59  = CARRY((\portb~8_combout  & (!\porta~105_combout  & !\Add0~57 )) # (!\portb~8_combout  & ((!\Add0~57 ) # (!\porta~105_combout ))))

	.dataa(portb2),
	.datab(porta21),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add0~57 ),
	.combout(\Add0~58_combout ),
	.cout(\Add0~59 ));
// synopsys translate_off
defparam \Add0~58 .lut_mask = 16'h9617;
defparam \Add0~58 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X50_Y39_N22
cycloneive_lcell_comb \Selector2~10 (
// Equation(s):
// \Selector2~10_combout  = (\Selector0~9_combout  & \Add0~58_combout )

	.dataa(gnd),
	.datab(\Selector0~9_combout ),
	.datac(gnd),
	.datad(\Add0~58_combout ),
	.cin(gnd),
	.combout(\Selector2~10_combout ),
	.cout());
// synopsys translate_off
defparam \Selector2~10 .lut_mask = 16'hCC00;
defparam \Selector2~10 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y33_N28
cycloneive_lcell_comb \Selector2~0 (
// Equation(s):
// \Selector2~0_combout  = (\portb~8_combout  & ((\Selector0~10_combout ) # ((\Selector0~11_combout  & \porta~105_combout ))))

	.dataa(\Selector0~10_combout ),
	.datab(portb2),
	.datac(\Selector0~11_combout ),
	.datad(porta21),
	.cin(gnd),
	.combout(\Selector2~0_combout ),
	.cout());
// synopsys translate_off
defparam \Selector2~0 .lut_mask = 16'hC888;
defparam \Selector2~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y33_N26
cycloneive_lcell_comb \Selector2~1 (
// Equation(s):
// \Selector2~1_combout  = (\porta~105_combout  & (\Selector0~10_combout )) # (!\porta~105_combout  & (((!\portb~8_combout  & \Selector0~12_combout ))))

	.dataa(\Selector0~10_combout ),
	.datab(portb2),
	.datac(\Selector0~12_combout ),
	.datad(porta21),
	.cin(gnd),
	.combout(\Selector2~1_combout ),
	.cout());
// synopsys translate_off
defparam \Selector2~1 .lut_mask = 16'hAA30;
defparam \Selector2~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y33_N0
cycloneive_lcell_comb \porto~1 (
// Equation(s):
// \porto~1_combout  = \portb~8_combout  $ (((\porta~76_combout ) # ((!\porta~63_combout  & plif_idexrdat1_l_29))))

	.dataa(porta4),
	.datab(porta5),
	.datac(plif_idexrdat1_l_29),
	.datad(portb2),
	.cin(gnd),
	.combout(\porto~1_combout ),
	.cout());
// synopsys translate_off
defparam \porto~1 .lut_mask = 16'h23DC;
defparam \porto~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y33_N30
cycloneive_lcell_comb \Selector2~2 (
// Equation(s):
// \Selector2~2_combout  = (\Selector2~0_combout ) # ((\Selector2~1_combout ) # ((\Selector0~13_combout  & \porto~1_combout )))

	.dataa(\Selector0~13_combout ),
	.datab(\Selector2~0_combout ),
	.datac(\Selector2~1_combout ),
	.datad(\porto~1_combout ),
	.cin(gnd),
	.combout(\Selector2~2_combout ),
	.cout());
// synopsys translate_off
defparam \Selector2~2 .lut_mask = 16'hFEFC;
defparam \Selector2~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X50_Y37_N30
cycloneive_lcell_comb \Selector2~3 (
// Equation(s):
// \Selector2~3_combout  = (\portb~66_combout  & (!plif_idexaluop_l_0 & (\Selector1~3_combout  & \ShiftLeft0~39_combout )))

	.dataa(portb31),
	.datab(plif_idexaluop_l_0),
	.datac(\Selector1~3_combout ),
	.datad(\ShiftLeft0~39_combout ),
	.cin(gnd),
	.combout(\Selector2~3_combout ),
	.cout());
// synopsys translate_off
defparam \Selector2~3 .lut_mask = 16'h2000;
defparam \Selector2~3 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X50_Y37_N0
cycloneive_lcell_comb \Selector2~4 (
// Equation(s):
// \Selector2~4_combout  = (!\portb~66_combout  & (\Selector0~20_combout  & (\ShiftRight0~74_combout  & !\ShiftRight0~72_combout )))

	.dataa(portb31),
	.datab(\Selector0~20_combout ),
	.datac(\ShiftRight0~74_combout ),
	.datad(\ShiftRight0~72_combout ),
	.cin(gnd),
	.combout(\Selector2~4_combout ),
	.cout());
// synopsys translate_off
defparam \Selector2~4 .lut_mask = 16'h0040;
defparam \Selector2~4 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X50_Y37_N24
cycloneive_lcell_comb \ShiftLeft0~78 (
// Equation(s):
// \ShiftLeft0~78_combout  = (\portb~58_combout  & (\porta~107_combout )) # (!\portb~58_combout  & ((\porta~105_combout )))

	.dataa(portb27),
	.datab(gnd),
	.datac(porta23),
	.datad(porta21),
	.cin(gnd),
	.combout(\ShiftLeft0~78_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftLeft0~78 .lut_mask = 16'hF5A0;
defparam \ShiftLeft0~78 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X50_Y37_N18
cycloneive_lcell_comb \Selector2~6 (
// Equation(s):
// \Selector2~6_combout  = (\ShiftRight0~74_combout  & (\ShiftLeft0~78_combout  & ((!\Selector3~1_combout )))) # (!\ShiftRight0~74_combout  & (((\ShiftLeft0~71_combout ) # (\Selector3~1_combout ))))

	.dataa(\ShiftRight0~74_combout ),
	.datab(\ShiftLeft0~78_combout ),
	.datac(\ShiftLeft0~71_combout ),
	.datad(\Selector3~1_combout ),
	.cin(gnd),
	.combout(\Selector2~6_combout ),
	.cout());
// synopsys translate_off
defparam \Selector2~6 .lut_mask = 16'h55D8;
defparam \Selector2~6 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X50_Y37_N4
cycloneive_lcell_comb \Selector2~7 (
// Equation(s):
// \Selector2~7_combout  = (\Selector3~1_combout  & ((\Selector2~6_combout  & ((\ShiftLeft0~62_combout ))) # (!\Selector2~6_combout  & (\ShiftLeft0~74_combout )))) # (!\Selector3~1_combout  & (((\Selector2~6_combout ))))

	.dataa(\ShiftLeft0~74_combout ),
	.datab(\Selector3~1_combout ),
	.datac(\Selector2~6_combout ),
	.datad(\ShiftLeft0~62_combout ),
	.cin(gnd),
	.combout(\Selector2~7_combout ),
	.cout());
// synopsys translate_off
defparam \Selector2~7 .lut_mask = 16'hF838;
defparam \Selector2~7 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X50_Y37_N6
cycloneive_lcell_comb \Selector2~5 (
// Equation(s):
// \Selector2~5_combout  = (!plif_idexaluop_l_0 & (!plif_idexaluop_l_1 & (!\Selector3~0_combout  & !\ShiftRight0~72_combout )))

	.dataa(plif_idexaluop_l_0),
	.datab(plif_idexaluop_l_1),
	.datac(\Selector3~0_combout ),
	.datad(\ShiftRight0~72_combout ),
	.cin(gnd),
	.combout(\Selector2~5_combout ),
	.cout());
// synopsys translate_off
defparam \Selector2~5 .lut_mask = 16'h0001;
defparam \Selector2~5 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X50_Y37_N10
cycloneive_lcell_comb \Selector2~8 (
// Equation(s):
// \Selector2~8_combout  = (\ShiftRight0~28_combout  & ((\Selector2~4_combout ) # ((\Selector2~7_combout  & \Selector2~5_combout )))) # (!\ShiftRight0~28_combout  & (((\Selector2~7_combout  & \Selector2~5_combout ))))

	.dataa(\ShiftRight0~28_combout ),
	.datab(\Selector2~4_combout ),
	.datac(\Selector2~7_combout ),
	.datad(\Selector2~5_combout ),
	.cin(gnd),
	.combout(\Selector2~8_combout ),
	.cout());
// synopsys translate_off
defparam \Selector2~8 .lut_mask = 16'hF888;
defparam \Selector2~8 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X50_Y37_N16
cycloneive_lcell_comb \Selector2~9 (
// Equation(s):
// \Selector2~9_combout  = (\Selector2~2_combout ) # ((\Selector2~3_combout ) # (\Selector2~8_combout ))

	.dataa(gnd),
	.datab(\Selector2~2_combout ),
	.datac(\Selector2~3_combout ),
	.datad(\Selector2~8_combout ),
	.cin(gnd),
	.combout(\Selector2~9_combout ),
	.cout());
// synopsys translate_off
defparam \Selector2~9 .lut_mask = 16'hFFFC;
defparam \Selector2~9 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X50_Y37_N12
cycloneive_lcell_comb \Selector3~10 (
// Equation(s):
// \Selector3~10_combout  = (\Add0~56_combout  & \Selector0~9_combout )

	.dataa(gnd),
	.datab(gnd),
	.datac(\Add0~56_combout ),
	.datad(\Selector0~9_combout ),
	.cin(gnd),
	.combout(\Selector3~10_combout ),
	.cout());
// synopsys translate_off
defparam \Selector3~10 .lut_mask = 16'hF000;
defparam \Selector3~10 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X50_Y39_N24
cycloneive_lcell_comb \Selector3~3 (
// Equation(s):
// \Selector3~3_combout  = (\porta~107_combout  & (\Selector0~10_combout )) # (!\porta~107_combout  & (((!\portb~10_combout  & \Selector0~12_combout ))))

	.dataa(porta23),
	.datab(\Selector0~10_combout ),
	.datac(portb3),
	.datad(\Selector0~12_combout ),
	.cin(gnd),
	.combout(\Selector3~3_combout ),
	.cout());
// synopsys translate_off
defparam \Selector3~3 .lut_mask = 16'h8D88;
defparam \Selector3~3 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X50_Y39_N26
cycloneive_lcell_comb \Selector3~4 (
// Equation(s):
// \Selector3~4_combout  = (\Selector3~3_combout ) # ((\Selector0~13_combout  & (\portb~10_combout  $ (\porta~107_combout ))))

	.dataa(portb3),
	.datab(\Selector3~3_combout ),
	.datac(\Selector0~13_combout ),
	.datad(porta23),
	.cin(gnd),
	.combout(\Selector3~4_combout ),
	.cout());
// synopsys translate_off
defparam \Selector3~4 .lut_mask = 16'hDCEC;
defparam \Selector3~4 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X50_Y39_N2
cycloneive_lcell_comb \Selector3~2 (
// Equation(s):
// \Selector3~2_combout  = (\portb~10_combout  & ((\Selector0~10_combout ) # ((\porta~107_combout  & \Selector0~11_combout ))))

	.dataa(porta23),
	.datab(\Selector0~10_combout ),
	.datac(portb3),
	.datad(\Selector0~11_combout ),
	.cin(gnd),
	.combout(\Selector3~2_combout ),
	.cout());
// synopsys translate_off
defparam \Selector3~2 .lut_mask = 16'hE0C0;
defparam \Selector3~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X50_Y39_N4
cycloneive_lcell_comb \Selector3~5 (
// Equation(s):
// \Selector3~5_combout  = (\Selector1~4_combout  & ((\portb~64_combout  & (\ShiftLeft0~14_combout )) # (!\portb~64_combout  & ((\Selector11~0_combout )))))

	.dataa(portb30),
	.datab(\ShiftLeft0~14_combout ),
	.datac(\Selector11~0_combout ),
	.datad(\Selector1~4_combout ),
	.cin(gnd),
	.combout(\Selector3~5_combout ),
	.cout());
// synopsys translate_off
defparam \Selector3~5 .lut_mask = 16'hD800;
defparam \Selector3~5 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X50_Y37_N22
cycloneive_lcell_comb \Selector3~6 (
// Equation(s):
// \Selector3~6_combout  = (\Selector3~1_combout  & (((!\ShiftRight0~74_combout )))) # (!\Selector3~1_combout  & ((\ShiftRight0~74_combout  & (\ShiftLeft0~79_combout )) # (!\ShiftRight0~74_combout  & ((\ShiftLeft0~73_combout )))))

	.dataa(\ShiftLeft0~79_combout ),
	.datab(\Selector3~1_combout ),
	.datac(\ShiftLeft0~73_combout ),
	.datad(\ShiftRight0~74_combout ),
	.cin(gnd),
	.combout(\Selector3~6_combout ),
	.cout());
// synopsys translate_off
defparam \Selector3~6 .lut_mask = 16'h22FC;
defparam \Selector3~6 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y40_N8
cycloneive_lcell_comb \ShiftLeft0~65 (
// Equation(s):
// \ShiftLeft0~65_combout  = (\portb~62_combout  & (\ShiftLeft0~52_combout )) # (!\portb~62_combout  & ((\ShiftLeft0~64_combout )))

	.dataa(gnd),
	.datab(portb29),
	.datac(\ShiftLeft0~52_combout ),
	.datad(\ShiftLeft0~64_combout ),
	.cin(gnd),
	.combout(\ShiftLeft0~65_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftLeft0~65 .lut_mask = 16'hF3C0;
defparam \ShiftLeft0~65 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X50_Y37_N8
cycloneive_lcell_comb \Selector3~7 (
// Equation(s):
// \Selector3~7_combout  = (\Selector3~1_combout  & ((\Selector3~6_combout  & ((\ShiftLeft0~65_combout ))) # (!\Selector3~6_combout  & (\ShiftLeft0~76_combout )))) # (!\Selector3~1_combout  & (((\Selector3~6_combout ))))

	.dataa(\ShiftLeft0~76_combout ),
	.datab(\Selector3~1_combout ),
	.datac(\Selector3~6_combout ),
	.datad(\ShiftLeft0~65_combout ),
	.cin(gnd),
	.combout(\Selector3~7_combout ),
	.cout());
// synopsys translate_off
defparam \Selector3~7 .lut_mask = 16'hF838;
defparam \Selector3~7 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X50_Y37_N14
cycloneive_lcell_comb \Selector3~8 (
// Equation(s):
// \Selector3~8_combout  = (\ShiftRight0~59_combout  & ((\Selector2~4_combout ) # ((\Selector3~7_combout  & \Selector2~5_combout )))) # (!\ShiftRight0~59_combout  & (((\Selector3~7_combout  & \Selector2~5_combout ))))

	.dataa(\ShiftRight0~59_combout ),
	.datab(\Selector2~4_combout ),
	.datac(\Selector3~7_combout ),
	.datad(\Selector2~5_combout ),
	.cin(gnd),
	.combout(\Selector3~8_combout ),
	.cout());
// synopsys translate_off
defparam \Selector3~8 .lut_mask = 16'hF888;
defparam \Selector3~8 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X50_Y39_N18
cycloneive_lcell_comb \Selector3~9 (
// Equation(s):
// \Selector3~9_combout  = (\Selector3~4_combout ) # ((\Selector3~2_combout ) # ((\Selector3~5_combout ) # (\Selector3~8_combout )))

	.dataa(\Selector3~4_combout ),
	.datab(\Selector3~2_combout ),
	.datac(\Selector3~5_combout ),
	.datad(\Selector3~8_combout ),
	.cin(gnd),
	.combout(\Selector3~9_combout ),
	.cout());
// synopsys translate_off
defparam \Selector3~9 .lut_mask = 16'hFFFE;
defparam \Selector3~9 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X52_Y42_N28
cycloneive_lcell_comb \Selector0~23 (
// Equation(s):
// \Selector0~23_combout  = (\Selector0~13_combout  & (\porta~104_combout  $ (\portb~4_combout )))

	.dataa(porta20),
	.datab(\Selector0~13_combout ),
	.datac(gnd),
	.datad(portb),
	.cin(gnd),
	.combout(\Selector0~23_combout ),
	.cout());
// synopsys translate_off
defparam \Selector0~23 .lut_mask = 16'h4488;
defparam \Selector0~23 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y42_N12
cycloneive_lcell_comb \Selector0~24 (
// Equation(s):
// \Selector0~24_combout  = (\Selector0~10_combout  & \portb~4_combout )

	.dataa(gnd),
	.datab(gnd),
	.datac(\Selector0~10_combout ),
	.datad(portb),
	.cin(gnd),
	.combout(\Selector0~24_combout ),
	.cout());
// synopsys translate_off
defparam \Selector0~24 .lut_mask = 16'hF000;
defparam \Selector0~24 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X52_Y37_N28
cycloneive_lcell_comb \Add0~60 (
// Equation(s):
// \Add0~60_combout  = ((\portb~6_combout  $ (\porta~106_combout  $ (!\Add0~59 )))) # (GND)
// \Add0~61  = CARRY((\portb~6_combout  & ((\porta~106_combout ) # (!\Add0~59 ))) # (!\portb~6_combout  & (\porta~106_combout  & !\Add0~59 )))

	.dataa(portb1),
	.datab(porta22),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add0~59 ),
	.combout(\Add0~60_combout ),
	.cout(\Add0~61 ));
// synopsys translate_off
defparam \Add0~60 .lut_mask = 16'h698E;
defparam \Add0~60 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X52_Y37_N30
cycloneive_lcell_comb \Add0~62 (
// Equation(s):
// \Add0~62_combout  = \porta~104_combout  $ (\Add0~61  $ (\portb~4_combout ))

	.dataa(porta20),
	.datab(gnd),
	.datac(gnd),
	.datad(portb),
	.cin(\Add0~61 ),
	.combout(\Add0~62_combout ),
	.cout());
// synopsys translate_off
defparam \Add0~62 .lut_mask = 16'hA55A;
defparam \Add0~62 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X52_Y42_N2
cycloneive_lcell_comb \Selector0~25 (
// Equation(s):
// \Selector0~25_combout  = (\Selector0~19_combout  & ((\portb~62_combout  & ((\ShiftLeft0~55_combout ))) # (!\portb~62_combout  & (\ShiftLeft0~67_combout ))))

	.dataa(\Selector0~19_combout ),
	.datab(portb29),
	.datac(\ShiftLeft0~67_combout ),
	.datad(\ShiftLeft0~55_combout ),
	.cin(gnd),
	.combout(\Selector0~25_combout ),
	.cout());
// synopsys translate_off
defparam \Selector0~25 .lut_mask = 16'hA820;
defparam \Selector0~25 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X52_Y42_N8
cycloneive_lcell_comb \Selector0~26 (
// Equation(s):
// \Selector0~26_combout  = (\Selector0~24_combout ) # ((\Selector0~25_combout ) # ((\Selector0~9_combout  & \Add0~62_combout )))

	.dataa(\Selector0~24_combout ),
	.datab(\Selector0~9_combout ),
	.datac(\Add0~62_combout ),
	.datad(\Selector0~25_combout ),
	.cin(gnd),
	.combout(\Selector0~26_combout ),
	.cout());
// synopsys translate_off
defparam \Selector0~26 .lut_mask = 16'hFFEA;
defparam \Selector0~26 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y41_N8
cycloneive_lcell_comb \Selector0~27 (
// Equation(s):
// \Selector0~27_combout  = (\Selector0~10_combout ) # ((\portb~4_combout  & \Selector0~11_combout ))

	.dataa(portb),
	.datab(\Selector0~10_combout ),
	.datac(gnd),
	.datad(\Selector0~11_combout ),
	.cin(gnd),
	.combout(\Selector0~27_combout ),
	.cout());
// synopsys translate_off
defparam \Selector0~27 .lut_mask = 16'hEECC;
defparam \Selector0~27 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y41_N16
cycloneive_lcell_comb \Selector0~28 (
// Equation(s):
// \Selector0~28_combout  = (\porta~104_combout  & ((\Selector0~27_combout ) # ((\Selector8~1_combout  & !\ShiftRight0~71_combout ))))

	.dataa(porta20),
	.datab(\Selector0~27_combout ),
	.datac(\Selector8~1_combout ),
	.datad(\ShiftRight0~71_combout ),
	.cin(gnd),
	.combout(\Selector0~28_combout ),
	.cout());
// synopsys translate_off
defparam \Selector0~28 .lut_mask = 16'h88A8;
defparam \Selector0~28 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y41_N14
cycloneive_lcell_comb \Selector0~29 (
// Equation(s):
// \Selector0~29_combout  = (\Selector0~28_combout ) # ((!\porta~104_combout  & (\Selector0~12_combout  & !\portb~4_combout )))

	.dataa(porta20),
	.datab(\Selector0~12_combout ),
	.datac(portb),
	.datad(\Selector0~28_combout ),
	.cin(gnd),
	.combout(\Selector0~29_combout ),
	.cout());
// synopsys translate_off
defparam \Selector0~29 .lut_mask = 16'hFF04;
defparam \Selector0~29 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y39_N28
cycloneive_lcell_comb \Add1~60 (
// Equation(s):
// \Add1~60_combout  = ((\porta~106_combout  $ (\portb~6_combout  $ (\Add1~59 )))) # (GND)
// \Add1~61  = CARRY((\porta~106_combout  & ((!\Add1~59 ) # (!\portb~6_combout ))) # (!\porta~106_combout  & (!\portb~6_combout  & !\Add1~59 )))

	.dataa(porta22),
	.datab(portb1),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add1~59 ),
	.combout(\Add1~60_combout ),
	.cout(\Add1~61 ));
// synopsys translate_off
defparam \Add1~60 .lut_mask = 16'h962B;
defparam \Add1~60 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X57_Y39_N30
cycloneive_lcell_comb \Add1~62 (
// Equation(s):
// \Add1~62_combout  = \portb~4_combout  $ (\Add1~61  $ (!\porta~104_combout ))

	.dataa(gnd),
	.datab(portb),
	.datac(gnd),
	.datad(porta20),
	.cin(\Add1~61 ),
	.combout(\Add1~62_combout ),
	.cout());
// synopsys translate_off
defparam \Add1~62 .lut_mask = 16'h3CC3;
defparam \Add1~62 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X52_Y42_N6
cycloneive_lcell_comb \Selector1~6 (
// Equation(s):
// \Selector1~6_combout  = (\portb~62_combout ) # ((\portb~58_combout  & !\portb~60_combout ))

	.dataa(portb29),
	.datab(gnd),
	.datac(portb27),
	.datad(portb28),
	.cin(gnd),
	.combout(\Selector1~6_combout ),
	.cout());
// synopsys translate_off
defparam \Selector1~6 .lut_mask = 16'hAAFA;
defparam \Selector1~6 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X52_Y42_N16
cycloneive_lcell_comb \Selector0~30 (
// Equation(s):
// \Selector0~30_combout  = (\Selector1~0_combout  & (((\ShiftLeft0~78_combout ) # (\Selector1~6_combout )))) # (!\Selector1~0_combout  & (\porta~104_combout  & ((!\Selector1~6_combout ))))

	.dataa(porta20),
	.datab(\ShiftLeft0~78_combout ),
	.datac(\Selector1~0_combout ),
	.datad(\Selector1~6_combout ),
	.cin(gnd),
	.combout(\Selector0~30_combout ),
	.cout());
// synopsys translate_off
defparam \Selector0~30 .lut_mask = 16'hF0CA;
defparam \Selector0~30 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X52_Y42_N14
cycloneive_lcell_comb \Selector0~31 (
// Equation(s):
// \Selector0~31_combout  = (\Selector1~6_combout  & ((\Selector0~30_combout  & (\ShiftLeft0~75_combout )) # (!\Selector0~30_combout  & ((\porta~106_combout ))))) # (!\Selector1~6_combout  & (((\Selector0~30_combout ))))

	.dataa(\Selector1~6_combout ),
	.datab(\ShiftLeft0~75_combout ),
	.datac(porta22),
	.datad(\Selector0~30_combout ),
	.cin(gnd),
	.combout(\Selector0~31_combout ),
	.cout());
// synopsys translate_off
defparam \Selector0~31 .lut_mask = 16'hDDA0;
defparam \Selector0~31 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X52_Y42_N12
cycloneive_lcell_comb \Selector0~32 (
// Equation(s):
// \Selector0~32_combout  = (\Selector0~15_combout  & (\Selector0~31_combout  & (!\Selector1~2_combout  & !plif_idexaluop_l_0)))

	.dataa(\Selector0~15_combout ),
	.datab(\Selector0~31_combout ),
	.datac(\Selector1~2_combout ),
	.datad(plif_idexaluop_l_0),
	.cin(gnd),
	.combout(\Selector0~32_combout ),
	.cout());
// synopsys translate_off
defparam \Selector0~32 .lut_mask = 16'h0008;
defparam \Selector0~32 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X52_Y42_N26
cycloneive_lcell_comb \Selector0~33 (
// Equation(s):
// \Selector0~33_combout  = (\Selector0~29_combout ) # ((\Selector0~32_combout ) # ((\Selector0~8_combout  & \Add1~62_combout )))

	.dataa(\Selector0~29_combout ),
	.datab(\Selector0~8_combout ),
	.datac(\Add1~62_combout ),
	.datad(\Selector0~32_combout ),
	.cin(gnd),
	.combout(\Selector0~33_combout ),
	.cout());
// synopsys translate_off
defparam \Selector0~33 .lut_mask = 16'hFFEA;
defparam \Selector0~33 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X52_Y35_N12
cycloneive_lcell_comb \Selector0~22 (
// Equation(s):
// \Selector0~22_combout  = (!plif_idexaluop_l_0 & (\portb~66_combout  & (\ShiftLeft0~44_combout  & \Selector1~3_combout )))

	.dataa(plif_idexaluop_l_0),
	.datab(portb31),
	.datac(\ShiftLeft0~44_combout ),
	.datad(\Selector1~3_combout ),
	.cin(gnd),
	.combout(\Selector0~22_combout ),
	.cout());
// synopsys translate_off
defparam \Selector0~22 .lut_mask = 16'h4000;
defparam \Selector0~22 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y42_N26
cycloneive_lcell_comb \Selector1~7 (
// Equation(s):
// \Selector1~7_combout  = (\ShiftRight0~57_combout  & (!\portb~64_combout  & (!\Selector1~0_combout  & \Selector8~1_combout )))

	.dataa(\ShiftRight0~57_combout ),
	.datab(portb30),
	.datac(\Selector1~0_combout ),
	.datad(\Selector8~1_combout ),
	.cin(gnd),
	.combout(\Selector1~7_combout ),
	.cout());
// synopsys translate_off
defparam \Selector1~7 .lut_mask = 16'h0200;
defparam \Selector1~7 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y42_N18
cycloneive_lcell_comb \Selector1~8 (
// Equation(s):
// \Selector1~8_combout  = (\Selector1~7_combout ) # ((\Selector0~13_combout  & (\portb~6_combout  $ (\porta~106_combout ))))

	.dataa(\Selector0~13_combout ),
	.datab(portb1),
	.datac(porta22),
	.datad(\Selector1~7_combout ),
	.cin(gnd),
	.combout(\Selector1~8_combout ),
	.cout());
// synopsys translate_off
defparam \Selector1~8 .lut_mask = 16'hFF28;
defparam \Selector1~8 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X52_Y35_N6
cycloneive_lcell_comb \Selector1~18 (
// Equation(s):
// \Selector1~18_combout  = (\portb~6_combout  & ((\Selector0~10_combout ) # ((\Selector0~11_combout  & \porta~106_combout ))))

	.dataa(\Selector0~10_combout ),
	.datab(portb1),
	.datac(\Selector0~11_combout ),
	.datad(porta22),
	.cin(gnd),
	.combout(\Selector1~18_combout ),
	.cout());
// synopsys translate_off
defparam \Selector1~18 .lut_mask = 16'hC888;
defparam \Selector1~18 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y42_N18
cycloneive_lcell_comb \Selector1~9 (
// Equation(s):
// \Selector1~9_combout  = (\porta~106_combout  & (\Selector0~10_combout )) # (!\porta~106_combout  & (((!\portb~6_combout  & \Selector0~12_combout ))))

	.dataa(\Selector0~10_combout ),
	.datab(porta22),
	.datac(portb1),
	.datad(\Selector0~12_combout ),
	.cin(gnd),
	.combout(\Selector1~9_combout ),
	.cout());
// synopsys translate_off
defparam \Selector1~9 .lut_mask = 16'h8B88;
defparam \Selector1~9 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X52_Y42_N18
cycloneive_lcell_comb \Selector1~10 (
// Equation(s):
// \Selector1~10_combout  = (\Selector1~0_combout  & ((\ShiftLeft0~79_combout ) # ((\Selector1~6_combout )))) # (!\Selector1~0_combout  & (((\porta~106_combout  & !\Selector1~6_combout ))))

	.dataa(\ShiftLeft0~79_combout ),
	.datab(porta22),
	.datac(\Selector1~0_combout ),
	.datad(\Selector1~6_combout ),
	.cin(gnd),
	.combout(\Selector1~10_combout ),
	.cout());
// synopsys translate_off
defparam \Selector1~10 .lut_mask = 16'hF0AC;
defparam \Selector1~10 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X52_Y42_N22
cycloneive_lcell_comb \Selector1~14 (
// Equation(s):
// \Selector1~14_combout  = (plif_idexaluop_l_0 & ((\Selector1~10_combout ))) # (!plif_idexaluop_l_0 & (\porta~105_combout  & !\Selector1~10_combout ))

	.dataa(porta21),
	.datab(plif_idexaluop_l_0),
	.datac(gnd),
	.datad(\Selector1~10_combout ),
	.cin(gnd),
	.combout(\Selector1~14_combout ),
	.cout());
// synopsys translate_off
defparam \Selector1~14 .lut_mask = 16'hCC22;
defparam \Selector1~14 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y42_N26
cycloneive_lcell_comb \Selector1~15 (
// Equation(s):
// \Selector1~15_combout  = (\Selector1~10_combout  & (!\Selector1~14_combout  & ((\ShiftLeft0~77_combout ) # (!\Selector1~6_combout )))) # (!\Selector1~10_combout  & (\Selector1~6_combout  & ((\Selector1~14_combout ))))

	.dataa(\Selector1~6_combout ),
	.datab(\ShiftLeft0~77_combout ),
	.datac(\Selector1~10_combout ),
	.datad(\Selector1~14_combout ),
	.cin(gnd),
	.combout(\Selector1~15_combout ),
	.cout());
// synopsys translate_off
defparam \Selector1~15 .lut_mask = 16'h0AD0;
defparam \Selector1~15 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y42_N0
cycloneive_lcell_comb \Selector1~16 (
// Equation(s):
// \Selector1~16_combout  = (\Selector0~18_combout  & ((\Selector1~15_combout ) # ((\Selector0~19_combout  & \Selector1~5_combout )))) # (!\Selector0~18_combout  & (\Selector0~19_combout  & ((\Selector1~5_combout ))))

	.dataa(\Selector0~18_combout ),
	.datab(\Selector0~19_combout ),
	.datac(\Selector1~15_combout ),
	.datad(\Selector1~5_combout ),
	.cin(gnd),
	.combout(\Selector1~16_combout ),
	.cout());
// synopsys translate_off
defparam \Selector1~16 .lut_mask = 16'hECA0;
defparam \Selector1~16 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X52_Y42_N20
cycloneive_lcell_comb \Selector1~11 (
// Equation(s):
// \Selector1~11_combout  = (\Selector1~6_combout  & ((\Selector1~10_combout  & ((\ShiftLeft0~77_combout ))) # (!\Selector1~10_combout  & (\porta~105_combout )))) # (!\Selector1~6_combout  & (\Selector1~10_combout ))

	.dataa(\Selector1~6_combout ),
	.datab(\Selector1~10_combout ),
	.datac(porta21),
	.datad(\ShiftLeft0~77_combout ),
	.cin(gnd),
	.combout(\Selector1~11_combout ),
	.cout());
// synopsys translate_off
defparam \Selector1~11 .lut_mask = 16'hEC64;
defparam \Selector1~11 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y42_N4
cycloneive_lcell_comb \Selector1~12 (
// Equation(s):
// \Selector1~12_combout  = (\Selector0~18_combout  & \Selector1~11_combout )

	.dataa(gnd),
	.datab(gnd),
	.datac(\Selector0~18_combout ),
	.datad(\Selector1~11_combout ),
	.cin(gnd),
	.combout(\Selector1~12_combout ),
	.cout());
// synopsys translate_off
defparam \Selector1~12 .lut_mask = 16'hF000;
defparam \Selector1~12 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y42_N0
cycloneive_lcell_comb \Selector1~13 (
// Equation(s):
// \Selector1~13_combout  = (!plif_idexaluop_l_0 & ((\Selector1~12_combout ) # ((\Selector1~3_combout  & \ShiftLeft0~47_combout ))))

	.dataa(plif_idexaluop_l_0),
	.datab(\Selector1~3_combout ),
	.datac(\Selector1~12_combout ),
	.datad(\ShiftLeft0~47_combout ),
	.cin(gnd),
	.combout(\Selector1~13_combout ),
	.cout());
// synopsys translate_off
defparam \Selector1~13 .lut_mask = 16'h5450;
defparam \Selector1~13 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y42_N20
cycloneive_lcell_comb \Selector1~17 (
// Equation(s):
// \Selector1~17_combout  = (\Selector1~9_combout ) # ((\Selector1~16_combout ) # ((\portb~66_combout  & \Selector1~13_combout )))

	.dataa(portb31),
	.datab(\Selector1~9_combout ),
	.datac(\Selector1~16_combout ),
	.datad(\Selector1~13_combout ),
	.cin(gnd),
	.combout(\Selector1~17_combout ),
	.cout());
// synopsys translate_off
defparam \Selector1~17 .lut_mask = 16'hFEFC;
defparam \Selector1~17 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y42_N12
cycloneive_lcell_comb \Selector1~19 (
// Equation(s):
// \Selector1~19_combout  = (\Selector1~18_combout ) # ((\Selector1~17_combout ) # ((\Selector0~8_combout  & \Add1~60_combout )))

	.dataa(\Selector0~8_combout ),
	.datab(\Selector1~18_combout ),
	.datac(\Add1~60_combout ),
	.datad(\Selector1~17_combout ),
	.cin(gnd),
	.combout(\Selector1~19_combout ),
	.cout());
// synopsys translate_off
defparam \Selector1~19 .lut_mask = 16'hFFEC;
defparam \Selector1~19 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X50_Y39_N10
cycloneive_lcell_comb \WideOr1~0 (
// Equation(s):
// \WideOr1~0_combout  = (Selector26) # ((Selector2) # ((Selector3) # (Selector27)))

	.dataa(Selector26),
	.datab(Selector2),
	.datac(Selector3),
	.datad(Selector27),
	.cin(gnd),
	.combout(\WideOr1~0_combout ),
	.cout());
// synopsys translate_off
defparam \WideOr1~0 .lut_mask = 16'hFFFE;
defparam \WideOr1~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X52_Y39_N16
cycloneive_lcell_comb \WideOr1~6 (
// Equation(s):
// \WideOr1~6_combout  = (\WideOr1~5_combout ) # ((Selector7) # ((Selector8) # (Selector9)))

	.dataa(\WideOr1~5_combout ),
	.datab(Selector7),
	.datac(Selector8),
	.datad(Selector9),
	.cin(gnd),
	.combout(\WideOr1~6_combout ),
	.cout());
// synopsys translate_off
defparam \WideOr1~6 .lut_mask = 16'hFFFE;
defparam \WideOr1~6 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y36_N6
cycloneive_lcell_comb \WideOr1~7 (
// Equation(s):
// \WideOr1~7_combout  = (Selector5) # ((Selector4) # (Selector6))

	.dataa(Selector5),
	.datab(gnd),
	.datac(Selector4),
	.datad(Selector6),
	.cin(gnd),
	.combout(\WideOr1~7_combout ),
	.cout());
// synopsys translate_off
defparam \WideOr1~7 .lut_mask = 16'hFFFA;
defparam \WideOr1~7 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y39_N4
cycloneive_lcell_comb \WideOr1~8 (
// Equation(s):
// \WideOr1~8_combout  = (Selector12) # (Selector11)

	.dataa(gnd),
	.datab(gnd),
	.datac(Selector12),
	.datad(Selector11),
	.cin(gnd),
	.combout(\WideOr1~8_combout ),
	.cout());
// synopsys translate_off
defparam \WideOr1~8 .lut_mask = 16'hFFF0;
defparam \WideOr1~8 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y39_N24
cycloneive_lcell_comb \WideOr1~9 (
// Equation(s):
// \WideOr1~9_combout  = (Selector22) # ((\WideOr1~8_combout ) # ((Selector23) # (Selector10)))

	.dataa(Selector22),
	.datab(\WideOr1~8_combout ),
	.datac(Selector23),
	.datad(Selector10),
	.cin(gnd),
	.combout(\WideOr1~9_combout ),
	.cout());
// synopsys translate_off
defparam \WideOr1~9 .lut_mask = 16'hFFFE;
defparam \WideOr1~9 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y39_N20
cycloneive_lcell_comb \WideOr1~10 (
// Equation(s):
// \WideOr1~10_combout  = (Selector13) # ((Selector25) # ((Selector14) # (\WideOr1~9_combout )))

	.dataa(Selector13),
	.datab(Selector25),
	.datac(Selector14),
	.datad(\WideOr1~9_combout ),
	.cin(gnd),
	.combout(\WideOr1~10_combout ),
	.cout());
// synopsys translate_off
defparam \WideOr1~10 .lut_mask = 16'hFFFE;
defparam \WideOr1~10 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y39_N20
cycloneive_lcell_comb \WideOr1~1 (
// Equation(s):
// \WideOr1~1_combout  = (Selector19) # ((Selector18) # ((Selector17) # (Selector20)))

	.dataa(Selector19),
	.datab(Selector18),
	.datac(Selector17),
	.datad(Selector20),
	.cin(gnd),
	.combout(\WideOr1~1_combout ),
	.cout());
// synopsys translate_off
defparam \WideOr1~1 .lut_mask = 16'hFFFE;
defparam \WideOr1~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y39_N26
cycloneive_lcell_comb \WideOr1~2 (
// Equation(s):
// \WideOr1~2_combout  = (\Selector31~7_combout ) # ((\Selector31~0_combout ) # ((\Selector31~4_combout ) # (\WideOr1~1_combout )))

	.dataa(\Selector31~7_combout ),
	.datab(\Selector31~0_combout ),
	.datac(\Selector31~4_combout ),
	.datad(\WideOr1~1_combout ),
	.cin(gnd),
	.combout(\WideOr1~2_combout ),
	.cout());
// synopsys translate_off
defparam \WideOr1~2 .lut_mask = 16'hFFFE;
defparam \WideOr1~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y39_N12
cycloneive_lcell_comb \WideOr1~3 (
// Equation(s):
// \WideOr1~3_combout  = (Selector16) # ((\WideOr1~2_combout ) # (Selector21))

	.dataa(Selector16),
	.datab(gnd),
	.datac(\WideOr1~2_combout ),
	.datad(Selector21),
	.cin(gnd),
	.combout(\WideOr1~3_combout ),
	.cout());
// synopsys translate_off
defparam \WideOr1~3 .lut_mask = 16'hFFFA;
defparam \WideOr1~3 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y39_N10
cycloneive_lcell_comb \WideOr1~4 (
// Equation(s):
// \WideOr1~4_combout  = (\Selector31~2_combout ) # ((Selector15) # ((Selector30) # (\WideOr1~3_combout )))

	.dataa(\Selector31~2_combout ),
	.datab(Selector15),
	.datac(Selector30),
	.datad(\WideOr1~3_combout ),
	.cin(gnd),
	.combout(\WideOr1~4_combout ),
	.cout());
// synopsys translate_off
defparam \WideOr1~4 .lut_mask = 16'hFFFE;
defparam \WideOr1~4 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y39_N0
cycloneive_lcell_comb \WideOr1~11 (
// Equation(s):
// \WideOr1~11_combout  = (\WideOr1~6_combout ) # ((\WideOr1~7_combout ) # ((\WideOr1~10_combout ) # (\WideOr1~4_combout )))

	.dataa(\WideOr1~6_combout ),
	.datab(\WideOr1~7_combout ),
	.datac(\WideOr1~10_combout ),
	.datad(\WideOr1~4_combout ),
	.cin(gnd),
	.combout(\WideOr1~11_combout ),
	.cout());
// synopsys translate_off
defparam \WideOr1~11 .lut_mask = 16'hFFFE;
defparam \WideOr1~11 .sum_lutc_input = "datac";
// synopsys translate_on

endmodule

module control_unit (
	plif_ifidinstr_l_31,
	plif_ifidinstr_l_29,
	plif_ifidinstr_l_27,
	plif_ifidinstr_l_26,
	plif_ifidinstr_l_28,
	Equal16,
	plif_ifidinstr_l_30,
	Equal22,
	plif_ifidinstr_l_5,
	plif_ifidinstr_l_1,
	plif_ifidinstr_l_0,
	plif_ifidinstr_l_2,
	plif_ifidinstr_l_3,
	WideNor0,
	Equal11,
	Equal26,
	plif_ifidinstr_l_4,
	Equal21,
	WideOr141,
	Equal13,
	aluop_l,
	WideNor1,
	Selector22,
	Selector4,
	plif_ifidinstr_l_22,
	Selector41,
	plif_ifidinstr_l_21,
	Selector5,
	plif_ifidinstr_l_24,
	Selector2,
	plif_ifidinstr_l_23,
	Selector3,
	plif_ifidinstr_l_25,
	Selector1,
	Equal6,
	Selector11,
	Selector21,
	Selector9,
	plif_ifidinstr_l_17,
	Selector91,
	plif_ifidinstr_l_16,
	Selector10,
	plif_ifidinstr_l_19,
	Selector7,
	plif_ifidinstr_l_18,
	Selector8,
	plif_ifidinstr_l_20,
	Selector6,
	Equal23,
	pcsrc,
	Equal1,
	Equal20,
	WideNor11,
	Equal19,
	Equal12,
	Equal18,
	Selector221,
	WideOr142,
	WideOr151,
	WideOr161,
	plif_ifidinstr_l_10,
	plif_ifidinstr_l_9,
	plif_ifidinstr_l_8,
	plif_ifidinstr_l_7,
	plif_ifidinstr_l_6,
	Selector14,
	Selector15,
	Selector16,
	Selector17,
	Selector18,
	Selector24,
	Equal121,
	Selector0,
	Equal25,
	devpor,
	devclrn,
	devoe);
input 	plif_ifidinstr_l_31;
input 	plif_ifidinstr_l_29;
input 	plif_ifidinstr_l_27;
input 	plif_ifidinstr_l_26;
input 	plif_ifidinstr_l_28;
output 	Equal16;
input 	plif_ifidinstr_l_30;
output 	Equal22;
input 	plif_ifidinstr_l_5;
input 	plif_ifidinstr_l_1;
input 	plif_ifidinstr_l_0;
input 	plif_ifidinstr_l_2;
input 	plif_ifidinstr_l_3;
output 	WideNor0;
output 	Equal11;
output 	Equal26;
input 	plif_ifidinstr_l_4;
output 	Equal21;
output 	WideOr141;
output 	Equal13;
input 	aluop_l;
output 	WideNor1;
output 	Selector22;
output 	Selector4;
input 	plif_ifidinstr_l_22;
output 	Selector41;
input 	plif_ifidinstr_l_21;
output 	Selector5;
input 	plif_ifidinstr_l_24;
output 	Selector2;
input 	plif_ifidinstr_l_23;
output 	Selector3;
input 	plif_ifidinstr_l_25;
output 	Selector1;
output 	Equal6;
output 	Selector11;
output 	Selector21;
output 	Selector9;
input 	plif_ifidinstr_l_17;
output 	Selector91;
input 	plif_ifidinstr_l_16;
output 	Selector10;
input 	plif_ifidinstr_l_19;
output 	Selector7;
input 	plif_ifidinstr_l_18;
output 	Selector8;
input 	plif_ifidinstr_l_20;
output 	Selector6;
output 	Equal23;
output 	pcsrc;
output 	Equal1;
output 	Equal20;
output 	WideNor11;
output 	Equal19;
output 	Equal12;
output 	Equal18;
output 	Selector221;
output 	WideOr142;
output 	WideOr151;
output 	WideOr161;
input 	plif_ifidinstr_l_10;
input 	plif_ifidinstr_l_9;
input 	plif_ifidinstr_l_8;
input 	plif_ifidinstr_l_7;
input 	plif_ifidinstr_l_6;
output 	Selector14;
output 	Selector15;
output 	Selector16;
output 	Selector17;
output 	Selector18;
output 	Selector24;
output 	Equal121;
output 	Selector0;
output 	Equal25;

// Design Ports Information

input 	devpor;
input 	devclrn;
input 	devoe;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
assign unknown = 1'bx;

wire \Equal13~0_combout ;
wire \WideNor0~1_combout ;
wire \WideNor0~0_combout ;
wire \WideNor0~3_combout ;
wire \Selector5~0_combout ;
wire \WideOr15~0_combout ;
wire \Selector22~3_combout ;
wire \Selector22~8_combout ;
wire \WideOr16~combout ;


// Location: LCCOMB_X59_Y30_N28
cycloneive_lcell_comb \Equal16~0 (
// Equation(s):
// Equal16 = (plif_ifidinstr_l_27 & (!plif_ifidinstr_l_28 & plif_ifidinstr_l_26))

	.dataa(plif_ifidinstr_l_27),
	.datab(gnd),
	.datac(plif_ifidinstr_l_28),
	.datad(plif_ifidinstr_l_26),
	.cin(gnd),
	.combout(Equal16),
	.cout());
// synopsys translate_off
defparam \Equal16~0 .lut_mask = 16'h0A00;
defparam \Equal16~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y30_N0
cycloneive_lcell_comb \Equal22~0 (
// Equation(s):
// Equal22 = (plif_ifidinstr_l_31 & (plif_ifidinstr_l_29 & (!plif_ifidinstr_l_30 & Equal16)))

	.dataa(plif_ifidinstr_l_31),
	.datab(plif_ifidinstr_l_29),
	.datac(plif_ifidinstr_l_30),
	.datad(Equal16),
	.cin(gnd),
	.combout(Equal22),
	.cout());
// synopsys translate_off
defparam \Equal22~0 .lut_mask = 16'h0800;
defparam \Equal22~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y30_N2
cycloneive_lcell_comb \WideNor0~2 (
// Equation(s):
// WideNor0 = (plif_ifidinstr_l_3 & plif_ifidinstr_l_1)

	.dataa(gnd),
	.datab(gnd),
	.datac(plif_ifidinstr_l_3),
	.datad(plif_ifidinstr_l_1),
	.cin(gnd),
	.combout(WideNor0),
	.cout());
// synopsys translate_off
defparam \WideNor0~2 .lut_mask = 16'hF000;
defparam \WideNor0~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y30_N14
cycloneive_lcell_comb \Equal11~0 (
// Equation(s):
// Equal11 = (!plif_ifidinstr_l_29 & (!plif_ifidinstr_l_30 & !plif_ifidinstr_l_31))

	.dataa(gnd),
	.datab(plif_ifidinstr_l_29),
	.datac(plif_ifidinstr_l_30),
	.datad(plif_ifidinstr_l_31),
	.cin(gnd),
	.combout(Equal11),
	.cout());
// synopsys translate_off
defparam \Equal11~0 .lut_mask = 16'h0003;
defparam \Equal11~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y30_N26
cycloneive_lcell_comb \Equal26~0 (
// Equation(s):
// Equal26 = (!plif_ifidinstr_l_28 & (!plif_ifidinstr_l_26 & (!plif_ifidinstr_l_27 & Equal11)))

	.dataa(plif_ifidinstr_l_28),
	.datab(plif_ifidinstr_l_26),
	.datac(plif_ifidinstr_l_27),
	.datad(Equal11),
	.cin(gnd),
	.combout(Equal26),
	.cout());
// synopsys translate_off
defparam \Equal26~0 .lut_mask = 16'h0100;
defparam \Equal26~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y30_N22
cycloneive_lcell_comb \Equal21~0 (
// Equation(s):
// Equal21 = (plif_ifidinstr_l_31 & (!plif_ifidinstr_l_29 & (!plif_ifidinstr_l_30 & Equal16)))

	.dataa(plif_ifidinstr_l_31),
	.datab(plif_ifidinstr_l_29),
	.datac(plif_ifidinstr_l_30),
	.datad(Equal16),
	.cin(gnd),
	.combout(Equal21),
	.cout());
// synopsys translate_off
defparam \Equal21~0 .lut_mask = 16'h0200;
defparam \Equal21~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y30_N12
cycloneive_lcell_comb \WideOr14~0 (
// Equation(s):
// WideOr141 = (!Equal21 & (((plif_ifidinstr_l_27 & plif_ifidinstr_l_26)) # (!\Equal13~0_combout )))

	.dataa(plif_ifidinstr_l_27),
	.datab(plif_ifidinstr_l_26),
	.datac(Equal21),
	.datad(\Equal13~0_combout ),
	.cin(gnd),
	.combout(WideOr141),
	.cout());
// synopsys translate_off
defparam \WideOr14~0 .lut_mask = 16'h080F;
defparam \WideOr14~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y30_N26
cycloneive_lcell_comb \Equal13~1 (
// Equation(s):
// Equal13 = (plif_ifidinstr_l_29 & (!plif_ifidinstr_l_30 & !plif_ifidinstr_l_31))

	.dataa(gnd),
	.datab(plif_ifidinstr_l_29),
	.datac(plif_ifidinstr_l_30),
	.datad(plif_ifidinstr_l_31),
	.cin(gnd),
	.combout(Equal13),
	.cout());
// synopsys translate_off
defparam \Equal13~1 .lut_mask = 16'h000C;
defparam \Equal13~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y30_N18
cycloneive_lcell_comb \WideNor1~0 (
// Equation(s):
// WideNor1 = (aluop_l & (WideOr141 & ((!Equal16) # (!Equal13))))

	.dataa(Equal13),
	.datab(Equal16),
	.datac(aluop_l),
	.datad(WideOr141),
	.cin(gnd),
	.combout(WideNor1),
	.cout());
// synopsys translate_off
defparam \WideNor1~0 .lut_mask = 16'h7000;
defparam \WideNor1~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y30_N16
cycloneive_lcell_comb \Selector22~6 (
// Equation(s):
// Selector22 = ((plif_ifidinstr_l_27) # (!Equal11)) # (!plif_ifidinstr_l_28)

	.dataa(gnd),
	.datab(plif_ifidinstr_l_28),
	.datac(Equal11),
	.datad(plif_ifidinstr_l_27),
	.cin(gnd),
	.combout(Selector22),
	.cout());
// synopsys translate_off
defparam \Selector22~6 .lut_mask = 16'hFF3F;
defparam \Selector22~6 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y30_N30
cycloneive_lcell_comb \Selector4~0 (
// Equation(s):
// Selector4 = (Equal22) # ((\Selector5~0_combout ) # ((!WideNor1) # (!Selector22)))

	.dataa(Equal22),
	.datab(\Selector5~0_combout ),
	.datac(Selector22),
	.datad(WideNor1),
	.cin(gnd),
	.combout(Selector4),
	.cout());
// synopsys translate_off
defparam \Selector4~0 .lut_mask = 16'hEFFF;
defparam \Selector4~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y33_N26
cycloneive_lcell_comb \Selector4~1 (
// Equation(s):
// Selector41 = (Selector4 & plif_ifidinstr_l_22)

	.dataa(gnd),
	.datab(gnd),
	.datac(Selector4),
	.datad(plif_ifidinstr_l_22),
	.cin(gnd),
	.combout(Selector41),
	.cout());
// synopsys translate_off
defparam \Selector4~1 .lut_mask = 16'hF000;
defparam \Selector4~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X63_Y32_N24
cycloneive_lcell_comb \Selector5~1 (
// Equation(s):
// Selector5 = (plif_ifidinstr_l_21 & Selector4)

	.dataa(gnd),
	.datab(gnd),
	.datac(plif_ifidinstr_l_21),
	.datad(Selector4),
	.cin(gnd),
	.combout(Selector5),
	.cout());
// synopsys translate_off
defparam \Selector5~1 .lut_mask = 16'hF000;
defparam \Selector5~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y33_N16
cycloneive_lcell_comb \Selector2~0 (
// Equation(s):
// Selector2 = (Selector4 & plif_ifidinstr_l_24)

	.dataa(gnd),
	.datab(gnd),
	.datac(Selector4),
	.datad(plif_ifidinstr_l_24),
	.cin(gnd),
	.combout(Selector2),
	.cout());
// synopsys translate_off
defparam \Selector2~0 .lut_mask = 16'hF000;
defparam \Selector2~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y31_N12
cycloneive_lcell_comb \Selector3~0 (
// Equation(s):
// Selector3 = (plif_ifidinstr_l_23 & Selector4)

	.dataa(gnd),
	.datab(plif_ifidinstr_l_23),
	.datac(gnd),
	.datad(Selector4),
	.cin(gnd),
	.combout(Selector3),
	.cout());
// synopsys translate_off
defparam \Selector3~0 .lut_mask = 16'hCC00;
defparam \Selector3~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y32_N28
cycloneive_lcell_comb \Selector1~0 (
// Equation(s):
// Selector1 = (plif_ifidinstr_l_25 & Selector4)

	.dataa(plif_ifidinstr_l_25),
	.datab(gnd),
	.datac(gnd),
	.datad(Selector4),
	.cin(gnd),
	.combout(Selector1),
	.cout());
// synopsys translate_off
defparam \Selector1~0 .lut_mask = 16'hAA00;
defparam \Selector1~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y30_N20
cycloneive_lcell_comb \Equal6~0 (
// Equation(s):
// Equal6 = (!plif_ifidinstr_l_5 & (!plif_ifidinstr_l_2 & (!plif_ifidinstr_l_4 & !plif_ifidinstr_l_0)))

	.dataa(plif_ifidinstr_l_5),
	.datab(plif_ifidinstr_l_2),
	.datac(plif_ifidinstr_l_4),
	.datad(plif_ifidinstr_l_0),
	.cin(gnd),
	.combout(Equal6),
	.cout());
// synopsys translate_off
defparam \Equal6~0 .lut_mask = 16'h0001;
defparam \Equal6~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y30_N10
cycloneive_lcell_comb \Selector11~0 (
// Equation(s):
// Selector11 = (\Selector5~0_combout  & (((plif_ifidinstr_l_1) # (!Equal6)) # (!plif_ifidinstr_l_3)))

	.dataa(plif_ifidinstr_l_3),
	.datab(plif_ifidinstr_l_1),
	.datac(\Selector5~0_combout ),
	.datad(Equal6),
	.cin(gnd),
	.combout(Selector11),
	.cout());
// synopsys translate_off
defparam \Selector11~0 .lut_mask = 16'hD0F0;
defparam \Selector11~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y30_N0
cycloneive_lcell_comb \Selector21~0 (
// Equation(s):
// Selector21 = (plif_ifidinstr_l_3) # (!Equal6)

	.dataa(gnd),
	.datab(gnd),
	.datac(plif_ifidinstr_l_3),
	.datad(Equal6),
	.cin(gnd),
	.combout(Selector21),
	.cout());
// synopsys translate_off
defparam \Selector21~0 .lut_mask = 16'hF0FF;
defparam \Selector21~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y30_N22
cycloneive_lcell_comb \Selector9~0 (
// Equation(s):
// Selector9 = ((Equal22) # ((Selector21 & Selector11))) # (!Selector22)

	.dataa(Selector22),
	.datab(Selector21),
	.datac(Equal22),
	.datad(Selector11),
	.cin(gnd),
	.combout(Selector9),
	.cout());
// synopsys translate_off
defparam \Selector9~0 .lut_mask = 16'hFDF5;
defparam \Selector9~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y30_N28
cycloneive_lcell_comb \Selector9~1 (
// Equation(s):
// Selector91 = (plif_ifidinstr_l_17 & Selector9)

	.dataa(gnd),
	.datab(gnd),
	.datac(plif_ifidinstr_l_17),
	.datad(Selector9),
	.cin(gnd),
	.combout(Selector91),
	.cout());
// synopsys translate_off
defparam \Selector9~1 .lut_mask = 16'hF000;
defparam \Selector9~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y30_N14
cycloneive_lcell_comb \Selector10~0 (
// Equation(s):
// Selector10 = (plif_ifidinstr_l_16 & Selector9)

	.dataa(gnd),
	.datab(gnd),
	.datac(plif_ifidinstr_l_16),
	.datad(Selector9),
	.cin(gnd),
	.combout(Selector10),
	.cout());
// synopsys translate_off
defparam \Selector10~0 .lut_mask = 16'hF000;
defparam \Selector10~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y32_N16
cycloneive_lcell_comb \Selector7~0 (
// Equation(s):
// Selector7 = (plif_ifidinstr_l_19 & Selector9)

	.dataa(gnd),
	.datab(gnd),
	.datac(plif_ifidinstr_l_19),
	.datad(Selector9),
	.cin(gnd),
	.combout(Selector7),
	.cout());
// synopsys translate_off
defparam \Selector7~0 .lut_mask = 16'hF000;
defparam \Selector7~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y30_N4
cycloneive_lcell_comb \Selector8~0 (
// Equation(s):
// Selector8 = (plif_ifidinstr_l_18 & Selector9)

	.dataa(gnd),
	.datab(gnd),
	.datac(plif_ifidinstr_l_18),
	.datad(Selector9),
	.cin(gnd),
	.combout(Selector8),
	.cout());
// synopsys translate_off
defparam \Selector8~0 .lut_mask = 16'hF000;
defparam \Selector8~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y32_N6
cycloneive_lcell_comb \Selector6~0 (
// Equation(s):
// Selector6 = (plif_ifidinstr_l_20 & Selector9)

	.dataa(gnd),
	.datab(plif_ifidinstr_l_20),
	.datac(gnd),
	.datad(Selector9),
	.cin(gnd),
	.combout(Selector6),
	.cout());
// synopsys translate_off
defparam \Selector6~0 .lut_mask = 16'hCC00;
defparam \Selector6~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y29_N0
cycloneive_lcell_comb \Equal23~0 (
// Equation(s):
// Equal23 = (plif_ifidinstr_l_28 & (plif_ifidinstr_l_26 & (plif_ifidinstr_l_31 & plif_ifidinstr_l_27)))

	.dataa(plif_ifidinstr_l_28),
	.datab(plif_ifidinstr_l_26),
	.datac(plif_ifidinstr_l_31),
	.datad(plif_ifidinstr_l_27),
	.cin(gnd),
	.combout(Equal23),
	.cout());
// synopsys translate_off
defparam \Equal23~0 .lut_mask = 16'h8000;
defparam \Equal23~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y29_N24
cycloneive_lcell_comb \pcsrc~0 (
// Equation(s):
// pcsrc = ((plif_ifidinstr_l_28) # (!Equal11)) # (!plif_ifidinstr_l_27)

	.dataa(gnd),
	.datab(plif_ifidinstr_l_27),
	.datac(plif_ifidinstr_l_28),
	.datad(Equal11),
	.cin(gnd),
	.combout(pcsrc),
	.cout());
// synopsys translate_off
defparam \pcsrc~0 .lut_mask = 16'hF3FF;
defparam \pcsrc~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y30_N30
cycloneive_lcell_comb \Equal1~0 (
// Equation(s):
// Equal1 = (!plif_ifidinstr_l_4 & (plif_ifidinstr_l_5 & (plif_ifidinstr_l_2 & !plif_ifidinstr_l_3)))

	.dataa(plif_ifidinstr_l_4),
	.datab(plif_ifidinstr_l_5),
	.datac(plif_ifidinstr_l_2),
	.datad(plif_ifidinstr_l_3),
	.cin(gnd),
	.combout(Equal1),
	.cout());
// synopsys translate_off
defparam \Equal1~0 .lut_mask = 16'h0040;
defparam \Equal1~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y30_N20
cycloneive_lcell_comb \Equal20~0 (
// Equation(s):
// Equal20 = (plif_ifidinstr_l_28 & (Equal13 & (plif_ifidinstr_l_26 & plif_ifidinstr_l_27)))

	.dataa(plif_ifidinstr_l_28),
	.datab(Equal13),
	.datac(plif_ifidinstr_l_26),
	.datad(plif_ifidinstr_l_27),
	.cin(gnd),
	.combout(Equal20),
	.cout());
// synopsys translate_off
defparam \Equal20~0 .lut_mask = 16'h8000;
defparam \Equal20~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y33_N8
cycloneive_lcell_comb \WideNor1~1 (
// Equation(s):
// WideNor11 = (!Equal20 & (!Equal22 & (Selector22 & \WideOr15~0_combout )))

	.dataa(Equal20),
	.datab(Equal22),
	.datac(Selector22),
	.datad(\WideOr15~0_combout ),
	.cin(gnd),
	.combout(WideNor11),
	.cout());
// synopsys translate_off
defparam \WideNor1~1 .lut_mask = 16'h1000;
defparam \WideNor1~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y30_N2
cycloneive_lcell_comb \Equal19~0 (
// Equation(s):
// Equal19 = (plif_ifidinstr_l_28 & (Equal13 & (!plif_ifidinstr_l_26 & plif_ifidinstr_l_27)))

	.dataa(plif_ifidinstr_l_28),
	.datab(Equal13),
	.datac(plif_ifidinstr_l_26),
	.datad(plif_ifidinstr_l_27),
	.cin(gnd),
	.combout(Equal19),
	.cout());
// synopsys translate_off
defparam \Equal19~0 .lut_mask = 16'h0800;
defparam \Equal19~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y30_N16
cycloneive_lcell_comb \Equal1~1 (
// Equation(s):
// Equal12 = (Equal1 & !plif_ifidinstr_l_1)

	.dataa(Equal1),
	.datab(gnd),
	.datac(plif_ifidinstr_l_1),
	.datad(gnd),
	.cin(gnd),
	.combout(Equal12),
	.cout());
// synopsys translate_off
defparam \Equal1~1 .lut_mask = 16'h0A0A;
defparam \Equal1~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y30_N22
cycloneive_lcell_comb \Equal18~0 (
// Equation(s):
// Equal18 = (plif_ifidinstr_l_28 & (Equal13 & (plif_ifidinstr_l_26 & !plif_ifidinstr_l_27)))

	.dataa(plif_ifidinstr_l_28),
	.datab(Equal13),
	.datac(plif_ifidinstr_l_26),
	.datad(plif_ifidinstr_l_27),
	.cin(gnd),
	.combout(Equal18),
	.cout());
// synopsys translate_off
defparam \Equal18~0 .lut_mask = 16'h0080;
defparam \Equal18~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y30_N24
cycloneive_lcell_comb \Selector22~7 (
// Equation(s):
// Selector221 = (Equal26 & ((\Selector22~8_combout ) # ((Equal12 & plif_ifidinstr_l_0))))

	.dataa(\Selector22~8_combout ),
	.datab(Equal12),
	.datac(plif_ifidinstr_l_0),
	.datad(Equal26),
	.cin(gnd),
	.combout(Selector221),
	.cout());
// synopsys translate_off
defparam \Selector22~7 .lut_mask = 16'hEA00;
defparam \Selector22~7 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y33_N18
cycloneive_lcell_comb WideOr14(
// Equation(s):
// WideOr142 = (Equal22) # ((!WideOr141) # (!Selector22))

	.dataa(gnd),
	.datab(Equal22),
	.datac(Selector22),
	.datad(WideOr141),
	.cin(gnd),
	.combout(WideOr142),
	.cout());
// synopsys translate_off
defparam WideOr14.lut_mask = 16'hCFFF;
defparam WideOr14.sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y33_N4
cycloneive_lcell_comb WideOr15(
// Equation(s):
// WideOr151 = (Equal26) # (((WideNor1 & WideNor11)) # (!\WideOr15~0_combout ))

	.dataa(Equal26),
	.datab(WideNor1),
	.datac(WideNor11),
	.datad(\WideOr15~0_combout ),
	.cin(gnd),
	.combout(WideOr151),
	.cout());
// synopsys translate_off
defparam WideOr15.lut_mask = 16'hEAFF;
defparam WideOr15.sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y33_N12
cycloneive_lcell_comb \WideOr16~0 (
// Equation(s):
// WideOr161 = (!Equal20 & WideNor1)

	.dataa(gnd),
	.datab(gnd),
	.datac(Equal20),
	.datad(WideNor1),
	.cin(gnd),
	.combout(WideOr161),
	.cout());
// synopsys translate_off
defparam \WideOr16~0 .lut_mask = 16'h0F00;
defparam \WideOr16~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y33_N14
cycloneive_lcell_comb \Selector14~0 (
// Equation(s):
// Selector14 = (\WideOr16~combout  & ((plif_ifidinstr_l_4) # ((plif_ifidinstr_l_10 & Selector0)))) # (!\WideOr16~combout  & (plif_ifidinstr_l_10 & (Selector0)))

	.dataa(\WideOr16~combout ),
	.datab(plif_ifidinstr_l_10),
	.datac(Selector0),
	.datad(plif_ifidinstr_l_4),
	.cin(gnd),
	.combout(Selector14),
	.cout());
// synopsys translate_off
defparam \Selector14~0 .lut_mask = 16'hEAC0;
defparam \Selector14~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y33_N0
cycloneive_lcell_comb \Selector15~0 (
// Equation(s):
// Selector15 = (plif_ifidinstr_l_3 & ((\WideOr16~combout ) # ((plif_ifidinstr_l_9 & Selector0)))) # (!plif_ifidinstr_l_3 & (plif_ifidinstr_l_9 & (Selector0)))

	.dataa(plif_ifidinstr_l_3),
	.datab(plif_ifidinstr_l_9),
	.datac(Selector0),
	.datad(\WideOr16~combout ),
	.cin(gnd),
	.combout(Selector15),
	.cout());
// synopsys translate_off
defparam \Selector15~0 .lut_mask = 16'hEAC0;
defparam \Selector15~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y33_N6
cycloneive_lcell_comb \Selector16~0 (
// Equation(s):
// Selector16 = (Selector0 & ((plif_ifidinstr_l_8) # ((plif_ifidinstr_l_2 & \WideOr16~combout )))) # (!Selector0 & (plif_ifidinstr_l_2 & ((\WideOr16~combout ))))

	.dataa(Selector0),
	.datab(plif_ifidinstr_l_2),
	.datac(plif_ifidinstr_l_8),
	.datad(\WideOr16~combout ),
	.cin(gnd),
	.combout(Selector16),
	.cout());
// synopsys translate_off
defparam \Selector16~0 .lut_mask = 16'hECA0;
defparam \Selector16~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y32_N0
cycloneive_lcell_comb \Selector17~0 (
// Equation(s):
// Selector17 = (plif_ifidinstr_l_7 & ((Selector0) # ((plif_ifidinstr_l_1 & \WideOr16~combout )))) # (!plif_ifidinstr_l_7 & (plif_ifidinstr_l_1 & (\WideOr16~combout )))

	.dataa(plif_ifidinstr_l_7),
	.datab(plif_ifidinstr_l_1),
	.datac(\WideOr16~combout ),
	.datad(Selector0),
	.cin(gnd),
	.combout(Selector17),
	.cout());
// synopsys translate_off
defparam \Selector17~0 .lut_mask = 16'hEAC0;
defparam \Selector17~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y33_N20
cycloneive_lcell_comb \Selector18~0 (
// Equation(s):
// Selector18 = (plif_ifidinstr_l_6 & ((Selector0) # ((plif_ifidinstr_l_0 & \WideOr16~combout )))) # (!plif_ifidinstr_l_6 & (plif_ifidinstr_l_0 & ((\WideOr16~combout ))))

	.dataa(plif_ifidinstr_l_6),
	.datab(plif_ifidinstr_l_0),
	.datac(Selector0),
	.datad(\WideOr16~combout ),
	.cin(gnd),
	.combout(Selector18),
	.cout());
// synopsys translate_off
defparam \Selector18~0 .lut_mask = 16'hECA0;
defparam \Selector18~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y30_N2
cycloneive_lcell_comb \Selector24~0 (
// Equation(s):
// Selector24 = (!plif_ifidinstr_l_30 & ((plif_ifidinstr_l_31 & (Equal16 & !plif_ifidinstr_l_29)) # (!plif_ifidinstr_l_31 & ((plif_ifidinstr_l_29)))))

	.dataa(plif_ifidinstr_l_31),
	.datab(Equal16),
	.datac(plif_ifidinstr_l_30),
	.datad(plif_ifidinstr_l_29),
	.cin(gnd),
	.combout(Selector24),
	.cout());
// synopsys translate_off
defparam \Selector24~0 .lut_mask = 16'h0508;
defparam \Selector24~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y30_N6
cycloneive_lcell_comb \Equal12~0 (
// Equation(s):
// Equal121 = (plif_ifidinstr_l_28 & (plif_ifidinstr_l_26 & !plif_ifidinstr_l_27))

	.dataa(plif_ifidinstr_l_28),
	.datab(gnd),
	.datac(plif_ifidinstr_l_26),
	.datad(plif_ifidinstr_l_27),
	.cin(gnd),
	.combout(Equal121),
	.cout());
// synopsys translate_off
defparam \Equal12~0 .lut_mask = 16'h00A0;
defparam \Equal12~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y33_N30
cycloneive_lcell_comb \Selector0~2 (
// Equation(s):
// Selector0 = (Equal26 & (!plif_ifidinstr_l_3 & Equal6))

	.dataa(Equal26),
	.datab(gnd),
	.datac(plif_ifidinstr_l_3),
	.datad(Equal6),
	.cin(gnd),
	.combout(Selector0),
	.cout());
// synopsys translate_off
defparam \Selector0~2 .lut_mask = 16'h0A00;
defparam \Selector0~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y29_N26
cycloneive_lcell_comb \Equal25~4 (
// Equation(s):
// Equal25 = (!plif_ifidinstr_l_28 & (plif_ifidinstr_l_26 & (Equal11 & plif_ifidinstr_l_27)))

	.dataa(plif_ifidinstr_l_28),
	.datab(plif_ifidinstr_l_26),
	.datac(Equal11),
	.datad(plif_ifidinstr_l_27),
	.cin(gnd),
	.combout(Equal25),
	.cout());
// synopsys translate_off
defparam \Equal25~4 .lut_mask = 16'h4000;
defparam \Equal25~4 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y30_N20
cycloneive_lcell_comb \Equal13~0 (
// Equation(s):
// \Equal13~0_combout  = (!plif_ifidinstr_l_30 & (plif_ifidinstr_l_29 & (!plif_ifidinstr_l_28 & !plif_ifidinstr_l_31)))

	.dataa(plif_ifidinstr_l_30),
	.datab(plif_ifidinstr_l_29),
	.datac(plif_ifidinstr_l_28),
	.datad(plif_ifidinstr_l_31),
	.cin(gnd),
	.combout(\Equal13~0_combout ),
	.cout());
// synopsys translate_off
defparam \Equal13~0 .lut_mask = 16'h0004;
defparam \Equal13~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y30_N4
cycloneive_lcell_comb \WideNor0~1 (
// Equation(s):
// \WideNor0~1_combout  = (!plif_ifidinstr_l_2 & (!plif_ifidinstr_l_5 & !plif_ifidinstr_l_0))

	.dataa(gnd),
	.datab(plif_ifidinstr_l_2),
	.datac(plif_ifidinstr_l_5),
	.datad(plif_ifidinstr_l_0),
	.cin(gnd),
	.combout(\WideNor0~1_combout ),
	.cout());
// synopsys translate_off
defparam \WideNor0~1 .lut_mask = 16'h0003;
defparam \WideNor0~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y30_N18
cycloneive_lcell_comb \WideNor0~0 (
// Equation(s):
// \WideNor0~0_combout  = (plif_ifidinstr_l_2 & (((!plif_ifidinstr_l_3)))) # (!plif_ifidinstr_l_2 & ((plif_ifidinstr_l_3 & ((plif_ifidinstr_l_1))) # (!plif_ifidinstr_l_3 & (plif_ifidinstr_l_0))))

	.dataa(plif_ifidinstr_l_0),
	.datab(plif_ifidinstr_l_2),
	.datac(plif_ifidinstr_l_3),
	.datad(plif_ifidinstr_l_1),
	.cin(gnd),
	.combout(\WideNor0~0_combout ),
	.cout());
// synopsys translate_off
defparam \WideNor0~0 .lut_mask = 16'h3E0E;
defparam \WideNor0~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y30_N16
cycloneive_lcell_comb \WideNor0~3 (
// Equation(s):
// \WideNor0~3_combout  = (plif_ifidinstr_l_5 & ((\WideNor0~0_combout ) # ((!WideNor0 & \WideNor0~1_combout )))) # (!plif_ifidinstr_l_5 & (!WideNor0 & (\WideNor0~1_combout )))

	.dataa(plif_ifidinstr_l_5),
	.datab(WideNor0),
	.datac(\WideNor0~1_combout ),
	.datad(\WideNor0~0_combout ),
	.cin(gnd),
	.combout(\WideNor0~3_combout ),
	.cout());
// synopsys translate_off
defparam \WideNor0~3 .lut_mask = 16'hBA30;
defparam \WideNor0~3 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y30_N8
cycloneive_lcell_comb \Selector5~0 (
// Equation(s):
// \Selector5~0_combout  = (!plif_ifidinstr_l_4 & (Equal26 & \WideNor0~3_combout ))

	.dataa(plif_ifidinstr_l_4),
	.datab(gnd),
	.datac(Equal26),
	.datad(\WideNor0~3_combout ),
	.cin(gnd),
	.combout(\Selector5~0_combout ),
	.cout());
// synopsys translate_off
defparam \Selector5~0 .lut_mask = 16'h5000;
defparam \Selector5~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y29_N6
cycloneive_lcell_comb \WideOr15~0 (
// Equation(s):
// \WideOr15~0_combout  = (pcsrc & (((!plif_ifidinstr_l_29) # (!plif_ifidinstr_l_30)) # (!Equal23)))

	.dataa(Equal23),
	.datab(pcsrc),
	.datac(plif_ifidinstr_l_30),
	.datad(plif_ifidinstr_l_29),
	.cin(gnd),
	.combout(\WideOr15~0_combout ),
	.cout());
// synopsys translate_off
defparam \WideOr15~0 .lut_mask = 16'h4CCC;
defparam \WideOr15~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y29_N0
cycloneive_lcell_comb \Selector22~3 (
// Equation(s):
// \Selector22~3_combout  = (plif_ifidinstr_l_5 & (plif_ifidinstr_l_0 & ((!plif_ifidinstr_l_3) # (!plif_ifidinstr_l_2)))) # (!plif_ifidinstr_l_5 & (!plif_ifidinstr_l_2 & (!plif_ifidinstr_l_0 & !plif_ifidinstr_l_3)))

	.dataa(plif_ifidinstr_l_5),
	.datab(plif_ifidinstr_l_2),
	.datac(plif_ifidinstr_l_0),
	.datad(plif_ifidinstr_l_3),
	.cin(gnd),
	.combout(\Selector22~3_combout ),
	.cout());
// synopsys translate_off
defparam \Selector22~3 .lut_mask = 16'h20A1;
defparam \Selector22~3 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y30_N6
cycloneive_lcell_comb \Selector22~8 (
// Equation(s):
// \Selector22~8_combout  = (plif_ifidinstr_l_1 & (!plif_ifidinstr_l_4 & \Selector22~3_combout ))

	.dataa(gnd),
	.datab(plif_ifidinstr_l_1),
	.datac(plif_ifidinstr_l_4),
	.datad(\Selector22~3_combout ),
	.cin(gnd),
	.combout(\Selector22~8_combout ),
	.cout());
// synopsys translate_off
defparam \Selector22~8 .lut_mask = 16'h0C00;
defparam \Selector22~8 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y30_N14
cycloneive_lcell_comb WideOr16(
// Equation(s):
// \WideOr16~combout  = (((Equal22) # (Equal20)) # (!Selector22)) # (!WideNor1)

	.dataa(WideNor1),
	.datab(Selector22),
	.datac(Equal22),
	.datad(Equal20),
	.cin(gnd),
	.combout(\WideOr16~combout ),
	.cout());
// synopsys translate_off
defparam WideOr16.lut_mask = 16'hFFF7;
defparam WideOr16.sum_lutc_input = "datac";
// synopsys translate_on

endmodule

module forwarding_unit (
	plif_exmemregen_l,
	plif_exmemwsel_l_0,
	plif_exmemwsel_l_1,
	plif_idexrsel2_l_1,
	plif_idexrsel2_l_0,
	plif_exmemwsel_l_4,
	plif_exmemwsel_l_3,
	plif_exmemwsel_l_2,
	always0,
	plif_idexrsel2_l_2,
	plif_idexrsel2_l_3,
	always01,
	plif_idexrsel2_l_4,
	always02,
	plif_memwbwsel_l_4,
	plif_memwbwsel_l_3,
	plif_memwbwsel_l_0,
	plif_memwbwsel_l_2,
	plif_memwbwsel_l_1,
	Decoder0,
	WideOr01,
	fwdc,
	plif_memwbregen_l,
	plif_idexrsel1_l_4,
	plif_idexrsel1_l_1,
	plif_idexrsel1_l_0,
	plif_idexrsel1_l_2,
	plif_idexrsel1_l_3,
	fwda,
	always03,
	devpor,
	devclrn,
	devoe);
input 	plif_exmemregen_l;
input 	plif_exmemwsel_l_0;
input 	plif_exmemwsel_l_1;
input 	plif_idexrsel2_l_1;
input 	plif_idexrsel2_l_0;
input 	plif_exmemwsel_l_4;
input 	plif_exmemwsel_l_3;
input 	plif_exmemwsel_l_2;
output 	always0;
input 	plif_idexrsel2_l_2;
input 	plif_idexrsel2_l_3;
output 	always01;
input 	plif_idexrsel2_l_4;
output 	always02;
input 	plif_memwbwsel_l_4;
input 	plif_memwbwsel_l_3;
input 	plif_memwbwsel_l_0;
input 	plif_memwbwsel_l_2;
input 	plif_memwbwsel_l_1;
input 	Decoder0;
output 	WideOr01;
output 	fwdc;
input 	plif_memwbregen_l;
input 	plif_idexrsel1_l_4;
input 	plif_idexrsel1_l_1;
input 	plif_idexrsel1_l_0;
input 	plif_idexrsel1_l_2;
input 	plif_idexrsel1_l_3;
output 	fwda;
output 	always03;

// Design Ports Information

input 	devpor;
input 	devclrn;
input 	devoe;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
assign unknown = 1'bx;

wire \always0~1_combout ;
wire \always0~0_combout ;
wire \fwdc~1_combout ;
wire \fwdc~0_combout ;
wire \Equal5~0_combout ;
wire \fwda~2_combout ;
wire \fwda~0_combout ;
wire \fwda~1_combout ;
wire \always0~7_combout ;
wire \always0~5_combout ;
wire \always0~6_combout ;


// Location: LCCOMB_X57_Y37_N14
cycloneive_lcell_comb \always0~2 (
// Equation(s):
// always0 = (plif_exmemregen_l & (\always0~0_combout  & ((plif_exmemwsel_l_0) # (\always0~1_combout ))))

	.dataa(plif_exmemwsel_l_0),
	.datab(\always0~1_combout ),
	.datac(plif_exmemregen_l),
	.datad(\always0~0_combout ),
	.cin(gnd),
	.combout(always0),
	.cout());
// synopsys translate_off
defparam \always0~2 .lut_mask = 16'hE000;
defparam \always0~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y37_N22
cycloneive_lcell_comb \always0~3 (
// Equation(s):
// always01 = (plif_exmemwsel_l_2 & (plif_idexrsel2_l_2 & (plif_exmemwsel_l_3 $ (!plif_idexrsel2_l_3)))) # (!plif_exmemwsel_l_2 & (!plif_idexrsel2_l_2 & (plif_exmemwsel_l_3 $ (!plif_idexrsel2_l_3))))

	.dataa(plif_exmemwsel_l_2),
	.datab(plif_idexrsel2_l_2),
	.datac(plif_exmemwsel_l_3),
	.datad(plif_idexrsel2_l_3),
	.cin(gnd),
	.combout(always01),
	.cout());
// synopsys translate_off
defparam \always0~3 .lut_mask = 16'h9009;
defparam \always0~3 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y37_N30
cycloneive_lcell_comb \always0~4 (
// Equation(s):
// always02 = (always01 & (always0 & (plif_idexrsel2_l_4 $ (!plif_exmemwsel_l_4))))

	.dataa(always01),
	.datab(plif_idexrsel2_l_4),
	.datac(plif_exmemwsel_l_4),
	.datad(always0),
	.cin(gnd),
	.combout(always02),
	.cout());
// synopsys translate_off
defparam \always0~4 .lut_mask = 16'h8200;
defparam \always0~4 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y37_N28
cycloneive_lcell_comb WideOr0(
// Equation(s):
// WideOr01 = (plif_memwbwsel_l_0) # ((plif_memwbwsel_l_3) # ((plif_memwbwsel_l_4) # (!Decoder0)))

	.dataa(plif_memwbwsel_l_0),
	.datab(plif_memwbwsel_l_3),
	.datac(plif_memwbwsel_l_4),
	.datad(Decoder0),
	.cin(gnd),
	.combout(WideOr01),
	.cout());
// synopsys translate_off
defparam WideOr0.lut_mask = 16'hFEFF;
defparam WideOr0.sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y37_N12
cycloneive_lcell_comb \fwdc~2 (
// Equation(s):
// fwdc = (\fwdc~1_combout  & (\fwdc~0_combout  & (!\Equal5~0_combout  & WideOr01)))

	.dataa(\fwdc~1_combout ),
	.datab(\fwdc~0_combout ),
	.datac(\Equal5~0_combout ),
	.datad(WideOr01),
	.cin(gnd),
	.combout(fwdc),
	.cout());
// synopsys translate_off
defparam \fwdc~2 .lut_mask = 16'h0800;
defparam \fwdc~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y37_N28
cycloneive_lcell_comb \fwda~3 (
// Equation(s):
// fwda = (\fwda~2_combout  & (\fwda~0_combout  & (\fwda~1_combout  & WideOr01)))

	.dataa(\fwda~2_combout ),
	.datab(\fwda~0_combout ),
	.datac(\fwda~1_combout ),
	.datad(WideOr01),
	.cin(gnd),
	.combout(fwda),
	.cout());
// synopsys translate_off
defparam \fwda~3 .lut_mask = 16'h8000;
defparam \fwda~3 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y37_N0
cycloneive_lcell_comb \always0~8 (
// Equation(s):
// always03 = (\always0~7_combout  & (\always0~6_combout  & (plif_idexrsel1_l_4 $ (!plif_exmemwsel_l_4))))

	.dataa(plif_idexrsel1_l_4),
	.datab(plif_exmemwsel_l_4),
	.datac(\always0~7_combout ),
	.datad(\always0~6_combout ),
	.cin(gnd),
	.combout(always03),
	.cout());
// synopsys translate_off
defparam \always0~8 .lut_mask = 16'h9000;
defparam \always0~8 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y37_N0
cycloneive_lcell_comb \always0~1 (
// Equation(s):
// \always0~1_combout  = (plif_exmemwsel_l_1) # ((plif_exmemwsel_l_3) # ((plif_exmemwsel_l_2) # (plif_exmemwsel_l_4)))

	.dataa(plif_exmemwsel_l_1),
	.datab(plif_exmemwsel_l_3),
	.datac(plif_exmemwsel_l_2),
	.datad(plif_exmemwsel_l_4),
	.cin(gnd),
	.combout(\always0~1_combout ),
	.cout());
// synopsys translate_off
defparam \always0~1 .lut_mask = 16'hFFFE;
defparam \always0~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y37_N26
cycloneive_lcell_comb \always0~0 (
// Equation(s):
// \always0~0_combout  = (plif_exmemwsel_l_1 & (plif_idexrsel2_l_1 & (plif_exmemwsel_l_0 $ (!plif_idexrsel2_l_0)))) # (!plif_exmemwsel_l_1 & (!plif_idexrsel2_l_1 & (plif_exmemwsel_l_0 $ (!plif_idexrsel2_l_0))))

	.dataa(plif_exmemwsel_l_1),
	.datab(plif_idexrsel2_l_1),
	.datac(plif_exmemwsel_l_0),
	.datad(plif_idexrsel2_l_0),
	.cin(gnd),
	.combout(\always0~0_combout ),
	.cout());
// synopsys translate_off
defparam \always0~0 .lut_mask = 16'h9009;
defparam \always0~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y37_N20
cycloneive_lcell_comb \fwdc~1 (
// Equation(s):
// \fwdc~1_combout  = (plif_memwbwsel_l_2 & (plif_idexrsel2_l_2 & (plif_memwbwsel_l_3 $ (!plif_idexrsel2_l_3)))) # (!plif_memwbwsel_l_2 & (!plif_idexrsel2_l_2 & (plif_memwbwsel_l_3 $ (!plif_idexrsel2_l_3))))

	.dataa(plif_memwbwsel_l_2),
	.datab(plif_idexrsel2_l_2),
	.datac(plif_memwbwsel_l_3),
	.datad(plif_idexrsel2_l_3),
	.cin(gnd),
	.combout(\fwdc~1_combout ),
	.cout());
// synopsys translate_off
defparam \fwdc~1 .lut_mask = 16'h9009;
defparam \fwdc~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y37_N8
cycloneive_lcell_comb \fwdc~0 (
// Equation(s):
// \fwdc~0_combout  = (plif_idexrsel2_l_0 & (plif_memwbwsel_l_0 & (plif_memwbwsel_l_1 $ (!plif_idexrsel2_l_1)))) # (!plif_idexrsel2_l_0 & (!plif_memwbwsel_l_0 & (plif_memwbwsel_l_1 $ (!plif_idexrsel2_l_1))))

	.dataa(plif_idexrsel2_l_0),
	.datab(plif_memwbwsel_l_1),
	.datac(plif_memwbwsel_l_0),
	.datad(plif_idexrsel2_l_1),
	.cin(gnd),
	.combout(\fwdc~0_combout ),
	.cout());
// synopsys translate_off
defparam \fwdc~0 .lut_mask = 16'h8421;
defparam \fwdc~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y37_N4
cycloneive_lcell_comb \Equal5~0 (
// Equation(s):
// \Equal5~0_combout  = plif_idexrsel2_l_4 $ (plif_memwbwsel_l_4)

	.dataa(gnd),
	.datab(plif_idexrsel2_l_4),
	.datac(gnd),
	.datad(plif_memwbwsel_l_4),
	.cin(gnd),
	.combout(\Equal5~0_combout ),
	.cout());
// synopsys translate_off
defparam \Equal5~0 .lut_mask = 16'h33CC;
defparam \Equal5~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y37_N10
cycloneive_lcell_comb \fwda~2 (
// Equation(s):
// \fwda~2_combout  = (plif_memwbwsel_l_3 & (plif_idexrsel1_l_3 & (plif_idexrsel1_l_2 $ (!plif_memwbwsel_l_2)))) # (!plif_memwbwsel_l_3 & (!plif_idexrsel1_l_3 & (plif_idexrsel1_l_2 $ (!plif_memwbwsel_l_2))))

	.dataa(plif_memwbwsel_l_3),
	.datab(plif_idexrsel1_l_2),
	.datac(plif_idexrsel1_l_3),
	.datad(plif_memwbwsel_l_2),
	.cin(gnd),
	.combout(\fwda~2_combout ),
	.cout());
// synopsys translate_off
defparam \fwda~2 .lut_mask = 16'h8421;
defparam \fwda~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y37_N2
cycloneive_lcell_comb \fwda~0 (
// Equation(s):
// \fwda~0_combout  = (plif_memwbregen_l & (plif_memwbwsel_l_4 $ (!plif_idexrsel1_l_4)))

	.dataa(plif_memwbregen_l),
	.datab(gnd),
	.datac(plif_memwbwsel_l_4),
	.datad(plif_idexrsel1_l_4),
	.cin(gnd),
	.combout(\fwda~0_combout ),
	.cout());
// synopsys translate_off
defparam \fwda~0 .lut_mask = 16'hA00A;
defparam \fwda~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y37_N4
cycloneive_lcell_comb \fwda~1 (
// Equation(s):
// \fwda~1_combout  = (plif_idexrsel1_l_0 & (plif_memwbwsel_l_0 & (plif_idexrsel1_l_1 $ (!plif_memwbwsel_l_1)))) # (!plif_idexrsel1_l_0 & (!plif_memwbwsel_l_0 & (plif_idexrsel1_l_1 $ (!plif_memwbwsel_l_1))))

	.dataa(plif_idexrsel1_l_0),
	.datab(plif_idexrsel1_l_1),
	.datac(plif_memwbwsel_l_0),
	.datad(plif_memwbwsel_l_1),
	.cin(gnd),
	.combout(\fwda~1_combout ),
	.cout());
// synopsys translate_off
defparam \fwda~1 .lut_mask = 16'h8421;
defparam \fwda~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y37_N14
cycloneive_lcell_comb \always0~7 (
// Equation(s):
// \always0~7_combout  = (plif_exmemwsel_l_3 & (plif_idexrsel1_l_3 & (plif_exmemwsel_l_2 $ (!plif_idexrsel1_l_2)))) # (!plif_exmemwsel_l_3 & (!plif_idexrsel1_l_3 & (plif_exmemwsel_l_2 $ (!plif_idexrsel1_l_2))))

	.dataa(plif_exmemwsel_l_3),
	.datab(plif_idexrsel1_l_3),
	.datac(plif_exmemwsel_l_2),
	.datad(plif_idexrsel1_l_2),
	.cin(gnd),
	.combout(\always0~7_combout ),
	.cout());
// synopsys translate_off
defparam \always0~7 .lut_mask = 16'h9009;
defparam \always0~7 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y37_N10
cycloneive_lcell_comb \always0~5 (
// Equation(s):
// \always0~5_combout  = (plif_exmemwsel_l_0 & (plif_idexrsel1_l_0 & (plif_exmemwsel_l_1 $ (!plif_idexrsel1_l_1)))) # (!plif_exmemwsel_l_0 & (!plif_idexrsel1_l_0 & (plif_exmemwsel_l_1 $ (!plif_idexrsel1_l_1))))

	.dataa(plif_exmemwsel_l_0),
	.datab(plif_idexrsel1_l_0),
	.datac(plif_exmemwsel_l_1),
	.datad(plif_idexrsel1_l_1),
	.cin(gnd),
	.combout(\always0~5_combout ),
	.cout());
// synopsys translate_off
defparam \always0~5 .lut_mask = 16'h9009;
defparam \always0~5 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y37_N16
cycloneive_lcell_comb \always0~6 (
// Equation(s):
// \always0~6_combout  = (plif_exmemregen_l & (\always0~5_combout  & ((plif_exmemwsel_l_0) # (\always0~1_combout ))))

	.dataa(plif_exmemwsel_l_0),
	.datab(\always0~1_combout ),
	.datac(plif_exmemregen_l),
	.datad(\always0~5_combout ),
	.cin(gnd),
	.combout(\always0~6_combout ),
	.cout());
// synopsys translate_off
defparam \always0~6 .lut_mask = 16'hE000;
defparam \always0~6 .sum_lutc_input = "datac";
// synopsys translate_on

endmodule

module hazard_unit (
	always1,
	plif_memwbpcsrc_l_1,
	plif_memwbpcsrc_l_0,
	always0,
	plif_idexpcsrc_l_1,
	plif_idexpcsrc_l_0,
	plif_exmempcsrc_l_1,
	plif_exmempcsrc_l_0,
	ifid_sRST,
	exmem_en,
	pcsrc,
	plif_idexdmemREN_l,
	plif_idexwsel_l_0,
	plif_idexwsel_l_1,
	Selector4,
	Selector5,
	plif_idexwsel_l_2,
	plif_idexwsel_l_3,
	Selector2,
	Selector3,
	plif_idexwsel_l_4,
	Selector1,
	Selector9,
	Selector10,
	Selector7,
	Selector8,
	Selector6,
	ifid_en,
	rambusy,
	idex_sRST,
	idex_sRST1,
	idex_sRST2,
	ifid_sRST1,
	devpor,
	devclrn,
	devoe);
input 	always1;
input 	plif_memwbpcsrc_l_1;
input 	plif_memwbpcsrc_l_0;
input 	always0;
input 	plif_idexpcsrc_l_1;
input 	plif_idexpcsrc_l_0;
input 	plif_exmempcsrc_l_1;
input 	plif_exmempcsrc_l_0;
output 	ifid_sRST;
output 	exmem_en;
input 	pcsrc;
input 	plif_idexdmemREN_l;
input 	plif_idexwsel_l_0;
input 	plif_idexwsel_l_1;
input 	Selector4;
input 	Selector5;
input 	plif_idexwsel_l_2;
input 	plif_idexwsel_l_3;
input 	Selector2;
input 	Selector3;
input 	plif_idexwsel_l_4;
input 	Selector1;
input 	Selector9;
input 	Selector10;
input 	Selector7;
input 	Selector8;
input 	Selector6;
output 	ifid_en;
output 	rambusy;
output 	idex_sRST;
output 	idex_sRST1;
output 	idex_sRST2;
output 	ifid_sRST1;

// Design Ports Information

input 	devpor;
input 	devclrn;
input 	devoe;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
assign unknown = 1'bx;

wire \Equal0~1_combout ;
wire \WideOr2~combout ;
wire \Equal0~0_combout ;
wire \Equal0~2_combout ;
wire \Equal1~1_combout ;
wire \Equal1~0_combout ;
wire \Equal1~2_combout ;
wire \idex_sRST~2_combout ;


// Location: LCCOMB_X60_Y32_N10
cycloneive_lcell_comb \Equal0~1 (
// Equation(s):
// \Equal0~1_combout  = (plif_idexwsel_l_2 & (Selector3 & (plif_idexwsel_l_3 $ (!Selector2)))) # (!plif_idexwsel_l_2 & (!Selector3 & (plif_idexwsel_l_3 $ (!Selector2))))

	.dataa(plif_idexwsel_l_2),
	.datab(plif_idexwsel_l_3),
	.datac(Selector3),
	.datad(Selector2),
	.cin(gnd),
	.combout(\Equal0~1_combout ),
	.cout());
// synopsys translate_off
defparam \Equal0~1 .lut_mask = 16'h8421;
defparam \Equal0~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y32_N18
cycloneive_lcell_comb \ifid_sRST~2 (
// Equation(s):
// ifid_sRST = (!plif_exmempcsrc_l_1 & (!plif_idexpcsrc_l_1 & (!plif_exmempcsrc_l_0 & !plif_idexpcsrc_l_0)))

	.dataa(plif_exmempcsrc_l_1),
	.datab(plif_idexpcsrc_l_1),
	.datac(plif_exmempcsrc_l_0),
	.datad(plif_idexpcsrc_l_0),
	.cin(gnd),
	.combout(ifid_sRST),
	.cout());
// synopsys translate_off
defparam \ifid_sRST~2 .lut_mask = 16'h0001;
defparam \ifid_sRST~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y32_N20
cycloneive_lcell_comb \exmem_en~0 (
// Equation(s):
// exmem_en = ((always1) # ((\WideOr2~combout ) # (!ifid_sRST))) # (!always0)

	.dataa(always0),
	.datab(always1),
	.datac(ifid_sRST),
	.datad(\WideOr2~combout ),
	.cin(gnd),
	.combout(exmem_en),
	.cout());
// synopsys translate_off
defparam \exmem_en~0 .lut_mask = 16'hFFDF;
defparam \exmem_en~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y33_N12
cycloneive_lcell_comb \ifid_en~0 (
// Equation(s):
// ifid_en = (ifid_sRST & ((\WideOr2~combout ) # ((!\idex_sRST~2_combout  & !always0))))

	.dataa(\WideOr2~combout ),
	.datab(ifid_sRST),
	.datac(\idex_sRST~2_combout ),
	.datad(always0),
	.cin(gnd),
	.combout(ifid_en),
	.cout());
// synopsys translate_off
defparam \ifid_en~0 .lut_mask = 16'h888C;
defparam \ifid_en~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y32_N10
cycloneive_lcell_comb \rambusy~0 (
// Equation(s):
// rambusy = (!always0 & (ifid_sRST & ((\WideOr2~combout ) # (!\idex_sRST~2_combout ))))

	.dataa(always0),
	.datab(ifid_sRST),
	.datac(\idex_sRST~2_combout ),
	.datad(\WideOr2~combout ),
	.cin(gnd),
	.combout(rambusy),
	.cout());
// synopsys translate_off
defparam \rambusy~0 .lut_mask = 16'h4404;
defparam \rambusy~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y32_N26
cycloneive_lcell_comb \idex_sRST~3 (
// Equation(s):
// idex_sRST = (!\WideOr2~combout  & ((always0 & (always1)) # (!always0 & ((\idex_sRST~2_combout )))))

	.dataa(always0),
	.datab(always1),
	.datac(\idex_sRST~2_combout ),
	.datad(\WideOr2~combout ),
	.cin(gnd),
	.combout(idex_sRST),
	.cout());
// synopsys translate_off
defparam \idex_sRST~3 .lut_mask = 16'h00D8;
defparam \idex_sRST~3 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y32_N24
cycloneive_lcell_comb \idex_sRST~4 (
// Equation(s):
// idex_sRST1 = (idex_sRST) # (idex_sRST2)

	.dataa(idex_sRST),
	.datab(idex_sRST2),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(idex_sRST1),
	.cout());
// synopsys translate_off
defparam \idex_sRST~4 .lut_mask = 16'hEEEE;
defparam \idex_sRST~4 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y32_N14
cycloneive_lcell_comb \idex_sRST~5 (
// Equation(s):
// idex_sRST2 = (plif_memwbpcsrc_l_1) # (((plif_memwbpcsrc_l_0 & \pcsrc~0_combout )) # (!ifid_sRST))

	.dataa(plif_memwbpcsrc_l_0),
	.datab(pcsrc),
	.datac(plif_memwbpcsrc_l_1),
	.datad(ifid_sRST),
	.cin(gnd),
	.combout(idex_sRST2),
	.cout());
// synopsys translate_off
defparam \idex_sRST~5 .lut_mask = 16'hF8FF;
defparam \idex_sRST~5 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y32_N0
cycloneive_lcell_comb \ifid_sRST~3 (
// Equation(s):
// ifid_sRST1 = (ifid_sRST & ((plif_memwbpcsrc_l_1) # ((plif_memwbpcsrc_l_0 & \pcsrc~0_combout ))))

	.dataa(plif_memwbpcsrc_l_0),
	.datab(pcsrc),
	.datac(plif_memwbpcsrc_l_1),
	.datad(ifid_sRST),
	.cin(gnd),
	.combout(ifid_sRST1),
	.cout());
// synopsys translate_off
defparam \ifid_sRST~3 .lut_mask = 16'hF800;
defparam \ifid_sRST~3 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y32_N2
cycloneive_lcell_comb WideOr2(
// Equation(s):
// \WideOr2~combout  = (plif_memwbpcsrc_l_1) # (plif_memwbpcsrc_l_0)

	.dataa(gnd),
	.datab(plif_memwbpcsrc_l_1),
	.datac(gnd),
	.datad(plif_memwbpcsrc_l_0),
	.cin(gnd),
	.combout(\WideOr2~combout ),
	.cout());
// synopsys translate_off
defparam WideOr2.lut_mask = 16'hFFCC;
defparam WideOr2.sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y32_N12
cycloneive_lcell_comb \Equal0~0 (
// Equation(s):
// \Equal0~0_combout  = (plif_idexwsel_l_1 & (Selector41 & (plif_idexwsel_l_0 $ (!Selector5)))) # (!plif_idexwsel_l_1 & (!Selector41 & (plif_idexwsel_l_0 $ (!Selector5))))

	.dataa(plif_idexwsel_l_1),
	.datab(plif_idexwsel_l_0),
	.datac(Selector5),
	.datad(Selector4),
	.cin(gnd),
	.combout(\Equal0~0_combout ),
	.cout());
// synopsys translate_off
defparam \Equal0~0 .lut_mask = 16'h8241;
defparam \Equal0~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y32_N14
cycloneive_lcell_comb \Equal0~2 (
// Equation(s):
// \Equal0~2_combout  = (\Equal0~1_combout  & (\Equal0~0_combout  & (Selector1 $ (!plif_idexwsel_l_4))))

	.dataa(\Equal0~1_combout ),
	.datab(Selector1),
	.datac(plif_idexwsel_l_4),
	.datad(\Equal0~0_combout ),
	.cin(gnd),
	.combout(\Equal0~2_combout ),
	.cout());
// synopsys translate_off
defparam \Equal0~2 .lut_mask = 16'h8200;
defparam \Equal0~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y32_N30
cycloneive_lcell_comb \Equal1~1 (
// Equation(s):
// \Equal1~1_combout  = (plif_idexwsel_l_3 & (Selector7 & (Selector8 $ (!plif_idexwsel_l_2)))) # (!plif_idexwsel_l_3 & (!Selector7 & (Selector8 $ (!plif_idexwsel_l_2))))

	.dataa(plif_idexwsel_l_3),
	.datab(Selector8),
	.datac(plif_idexwsel_l_2),
	.datad(Selector7),
	.cin(gnd),
	.combout(\Equal1~1_combout ),
	.cout());
// synopsys translate_off
defparam \Equal1~1 .lut_mask = 16'h8241;
defparam \Equal1~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y32_N16
cycloneive_lcell_comb \Equal1~0 (
// Equation(s):
// \Equal1~0_combout  = (plif_idexwsel_l_1 & (Selector91 & (plif_idexwsel_l_0 $ (!Selector10)))) # (!plif_idexwsel_l_1 & (!Selector91 & (plif_idexwsel_l_0 $ (!Selector10))))

	.dataa(plif_idexwsel_l_1),
	.datab(plif_idexwsel_l_0),
	.datac(Selector10),
	.datad(Selector9),
	.cin(gnd),
	.combout(\Equal1~0_combout ),
	.cout());
// synopsys translate_off
defparam \Equal1~0 .lut_mask = 16'h8241;
defparam \Equal1~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y32_N28
cycloneive_lcell_comb \Equal1~2 (
// Equation(s):
// \Equal1~2_combout  = (\Equal1~1_combout  & (\Equal1~0_combout  & (Selector6 $ (!plif_idexwsel_l_4))))

	.dataa(Selector6),
	.datab(plif_idexwsel_l_4),
	.datac(\Equal1~1_combout ),
	.datad(\Equal1~0_combout ),
	.cin(gnd),
	.combout(\Equal1~2_combout ),
	.cout());
// synopsys translate_off
defparam \Equal1~2 .lut_mask = 16'h9000;
defparam \Equal1~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y32_N6
cycloneive_lcell_comb \idex_sRST~2 (
// Equation(s):
// \idex_sRST~2_combout  = (plif_idexdmemREN_l & ((\Equal0~2_combout ) # (\Equal1~2_combout )))

	.dataa(gnd),
	.datab(plif_idexdmemREN_l),
	.datac(\Equal0~2_combout ),
	.datad(\Equal1~2_combout ),
	.cin(gnd),
	.combout(\idex_sRST~2_combout ),
	.cout());
// synopsys translate_off
defparam \idex_sRST~2 .lut_mask = 16'hCCC0;
defparam \idex_sRST~2 .sum_lutc_input = "datac";
// synopsys translate_on

endmodule

module pc (
	PCreg_1,
	PCreg_0,
	pcifrtnaddr_2,
	pcifrtnaddr_3,
	pcifrtnaddr_4,
	pcifrtnaddr_5,
	pcifrtnaddr_6,
	pcifrtnaddr_7,
	pcifrtnaddr_8,
	pcifrtnaddr_9,
	pcifrtnaddr_10,
	pcifrtnaddr_11,
	pcifrtnaddr_12,
	pcifrtnaddr_13,
	pcifrtnaddr_14,
	pcifrtnaddr_15,
	pcifrtnaddr_16,
	pcifrtnaddr_17,
	pcifrtnaddr_18,
	pcifrtnaddr_19,
	pcifrtnaddr_20,
	pcifrtnaddr_21,
	pcifrtnaddr_22,
	pcifrtnaddr_23,
	pcifrtnaddr_24,
	pcifrtnaddr_25,
	pcifrtnaddr_26,
	pcifrtnaddr_27,
	pcifrtnaddr_28,
	pcifrtnaddr_29,
	pcifrtnaddr_30,
	pcifrtnaddr_31,
	PCreg_3,
	PCreg_2,
	PCreg_5,
	PCreg_4,
	PCreg_7,
	PCreg_6,
	PCreg_9,
	PCreg_8,
	PCreg_11,
	PCreg_10,
	PCreg_13,
	PCreg_12,
	PCreg_15,
	PCreg_14,
	PCreg_17,
	PCreg_16,
	PCreg_19,
	PCreg_18,
	PCreg_21,
	PCreg_20,
	PCreg_23,
	PCreg_22,
	PCreg_25,
	PCreg_24,
	PCreg_27,
	PCreg_26,
	PCreg_29,
	PCreg_28,
	PCreg_31,
	PCreg_30,
	plif_memwbpcsrc_l_1,
	always0,
	plif_memwbporto_l_31,
	plif_memwbrtnaddr_l_31,
	plif_memwbporto_l_30,
	plif_memwbrtnaddr_l_30,
	plif_memwbporto_l_29,
	plif_memwbrtnaddr_l_29,
	plif_memwbporto_l_28,
	plif_memwbrtnaddr_l_28,
	plif_memwbporto_l_27,
	plif_memwbrtnaddr_l_27,
	plif_memwbporto_l_26,
	plif_memwbrtnaddr_l_26,
	plif_memwbporto_l_25,
	plif_memwbrtnaddr_l_25,
	plif_memwbporto_l_24,
	plif_memwbrtnaddr_l_24,
	plif_memwbporto_l_23,
	plif_memwbrtnaddr_l_23,
	plif_memwbporto_l_22,
	plif_memwbrtnaddr_l_22,
	plif_memwbporto_l_21,
	plif_memwbrtnaddr_l_21,
	plif_memwbporto_l_20,
	plif_memwbrtnaddr_l_20,
	plif_memwbporto_l_19,
	plif_memwbrtnaddr_l_19,
	plif_memwbporto_l_18,
	plif_memwbrtnaddr_l_18,
	plif_memwbporto_l_17,
	plif_memwbrtnaddr_l_17,
	plif_memwbporto_l_16,
	plif_memwbrtnaddr_l_16,
	plif_memwbporto_l_15,
	plif_memwbrtnaddr_l_15,
	plif_memwbporto_l_14,
	plif_memwbrtnaddr_l_14,
	plif_memwbporto_l_13,
	plif_memwbrtnaddr_l_13,
	plif_memwbporto_l_12,
	plif_memwbrtnaddr_l_12,
	plif_memwbporto_l_11,
	plif_memwbrtnaddr_l_11,
	plif_memwbporto_l_10,
	plif_memwbrtnaddr_l_10,
	plif_memwbporto_l_9,
	plif_memwbrtnaddr_l_9,
	plif_memwbporto_l_8,
	plif_memwbrtnaddr_l_8,
	plif_memwbporto_l_7,
	plif_memwbrtnaddr_l_7,
	plif_memwbporto_l_6,
	plif_memwbrtnaddr_l_6,
	plif_memwbporto_l_5,
	plif_memwbrtnaddr_l_5,
	plif_memwbporto_l_2,
	plif_memwbrtnaddr_l_2,
	plif_memwbporto_l_1,
	plif_memwbrtnaddr_l_1,
	plif_memwbporto_l_0,
	plif_memwbrtnaddr_l_0,
	plif_memwbporto_l_4,
	plif_memwbrtnaddr_l_4,
	plif_memwbporto_l_3,
	plif_memwbrtnaddr_l_3,
	pcsrc,
	ifid_en,
	plif_memwbjaddr_l_1,
	plif_memwbextimm_l_1,
	plif_memwbextimm_l_0,
	\pcif.rambusy ,
	plif_memwbjaddr_l_0,
	plif_memwbjaddr_l_3,
	plif_memwbextimm_l_3,
	plif_memwbextimm_l_2,
	plif_memwbjaddr_l_2,
	plif_memwbjaddr_l_5,
	plif_memwbextimm_l_5,
	plif_memwbextimm_l_4,
	plif_memwbjaddr_l_4,
	plif_memwbjaddr_l_7,
	plif_memwbextimm_l_7,
	plif_memwbextimm_l_6,
	plif_memwbjaddr_l_6,
	plif_memwbjaddr_l_9,
	plif_memwbextimm_l_9,
	plif_memwbextimm_l_8,
	plif_memwbjaddr_l_8,
	plif_memwbjaddr_l_11,
	plif_memwbextimm_l_11,
	plif_memwbextimm_l_10,
	plif_memwbjaddr_l_10,
	plif_memwbjaddr_l_13,
	plif_memwbextimm_l_13,
	plif_memwbextimm_l_12,
	plif_memwbjaddr_l_12,
	plif_memwbjaddr_l_15,
	plif_memwbextimm_l_15,
	plif_memwbextimm_l_14,
	plif_memwbjaddr_l_14,
	plif_memwbjaddr_l_17,
	plif_memwbextimm_l_17,
	plif_memwbextimm_l_16,
	plif_memwbjaddr_l_16,
	plif_memwbjaddr_l_19,
	plif_memwbextimm_l_19,
	plif_memwbextimm_l_18,
	plif_memwbjaddr_l_18,
	plif_memwbjaddr_l_21,
	plif_memwbextimm_l_21,
	plif_memwbextimm_l_20,
	plif_memwbjaddr_l_20,
	plif_memwbjaddr_l_23,
	plif_memwbextimm_l_23,
	plif_memwbextimm_l_22,
	plif_memwbjaddr_l_22,
	plif_memwbjaddr_l_25,
	plif_memwbextimm_l_25,
	plif_memwbextimm_l_24,
	plif_memwbjaddr_l_24,
	plif_memwbextimm_l_27,
	plif_memwbextimm_l_26,
	plif_memwbextimm_l_29,
	plif_memwbextimm_l_28,
	CLK,
	nRST,
	devpor,
	devclrn,
	devoe);
output 	PCreg_1;
output 	PCreg_0;
output 	pcifrtnaddr_2;
output 	pcifrtnaddr_3;
output 	pcifrtnaddr_4;
output 	pcifrtnaddr_5;
output 	pcifrtnaddr_6;
output 	pcifrtnaddr_7;
output 	pcifrtnaddr_8;
output 	pcifrtnaddr_9;
output 	pcifrtnaddr_10;
output 	pcifrtnaddr_11;
output 	pcifrtnaddr_12;
output 	pcifrtnaddr_13;
output 	pcifrtnaddr_14;
output 	pcifrtnaddr_15;
output 	pcifrtnaddr_16;
output 	pcifrtnaddr_17;
output 	pcifrtnaddr_18;
output 	pcifrtnaddr_19;
output 	pcifrtnaddr_20;
output 	pcifrtnaddr_21;
output 	pcifrtnaddr_22;
output 	pcifrtnaddr_23;
output 	pcifrtnaddr_24;
output 	pcifrtnaddr_25;
output 	pcifrtnaddr_26;
output 	pcifrtnaddr_27;
output 	pcifrtnaddr_28;
output 	pcifrtnaddr_29;
output 	pcifrtnaddr_30;
output 	pcifrtnaddr_31;
output 	PCreg_3;
output 	PCreg_2;
output 	PCreg_5;
output 	PCreg_4;
output 	PCreg_7;
output 	PCreg_6;
output 	PCreg_9;
output 	PCreg_8;
output 	PCreg_11;
output 	PCreg_10;
output 	PCreg_13;
output 	PCreg_12;
output 	PCreg_15;
output 	PCreg_14;
output 	PCreg_17;
output 	PCreg_16;
output 	PCreg_19;
output 	PCreg_18;
output 	PCreg_21;
output 	PCreg_20;
output 	PCreg_23;
output 	PCreg_22;
output 	PCreg_25;
output 	PCreg_24;
output 	PCreg_27;
output 	PCreg_26;
output 	PCreg_29;
output 	PCreg_28;
output 	PCreg_31;
output 	PCreg_30;
input 	plif_memwbpcsrc_l_1;
input 	always0;
input 	plif_memwbporto_l_31;
input 	plif_memwbrtnaddr_l_31;
input 	plif_memwbporto_l_30;
input 	plif_memwbrtnaddr_l_30;
input 	plif_memwbporto_l_29;
input 	plif_memwbrtnaddr_l_29;
input 	plif_memwbporto_l_28;
input 	plif_memwbrtnaddr_l_28;
input 	plif_memwbporto_l_27;
input 	plif_memwbrtnaddr_l_27;
input 	plif_memwbporto_l_26;
input 	plif_memwbrtnaddr_l_26;
input 	plif_memwbporto_l_25;
input 	plif_memwbrtnaddr_l_25;
input 	plif_memwbporto_l_24;
input 	plif_memwbrtnaddr_l_24;
input 	plif_memwbporto_l_23;
input 	plif_memwbrtnaddr_l_23;
input 	plif_memwbporto_l_22;
input 	plif_memwbrtnaddr_l_22;
input 	plif_memwbporto_l_21;
input 	plif_memwbrtnaddr_l_21;
input 	plif_memwbporto_l_20;
input 	plif_memwbrtnaddr_l_20;
input 	plif_memwbporto_l_19;
input 	plif_memwbrtnaddr_l_19;
input 	plif_memwbporto_l_18;
input 	plif_memwbrtnaddr_l_18;
input 	plif_memwbporto_l_17;
input 	plif_memwbrtnaddr_l_17;
input 	plif_memwbporto_l_16;
input 	plif_memwbrtnaddr_l_16;
input 	plif_memwbporto_l_15;
input 	plif_memwbrtnaddr_l_15;
input 	plif_memwbporto_l_14;
input 	plif_memwbrtnaddr_l_14;
input 	plif_memwbporto_l_13;
input 	plif_memwbrtnaddr_l_13;
input 	plif_memwbporto_l_12;
input 	plif_memwbrtnaddr_l_12;
input 	plif_memwbporto_l_11;
input 	plif_memwbrtnaddr_l_11;
input 	plif_memwbporto_l_10;
input 	plif_memwbrtnaddr_l_10;
input 	plif_memwbporto_l_9;
input 	plif_memwbrtnaddr_l_9;
input 	plif_memwbporto_l_8;
input 	plif_memwbrtnaddr_l_8;
input 	plif_memwbporto_l_7;
input 	plif_memwbrtnaddr_l_7;
input 	plif_memwbporto_l_6;
input 	plif_memwbrtnaddr_l_6;
input 	plif_memwbporto_l_5;
input 	plif_memwbrtnaddr_l_5;
input 	plif_memwbporto_l_2;
input 	plif_memwbrtnaddr_l_2;
input 	plif_memwbporto_l_1;
input 	plif_memwbrtnaddr_l_1;
input 	plif_memwbporto_l_0;
input 	plif_memwbrtnaddr_l_0;
input 	plif_memwbporto_l_4;
input 	plif_memwbrtnaddr_l_4;
input 	plif_memwbporto_l_3;
input 	plif_memwbrtnaddr_l_3;
input 	pcsrc;
input 	ifid_en;
input 	plif_memwbjaddr_l_1;
input 	plif_memwbextimm_l_1;
input 	plif_memwbextimm_l_0;
input 	\pcif.rambusy ;
input 	plif_memwbjaddr_l_0;
input 	plif_memwbjaddr_l_3;
input 	plif_memwbextimm_l_3;
input 	plif_memwbextimm_l_2;
input 	plif_memwbjaddr_l_2;
input 	plif_memwbjaddr_l_5;
input 	plif_memwbextimm_l_5;
input 	plif_memwbextimm_l_4;
input 	plif_memwbjaddr_l_4;
input 	plif_memwbjaddr_l_7;
input 	plif_memwbextimm_l_7;
input 	plif_memwbextimm_l_6;
input 	plif_memwbjaddr_l_6;
input 	plif_memwbjaddr_l_9;
input 	plif_memwbextimm_l_9;
input 	plif_memwbextimm_l_8;
input 	plif_memwbjaddr_l_8;
input 	plif_memwbjaddr_l_11;
input 	plif_memwbextimm_l_11;
input 	plif_memwbextimm_l_10;
input 	plif_memwbjaddr_l_10;
input 	plif_memwbjaddr_l_13;
input 	plif_memwbextimm_l_13;
input 	plif_memwbextimm_l_12;
input 	plif_memwbjaddr_l_12;
input 	plif_memwbjaddr_l_15;
input 	plif_memwbextimm_l_15;
input 	plif_memwbextimm_l_14;
input 	plif_memwbjaddr_l_14;
input 	plif_memwbjaddr_l_17;
input 	plif_memwbextimm_l_17;
input 	plif_memwbextimm_l_16;
input 	plif_memwbjaddr_l_16;
input 	plif_memwbjaddr_l_19;
input 	plif_memwbextimm_l_19;
input 	plif_memwbextimm_l_18;
input 	plif_memwbjaddr_l_18;
input 	plif_memwbjaddr_l_21;
input 	plif_memwbextimm_l_21;
input 	plif_memwbextimm_l_20;
input 	plif_memwbjaddr_l_20;
input 	plif_memwbjaddr_l_23;
input 	plif_memwbextimm_l_23;
input 	plif_memwbextimm_l_22;
input 	plif_memwbjaddr_l_22;
input 	plif_memwbjaddr_l_25;
input 	plif_memwbextimm_l_25;
input 	plif_memwbextimm_l_24;
input 	plif_memwbjaddr_l_24;
input 	plif_memwbextimm_l_27;
input 	plif_memwbextimm_l_26;
input 	plif_memwbextimm_l_29;
input 	plif_memwbextimm_l_28;
input 	CLK;
input 	nRST;

// Design Ports Information

input 	devpor;
input 	devclrn;
input 	devoe;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
assign unknown = 1'bx;

wire \Add1~14_combout ;
wire \Add1~24_combout ;
wire \Add1~54_combout ;
wire \pcif.rtnaddr[2]~1 ;
wire \pcif.rtnaddr[3]~3 ;
wire \pcif.rtnaddr[4]~5 ;
wire \pcif.rtnaddr[5]~7 ;
wire \pcif.rtnaddr[6]~9 ;
wire \pcif.rtnaddr[7]~11 ;
wire \pcif.rtnaddr[8]~13 ;
wire \pcif.rtnaddr[9]~15 ;
wire \pcif.rtnaddr[10]~17 ;
wire \pcif.rtnaddr[11]~19 ;
wire \pcif.rtnaddr[12]~21 ;
wire \pcif.rtnaddr[13]~23 ;
wire \pcif.rtnaddr[14]~25 ;
wire \pcif.rtnaddr[15]~27 ;
wire \pcif.rtnaddr[16]~29 ;
wire \pcif.rtnaddr[17]~31 ;
wire \pcif.rtnaddr[18]~33 ;
wire \pcif.rtnaddr[19]~35 ;
wire \pcif.rtnaddr[20]~37 ;
wire \pcif.rtnaddr[21]~39 ;
wire \pcif.rtnaddr[22]~41 ;
wire \pcif.rtnaddr[23]~43 ;
wire \pcif.rtnaddr[24]~45 ;
wire \pcif.rtnaddr[25]~47 ;
wire \pcif.rtnaddr[26]~49 ;
wire \pcif.rtnaddr[27]~51 ;
wire \pcif.rtnaddr[28]~53 ;
wire \pcif.rtnaddr[29]~55 ;
wire \pcif.rtnaddr[30]~57 ;
wire \PCregN~0_combout ;
wire \PCreg[1]~feeder_combout ;
wire \PCreg[1]~0_combout ;
wire \PCregN~1_combout ;
wire \PCreg[0]~feeder_combout ;
wire \Add1~1 ;
wire \Add1~2_combout ;
wire \PCregN~2_combout ;
wire \PCregN~3_combout ;
wire \PCregN~4_combout ;
wire \Add1~0_combout ;
wire \PCregN~5_combout ;
wire \Add1~3 ;
wire \Add1~5 ;
wire \Add1~6_combout ;
wire \PCregN~6_combout ;
wire \PCregN~7_combout ;
wire \Add1~4_combout ;
wire \PCregN~8_combout ;
wire \PCregN~9_combout ;
wire \Add1~7 ;
wire \Add1~9 ;
wire \Add1~10_combout ;
wire \PCregN~10_combout ;
wire \PCregN~11_combout ;
wire \Add1~8_combout ;
wire \PCregN~12_combout ;
wire \PCregN~13_combout ;
wire \PCregN~14_combout ;
wire \PCregN~15_combout ;
wire \PCregN~16_combout ;
wire \Add1~11 ;
wire \Add1~12_combout ;
wire \PCregN~17_combout ;
wire \Add1~13 ;
wire \Add1~15 ;
wire \Add1~17 ;
wire \Add1~18_combout ;
wire \PCregN~18_combout ;
wire \PCregN~19_combout ;
wire \Add1~16_combout ;
wire \PCregN~20_combout ;
wire \PCregN~21_combout ;
wire \Add1~19 ;
wire \Add1~21 ;
wire \Add1~22_combout ;
wire \PCregN~22_combout ;
wire \PCregN~23_combout ;
wire \PCregN~24_combout ;
wire \Add1~20_combout ;
wire \PCregN~25_combout ;
wire \Add1~23 ;
wire \Add1~25 ;
wire \Add1~26_combout ;
wire \PCregN~26_combout ;
wire \PCregN~27_combout ;
wire \PCregN~28_combout ;
wire \PCregN~29_combout ;
wire \PCreg[14]~feeder_combout ;
wire \Add1~27 ;
wire \Add1~29 ;
wire \Add1~30_combout ;
wire \PCregN~30_combout ;
wire \PCregN~31_combout ;
wire \Add1~28_combout ;
wire \PCregN~32_combout ;
wire \PCregN~33_combout ;
wire \Add1~31 ;
wire \Add1~33 ;
wire \Add1~34_combout ;
wire \PCregN~34_combout ;
wire \PCregN~35_combout ;
wire \PCregN~36_combout ;
wire \Add1~32_combout ;
wire \PCregN~37_combout ;
wire \Add1~35 ;
wire \Add1~37 ;
wire \Add1~38_combout ;
wire \PCregN~38_combout ;
wire \PCregN~39_combout ;
wire \PCregN~40_combout ;
wire \Add1~36_combout ;
wire \PCregN~41_combout ;
wire \Add1~39 ;
wire \Add1~41 ;
wire \Add1~42_combout ;
wire \PCregN~42_combout ;
wire \PCregN~43_combout ;
wire \PCregN~44_combout ;
wire \Add1~40_combout ;
wire \PCregN~45_combout ;
wire \Add1~43 ;
wire \Add1~45 ;
wire \Add1~46_combout ;
wire \PCregN~46_combout ;
wire \PCregN~47_combout ;
wire \PCregN~48_combout ;
wire \Add1~44_combout ;
wire \PCregN~49_combout ;
wire \Add1~47 ;
wire \Add1~49 ;
wire \Add1~50_combout ;
wire \PCregN~50_combout ;
wire \PCregN~51_combout ;
wire \PCregN~52_combout ;
wire \Add1~48_combout ;
wire \PCregN~53_combout ;
wire \PCregN~54_combout ;
wire \PCregN~55_combout ;
wire \PCregN~56_combout ;
wire \Add1~51 ;
wire \Add1~52_combout ;
wire \PCregN~57_combout ;
wire \Add1~53 ;
wire \Add1~55 ;
wire \Add1~57 ;
wire \Add1~58_combout ;
wire \PCregN~58_combout ;
wire \PCregN~59_combout ;
wire \PCregN~60_combout ;
wire \Add1~56_combout ;
wire \PCregN~61_combout ;


// Location: LCCOMB_X56_Y32_N16
cycloneive_lcell_comb \Add1~14 (
// Equation(s):
// \Add1~14_combout  = (plif_memwbextimm_l_7 & ((plif_memwbrtnaddr_l_9 & (\Add1~13  & VCC)) # (!plif_memwbrtnaddr_l_9 & (!\Add1~13 )))) # (!plif_memwbextimm_l_7 & ((plif_memwbrtnaddr_l_9 & (!\Add1~13 )) # (!plif_memwbrtnaddr_l_9 & ((\Add1~13 ) # (GND)))))
// \Add1~15  = CARRY((plif_memwbextimm_l_7 & (!plif_memwbrtnaddr_l_9 & !\Add1~13 )) # (!plif_memwbextimm_l_7 & ((!\Add1~13 ) # (!plif_memwbrtnaddr_l_9))))

	.dataa(plif_memwbextimm_l_7),
	.datab(plif_memwbrtnaddr_l_9),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add1~13 ),
	.combout(\Add1~14_combout ),
	.cout(\Add1~15 ));
// synopsys translate_off
defparam \Add1~14 .lut_mask = 16'h9617;
defparam \Add1~14 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X56_Y32_N26
cycloneive_lcell_comb \Add1~24 (
// Equation(s):
// \Add1~24_combout  = ((plif_memwbextimm_l_12 $ (plif_memwbrtnaddr_l_14 $ (!\Add1~23 )))) # (GND)
// \Add1~25  = CARRY((plif_memwbextimm_l_12 & ((plif_memwbrtnaddr_l_14) # (!\Add1~23 ))) # (!plif_memwbextimm_l_12 & (plif_memwbrtnaddr_l_14 & !\Add1~23 )))

	.dataa(plif_memwbextimm_l_12),
	.datab(plif_memwbrtnaddr_l_14),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add1~23 ),
	.combout(\Add1~24_combout ),
	.cout(\Add1~25 ));
// synopsys translate_off
defparam \Add1~24 .lut_mask = 16'h698E;
defparam \Add1~24 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X56_Y31_N24
cycloneive_lcell_comb \Add1~54 (
// Equation(s):
// \Add1~54_combout  = (plif_memwbextimm_l_27 & ((plif_memwbrtnaddr_l_29 & (\Add1~53  & VCC)) # (!plif_memwbrtnaddr_l_29 & (!\Add1~53 )))) # (!plif_memwbextimm_l_27 & ((plif_memwbrtnaddr_l_29 & (!\Add1~53 )) # (!plif_memwbrtnaddr_l_29 & ((\Add1~53 ) # 
// (GND)))))
// \Add1~55  = CARRY((plif_memwbextimm_l_27 & (!plif_memwbrtnaddr_l_29 & !\Add1~53 )) # (!plif_memwbextimm_l_27 & ((!\Add1~53 ) # (!plif_memwbrtnaddr_l_29))))

	.dataa(plif_memwbextimm_l_27),
	.datab(plif_memwbrtnaddr_l_29),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add1~53 ),
	.combout(\Add1~54_combout ),
	.cout(\Add1~55 ));
// synopsys translate_off
defparam \Add1~54 .lut_mask = 16'h9617;
defparam \Add1~54 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: FF_X50_Y32_N25
dffeas \PCreg[1] (
	.clk(CLK),
	.d(\PCreg[1]~feeder_combout ),
	.asdata(plif_memwbrtnaddr_l_1),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(!plif_memwbpcsrc_l_1),
	.ena(\PCreg[1]~0_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(PCreg_1),
	.prn(vcc));
// synopsys translate_off
defparam \PCreg[1] .is_wysiwyg = "true";
defparam \PCreg[1] .power_up = "low";
// synopsys translate_on

// Location: FF_X50_Y32_N11
dffeas \PCreg[0] (
	.clk(CLK),
	.d(\PCreg[0]~feeder_combout ),
	.asdata(plif_memwbrtnaddr_l_0),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(!plif_memwbpcsrc_l_1),
	.ena(\PCreg[1]~0_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(PCreg_0),
	.prn(vcc));
// synopsys translate_off
defparam \PCreg[0] .is_wysiwyg = "true";
defparam \PCreg[0] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X52_Y33_N2
cycloneive_lcell_comb \pcif.rtnaddr[2]~0 (
// Equation(s):
// pcifrtnaddr_2 = PCreg_2 $ (VCC)
// \pcif.rtnaddr[2]~1  = CARRY(PCreg_2)

	.dataa(gnd),
	.datab(PCreg_2),
	.datac(gnd),
	.datad(vcc),
	.cin(gnd),
	.combout(pcifrtnaddr_2),
	.cout(\pcif.rtnaddr[2]~1 ));
// synopsys translate_off
defparam \pcif.rtnaddr[2]~0 .lut_mask = 16'h33CC;
defparam \pcif.rtnaddr[2]~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X52_Y33_N4
cycloneive_lcell_comb \pcif.rtnaddr[3]~2 (
// Equation(s):
// pcifrtnaddr_3 = (PCreg_3 & (!\pcif.rtnaddr[2]~1 )) # (!PCreg_3 & ((\pcif.rtnaddr[2]~1 ) # (GND)))
// \pcif.rtnaddr[3]~3  = CARRY((!\pcif.rtnaddr[2]~1 ) # (!PCreg_3))

	.dataa(gnd),
	.datab(PCreg_3),
	.datac(gnd),
	.datad(vcc),
	.cin(\pcif.rtnaddr[2]~1 ),
	.combout(pcifrtnaddr_3),
	.cout(\pcif.rtnaddr[3]~3 ));
// synopsys translate_off
defparam \pcif.rtnaddr[3]~2 .lut_mask = 16'h3C3F;
defparam \pcif.rtnaddr[3]~2 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X52_Y33_N6
cycloneive_lcell_comb \pcif.rtnaddr[4]~4 (
// Equation(s):
// pcifrtnaddr_4 = (PCreg_4 & (\pcif.rtnaddr[3]~3  $ (GND))) # (!PCreg_4 & (!\pcif.rtnaddr[3]~3  & VCC))
// \pcif.rtnaddr[4]~5  = CARRY((PCreg_4 & !\pcif.rtnaddr[3]~3 ))

	.dataa(gnd),
	.datab(PCreg_4),
	.datac(gnd),
	.datad(vcc),
	.cin(\pcif.rtnaddr[3]~3 ),
	.combout(pcifrtnaddr_4),
	.cout(\pcif.rtnaddr[4]~5 ));
// synopsys translate_off
defparam \pcif.rtnaddr[4]~4 .lut_mask = 16'hC30C;
defparam \pcif.rtnaddr[4]~4 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X52_Y33_N8
cycloneive_lcell_comb \pcif.rtnaddr[5]~6 (
// Equation(s):
// pcifrtnaddr_5 = (PCreg_5 & (!\pcif.rtnaddr[4]~5 )) # (!PCreg_5 & ((\pcif.rtnaddr[4]~5 ) # (GND)))
// \pcif.rtnaddr[5]~7  = CARRY((!\pcif.rtnaddr[4]~5 ) # (!PCreg_5))

	.dataa(PCreg_5),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\pcif.rtnaddr[4]~5 ),
	.combout(pcifrtnaddr_5),
	.cout(\pcif.rtnaddr[5]~7 ));
// synopsys translate_off
defparam \pcif.rtnaddr[5]~6 .lut_mask = 16'h5A5F;
defparam \pcif.rtnaddr[5]~6 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X52_Y33_N10
cycloneive_lcell_comb \pcif.rtnaddr[6]~8 (
// Equation(s):
// pcifrtnaddr_6 = (PCreg_6 & (\pcif.rtnaddr[5]~7  $ (GND))) # (!PCreg_6 & (!\pcif.rtnaddr[5]~7  & VCC))
// \pcif.rtnaddr[6]~9  = CARRY((PCreg_6 & !\pcif.rtnaddr[5]~7 ))

	.dataa(gnd),
	.datab(PCreg_6),
	.datac(gnd),
	.datad(vcc),
	.cin(\pcif.rtnaddr[5]~7 ),
	.combout(pcifrtnaddr_6),
	.cout(\pcif.rtnaddr[6]~9 ));
// synopsys translate_off
defparam \pcif.rtnaddr[6]~8 .lut_mask = 16'hC30C;
defparam \pcif.rtnaddr[6]~8 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X52_Y33_N12
cycloneive_lcell_comb \pcif.rtnaddr[7]~10 (
// Equation(s):
// pcifrtnaddr_7 = (PCreg_7 & (!\pcif.rtnaddr[6]~9 )) # (!PCreg_7 & ((\pcif.rtnaddr[6]~9 ) # (GND)))
// \pcif.rtnaddr[7]~11  = CARRY((!\pcif.rtnaddr[6]~9 ) # (!PCreg_7))

	.dataa(PCreg_7),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\pcif.rtnaddr[6]~9 ),
	.combout(pcifrtnaddr_7),
	.cout(\pcif.rtnaddr[7]~11 ));
// synopsys translate_off
defparam \pcif.rtnaddr[7]~10 .lut_mask = 16'h5A5F;
defparam \pcif.rtnaddr[7]~10 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X52_Y33_N14
cycloneive_lcell_comb \pcif.rtnaddr[8]~12 (
// Equation(s):
// pcifrtnaddr_8 = (PCreg_8 & (\pcif.rtnaddr[7]~11  $ (GND))) # (!PCreg_8 & (!\pcif.rtnaddr[7]~11  & VCC))
// \pcif.rtnaddr[8]~13  = CARRY((PCreg_8 & !\pcif.rtnaddr[7]~11 ))

	.dataa(gnd),
	.datab(PCreg_8),
	.datac(gnd),
	.datad(vcc),
	.cin(\pcif.rtnaddr[7]~11 ),
	.combout(pcifrtnaddr_8),
	.cout(\pcif.rtnaddr[8]~13 ));
// synopsys translate_off
defparam \pcif.rtnaddr[8]~12 .lut_mask = 16'hC30C;
defparam \pcif.rtnaddr[8]~12 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X52_Y33_N16
cycloneive_lcell_comb \pcif.rtnaddr[9]~14 (
// Equation(s):
// pcifrtnaddr_9 = (PCreg_9 & (!\pcif.rtnaddr[8]~13 )) # (!PCreg_9 & ((\pcif.rtnaddr[8]~13 ) # (GND)))
// \pcif.rtnaddr[9]~15  = CARRY((!\pcif.rtnaddr[8]~13 ) # (!PCreg_9))

	.dataa(gnd),
	.datab(PCreg_9),
	.datac(gnd),
	.datad(vcc),
	.cin(\pcif.rtnaddr[8]~13 ),
	.combout(pcifrtnaddr_9),
	.cout(\pcif.rtnaddr[9]~15 ));
// synopsys translate_off
defparam \pcif.rtnaddr[9]~14 .lut_mask = 16'h3C3F;
defparam \pcif.rtnaddr[9]~14 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X52_Y33_N18
cycloneive_lcell_comb \pcif.rtnaddr[10]~16 (
// Equation(s):
// pcifrtnaddr_10 = (PCreg_10 & (\pcif.rtnaddr[9]~15  $ (GND))) # (!PCreg_10 & (!\pcif.rtnaddr[9]~15  & VCC))
// \pcif.rtnaddr[10]~17  = CARRY((PCreg_10 & !\pcif.rtnaddr[9]~15 ))

	.dataa(PCreg_10),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\pcif.rtnaddr[9]~15 ),
	.combout(pcifrtnaddr_10),
	.cout(\pcif.rtnaddr[10]~17 ));
// synopsys translate_off
defparam \pcif.rtnaddr[10]~16 .lut_mask = 16'hA50A;
defparam \pcif.rtnaddr[10]~16 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X52_Y33_N20
cycloneive_lcell_comb \pcif.rtnaddr[11]~18 (
// Equation(s):
// pcifrtnaddr_11 = (PCreg_11 & (!\pcif.rtnaddr[10]~17 )) # (!PCreg_11 & ((\pcif.rtnaddr[10]~17 ) # (GND)))
// \pcif.rtnaddr[11]~19  = CARRY((!\pcif.rtnaddr[10]~17 ) # (!PCreg_11))

	.dataa(gnd),
	.datab(PCreg_11),
	.datac(gnd),
	.datad(vcc),
	.cin(\pcif.rtnaddr[10]~17 ),
	.combout(pcifrtnaddr_11),
	.cout(\pcif.rtnaddr[11]~19 ));
// synopsys translate_off
defparam \pcif.rtnaddr[11]~18 .lut_mask = 16'h3C3F;
defparam \pcif.rtnaddr[11]~18 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X52_Y33_N22
cycloneive_lcell_comb \pcif.rtnaddr[12]~20 (
// Equation(s):
// pcifrtnaddr_12 = (PCreg_12 & (\pcif.rtnaddr[11]~19  $ (GND))) # (!PCreg_12 & (!\pcif.rtnaddr[11]~19  & VCC))
// \pcif.rtnaddr[12]~21  = CARRY((PCreg_12 & !\pcif.rtnaddr[11]~19 ))

	.dataa(gnd),
	.datab(PCreg_12),
	.datac(gnd),
	.datad(vcc),
	.cin(\pcif.rtnaddr[11]~19 ),
	.combout(pcifrtnaddr_12),
	.cout(\pcif.rtnaddr[12]~21 ));
// synopsys translate_off
defparam \pcif.rtnaddr[12]~20 .lut_mask = 16'hC30C;
defparam \pcif.rtnaddr[12]~20 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X52_Y33_N24
cycloneive_lcell_comb \pcif.rtnaddr[13]~22 (
// Equation(s):
// pcifrtnaddr_13 = (PCreg_13 & (!\pcif.rtnaddr[12]~21 )) # (!PCreg_13 & ((\pcif.rtnaddr[12]~21 ) # (GND)))
// \pcif.rtnaddr[13]~23  = CARRY((!\pcif.rtnaddr[12]~21 ) # (!PCreg_13))

	.dataa(PCreg_13),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\pcif.rtnaddr[12]~21 ),
	.combout(pcifrtnaddr_13),
	.cout(\pcif.rtnaddr[13]~23 ));
// synopsys translate_off
defparam \pcif.rtnaddr[13]~22 .lut_mask = 16'h5A5F;
defparam \pcif.rtnaddr[13]~22 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X52_Y33_N26
cycloneive_lcell_comb \pcif.rtnaddr[14]~24 (
// Equation(s):
// pcifrtnaddr_14 = (PCreg_14 & (\pcif.rtnaddr[13]~23  $ (GND))) # (!PCreg_14 & (!\pcif.rtnaddr[13]~23  & VCC))
// \pcif.rtnaddr[14]~25  = CARRY((PCreg_14 & !\pcif.rtnaddr[13]~23 ))

	.dataa(PCreg_14),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\pcif.rtnaddr[13]~23 ),
	.combout(pcifrtnaddr_14),
	.cout(\pcif.rtnaddr[14]~25 ));
// synopsys translate_off
defparam \pcif.rtnaddr[14]~24 .lut_mask = 16'hA50A;
defparam \pcif.rtnaddr[14]~24 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X52_Y33_N28
cycloneive_lcell_comb \pcif.rtnaddr[15]~26 (
// Equation(s):
// pcifrtnaddr_15 = (PCreg_15 & (!\pcif.rtnaddr[14]~25 )) # (!PCreg_15 & ((\pcif.rtnaddr[14]~25 ) # (GND)))
// \pcif.rtnaddr[15]~27  = CARRY((!\pcif.rtnaddr[14]~25 ) # (!PCreg_15))

	.dataa(PCreg_15),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\pcif.rtnaddr[14]~25 ),
	.combout(pcifrtnaddr_15),
	.cout(\pcif.rtnaddr[15]~27 ));
// synopsys translate_off
defparam \pcif.rtnaddr[15]~26 .lut_mask = 16'h5A5F;
defparam \pcif.rtnaddr[15]~26 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X52_Y33_N30
cycloneive_lcell_comb \pcif.rtnaddr[16]~28 (
// Equation(s):
// pcifrtnaddr_16 = (PCreg_16 & (\pcif.rtnaddr[15]~27  $ (GND))) # (!PCreg_16 & (!\pcif.rtnaddr[15]~27  & VCC))
// \pcif.rtnaddr[16]~29  = CARRY((PCreg_16 & !\pcif.rtnaddr[15]~27 ))

	.dataa(PCreg_16),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\pcif.rtnaddr[15]~27 ),
	.combout(pcifrtnaddr_16),
	.cout(\pcif.rtnaddr[16]~29 ));
// synopsys translate_off
defparam \pcif.rtnaddr[16]~28 .lut_mask = 16'hA50A;
defparam \pcif.rtnaddr[16]~28 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X52_Y32_N0
cycloneive_lcell_comb \pcif.rtnaddr[17]~30 (
// Equation(s):
// pcifrtnaddr_17 = (PCreg_17 & (!\pcif.rtnaddr[16]~29 )) # (!PCreg_17 & ((\pcif.rtnaddr[16]~29 ) # (GND)))
// \pcif.rtnaddr[17]~31  = CARRY((!\pcif.rtnaddr[16]~29 ) # (!PCreg_17))

	.dataa(PCreg_17),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\pcif.rtnaddr[16]~29 ),
	.combout(pcifrtnaddr_17),
	.cout(\pcif.rtnaddr[17]~31 ));
// synopsys translate_off
defparam \pcif.rtnaddr[17]~30 .lut_mask = 16'h5A5F;
defparam \pcif.rtnaddr[17]~30 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X52_Y32_N2
cycloneive_lcell_comb \pcif.rtnaddr[18]~32 (
// Equation(s):
// pcifrtnaddr_18 = (PCreg_18 & (\pcif.rtnaddr[17]~31  $ (GND))) # (!PCreg_18 & (!\pcif.rtnaddr[17]~31  & VCC))
// \pcif.rtnaddr[18]~33  = CARRY((PCreg_18 & !\pcif.rtnaddr[17]~31 ))

	.dataa(gnd),
	.datab(PCreg_18),
	.datac(gnd),
	.datad(vcc),
	.cin(\pcif.rtnaddr[17]~31 ),
	.combout(pcifrtnaddr_18),
	.cout(\pcif.rtnaddr[18]~33 ));
// synopsys translate_off
defparam \pcif.rtnaddr[18]~32 .lut_mask = 16'hC30C;
defparam \pcif.rtnaddr[18]~32 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X52_Y32_N4
cycloneive_lcell_comb \pcif.rtnaddr[19]~34 (
// Equation(s):
// pcifrtnaddr_19 = (PCreg_19 & (!\pcif.rtnaddr[18]~33 )) # (!PCreg_19 & ((\pcif.rtnaddr[18]~33 ) # (GND)))
// \pcif.rtnaddr[19]~35  = CARRY((!\pcif.rtnaddr[18]~33 ) # (!PCreg_19))

	.dataa(gnd),
	.datab(PCreg_19),
	.datac(gnd),
	.datad(vcc),
	.cin(\pcif.rtnaddr[18]~33 ),
	.combout(pcifrtnaddr_19),
	.cout(\pcif.rtnaddr[19]~35 ));
// synopsys translate_off
defparam \pcif.rtnaddr[19]~34 .lut_mask = 16'h3C3F;
defparam \pcif.rtnaddr[19]~34 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X52_Y32_N6
cycloneive_lcell_comb \pcif.rtnaddr[20]~36 (
// Equation(s):
// pcifrtnaddr_20 = (PCreg_20 & (\pcif.rtnaddr[19]~35  $ (GND))) # (!PCreg_20 & (!\pcif.rtnaddr[19]~35  & VCC))
// \pcif.rtnaddr[20]~37  = CARRY((PCreg_20 & !\pcif.rtnaddr[19]~35 ))

	.dataa(gnd),
	.datab(PCreg_20),
	.datac(gnd),
	.datad(vcc),
	.cin(\pcif.rtnaddr[19]~35 ),
	.combout(pcifrtnaddr_20),
	.cout(\pcif.rtnaddr[20]~37 ));
// synopsys translate_off
defparam \pcif.rtnaddr[20]~36 .lut_mask = 16'hC30C;
defparam \pcif.rtnaddr[20]~36 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X52_Y32_N8
cycloneive_lcell_comb \pcif.rtnaddr[21]~38 (
// Equation(s):
// pcifrtnaddr_21 = (PCreg_21 & (!\pcif.rtnaddr[20]~37 )) # (!PCreg_21 & ((\pcif.rtnaddr[20]~37 ) # (GND)))
// \pcif.rtnaddr[21]~39  = CARRY((!\pcif.rtnaddr[20]~37 ) # (!PCreg_21))

	.dataa(PCreg_21),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\pcif.rtnaddr[20]~37 ),
	.combout(pcifrtnaddr_21),
	.cout(\pcif.rtnaddr[21]~39 ));
// synopsys translate_off
defparam \pcif.rtnaddr[21]~38 .lut_mask = 16'h5A5F;
defparam \pcif.rtnaddr[21]~38 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X52_Y32_N10
cycloneive_lcell_comb \pcif.rtnaddr[22]~40 (
// Equation(s):
// pcifrtnaddr_22 = (PCreg_22 & (\pcif.rtnaddr[21]~39  $ (GND))) # (!PCreg_22 & (!\pcif.rtnaddr[21]~39  & VCC))
// \pcif.rtnaddr[22]~41  = CARRY((PCreg_22 & !\pcif.rtnaddr[21]~39 ))

	.dataa(gnd),
	.datab(PCreg_22),
	.datac(gnd),
	.datad(vcc),
	.cin(\pcif.rtnaddr[21]~39 ),
	.combout(pcifrtnaddr_22),
	.cout(\pcif.rtnaddr[22]~41 ));
// synopsys translate_off
defparam \pcif.rtnaddr[22]~40 .lut_mask = 16'hC30C;
defparam \pcif.rtnaddr[22]~40 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X52_Y32_N12
cycloneive_lcell_comb \pcif.rtnaddr[23]~42 (
// Equation(s):
// pcifrtnaddr_23 = (PCreg_23 & (!\pcif.rtnaddr[22]~41 )) # (!PCreg_23 & ((\pcif.rtnaddr[22]~41 ) # (GND)))
// \pcif.rtnaddr[23]~43  = CARRY((!\pcif.rtnaddr[22]~41 ) # (!PCreg_23))

	.dataa(PCreg_23),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\pcif.rtnaddr[22]~41 ),
	.combout(pcifrtnaddr_23),
	.cout(\pcif.rtnaddr[23]~43 ));
// synopsys translate_off
defparam \pcif.rtnaddr[23]~42 .lut_mask = 16'h5A5F;
defparam \pcif.rtnaddr[23]~42 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X52_Y32_N14
cycloneive_lcell_comb \pcif.rtnaddr[24]~44 (
// Equation(s):
// pcifrtnaddr_24 = (PCreg_24 & (\pcif.rtnaddr[23]~43  $ (GND))) # (!PCreg_24 & (!\pcif.rtnaddr[23]~43  & VCC))
// \pcif.rtnaddr[24]~45  = CARRY((PCreg_24 & !\pcif.rtnaddr[23]~43 ))

	.dataa(gnd),
	.datab(PCreg_24),
	.datac(gnd),
	.datad(vcc),
	.cin(\pcif.rtnaddr[23]~43 ),
	.combout(pcifrtnaddr_24),
	.cout(\pcif.rtnaddr[24]~45 ));
// synopsys translate_off
defparam \pcif.rtnaddr[24]~44 .lut_mask = 16'hC30C;
defparam \pcif.rtnaddr[24]~44 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X52_Y32_N16
cycloneive_lcell_comb \pcif.rtnaddr[25]~46 (
// Equation(s):
// pcifrtnaddr_25 = (PCreg_25 & (!\pcif.rtnaddr[24]~45 )) # (!PCreg_25 & ((\pcif.rtnaddr[24]~45 ) # (GND)))
// \pcif.rtnaddr[25]~47  = CARRY((!\pcif.rtnaddr[24]~45 ) # (!PCreg_25))

	.dataa(gnd),
	.datab(PCreg_25),
	.datac(gnd),
	.datad(vcc),
	.cin(\pcif.rtnaddr[24]~45 ),
	.combout(pcifrtnaddr_25),
	.cout(\pcif.rtnaddr[25]~47 ));
// synopsys translate_off
defparam \pcif.rtnaddr[25]~46 .lut_mask = 16'h3C3F;
defparam \pcif.rtnaddr[25]~46 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X52_Y32_N18
cycloneive_lcell_comb \pcif.rtnaddr[26]~48 (
// Equation(s):
// pcifrtnaddr_26 = (PCreg_26 & (\pcif.rtnaddr[25]~47  $ (GND))) # (!PCreg_26 & (!\pcif.rtnaddr[25]~47  & VCC))
// \pcif.rtnaddr[26]~49  = CARRY((PCreg_26 & !\pcif.rtnaddr[25]~47 ))

	.dataa(PCreg_26),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\pcif.rtnaddr[25]~47 ),
	.combout(pcifrtnaddr_26),
	.cout(\pcif.rtnaddr[26]~49 ));
// synopsys translate_off
defparam \pcif.rtnaddr[26]~48 .lut_mask = 16'hA50A;
defparam \pcif.rtnaddr[26]~48 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X52_Y32_N20
cycloneive_lcell_comb \pcif.rtnaddr[27]~50 (
// Equation(s):
// pcifrtnaddr_27 = (PCreg_27 & (!\pcif.rtnaddr[26]~49 )) # (!PCreg_27 & ((\pcif.rtnaddr[26]~49 ) # (GND)))
// \pcif.rtnaddr[27]~51  = CARRY((!\pcif.rtnaddr[26]~49 ) # (!PCreg_27))

	.dataa(gnd),
	.datab(PCreg_27),
	.datac(gnd),
	.datad(vcc),
	.cin(\pcif.rtnaddr[26]~49 ),
	.combout(pcifrtnaddr_27),
	.cout(\pcif.rtnaddr[27]~51 ));
// synopsys translate_off
defparam \pcif.rtnaddr[27]~50 .lut_mask = 16'h3C3F;
defparam \pcif.rtnaddr[27]~50 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X52_Y32_N22
cycloneive_lcell_comb \pcif.rtnaddr[28]~52 (
// Equation(s):
// pcifrtnaddr_28 = (PCreg_28 & (\pcif.rtnaddr[27]~51  $ (GND))) # (!PCreg_28 & (!\pcif.rtnaddr[27]~51  & VCC))
// \pcif.rtnaddr[28]~53  = CARRY((PCreg_28 & !\pcif.rtnaddr[27]~51 ))

	.dataa(PCreg_28),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\pcif.rtnaddr[27]~51 ),
	.combout(pcifrtnaddr_28),
	.cout(\pcif.rtnaddr[28]~53 ));
// synopsys translate_off
defparam \pcif.rtnaddr[28]~52 .lut_mask = 16'hA50A;
defparam \pcif.rtnaddr[28]~52 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X52_Y32_N24
cycloneive_lcell_comb \pcif.rtnaddr[29]~54 (
// Equation(s):
// pcifrtnaddr_29 = (PCreg_29 & (!\pcif.rtnaddr[28]~53 )) # (!PCreg_29 & ((\pcif.rtnaddr[28]~53 ) # (GND)))
// \pcif.rtnaddr[29]~55  = CARRY((!\pcif.rtnaddr[28]~53 ) # (!PCreg_29))

	.dataa(gnd),
	.datab(PCreg_29),
	.datac(gnd),
	.datad(vcc),
	.cin(\pcif.rtnaddr[28]~53 ),
	.combout(pcifrtnaddr_29),
	.cout(\pcif.rtnaddr[29]~55 ));
// synopsys translate_off
defparam \pcif.rtnaddr[29]~54 .lut_mask = 16'h3C3F;
defparam \pcif.rtnaddr[29]~54 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X52_Y32_N26
cycloneive_lcell_comb \pcif.rtnaddr[30]~56 (
// Equation(s):
// pcifrtnaddr_30 = (PCreg_30 & (\pcif.rtnaddr[29]~55  $ (GND))) # (!PCreg_30 & (!\pcif.rtnaddr[29]~55  & VCC))
// \pcif.rtnaddr[30]~57  = CARRY((PCreg_30 & !\pcif.rtnaddr[29]~55 ))

	.dataa(PCreg_30),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\pcif.rtnaddr[29]~55 ),
	.combout(pcifrtnaddr_30),
	.cout(\pcif.rtnaddr[30]~57 ));
// synopsys translate_off
defparam \pcif.rtnaddr[30]~56 .lut_mask = 16'hA50A;
defparam \pcif.rtnaddr[30]~56 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X52_Y32_N28
cycloneive_lcell_comb \pcif.rtnaddr[31]~58 (
// Equation(s):
// pcifrtnaddr_31 = PCreg_31 $ (\pcif.rtnaddr[30]~57 )

	.dataa(PCreg_31),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.cin(\pcif.rtnaddr[30]~57 ),
	.combout(pcifrtnaddr_31),
	.cout());
// synopsys translate_off
defparam \pcif.rtnaddr[31]~58 .lut_mask = 16'h5A5A;
defparam \pcif.rtnaddr[31]~58 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: FF_X54_Y35_N1
dffeas \PCreg[3] (
	.clk(CLK),
	.d(\PCregN~3_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\pcif.rambusy ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(PCreg_3),
	.prn(vcc));
// synopsys translate_off
defparam \PCreg[3] .is_wysiwyg = "true";
defparam \PCreg[3] .power_up = "low";
// synopsys translate_on

// Location: FF_X54_Y35_N3
dffeas \PCreg[2] (
	.clk(CLK),
	.d(\PCregN~5_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\pcif.rambusy ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(PCreg_2),
	.prn(vcc));
// synopsys translate_off
defparam \PCreg[2] .is_wysiwyg = "true";
defparam \PCreg[2] .power_up = "low";
// synopsys translate_on

// Location: FF_X49_Y34_N31
dffeas \PCreg[5] (
	.clk(CLK),
	.d(\PCregN~7_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\pcif.rambusy ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(PCreg_5),
	.prn(vcc));
// synopsys translate_off
defparam \PCreg[5] .is_wysiwyg = "true";
defparam \PCreg[5] .power_up = "low";
// synopsys translate_on

// Location: FF_X49_Y34_N29
dffeas \PCreg[4] (
	.clk(CLK),
	.d(\PCregN~9_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\pcif.rambusy ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(PCreg_4),
	.prn(vcc));
// synopsys translate_off
defparam \PCreg[4] .is_wysiwyg = "true";
defparam \PCreg[4] .power_up = "low";
// synopsys translate_on

// Location: FF_X55_Y34_N21
dffeas \PCreg[7] (
	.clk(CLK),
	.d(\PCregN~11_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\pcif.rambusy ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(PCreg_7),
	.prn(vcc));
// synopsys translate_off
defparam \PCreg[7] .is_wysiwyg = "true";
defparam \PCreg[7] .power_up = "low";
// synopsys translate_on

// Location: FF_X55_Y34_N31
dffeas \PCreg[6] (
	.clk(CLK),
	.d(\PCregN~13_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\pcif.rambusy ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(PCreg_6),
	.prn(vcc));
// synopsys translate_off
defparam \PCreg[6] .is_wysiwyg = "true";
defparam \PCreg[6] .power_up = "low";
// synopsys translate_on

// Location: FF_X53_Y33_N13
dffeas \PCreg[9] (
	.clk(CLK),
	.d(\PCregN~15_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\pcif.rambusy ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(PCreg_9),
	.prn(vcc));
// synopsys translate_off
defparam \PCreg[9] .is_wysiwyg = "true";
defparam \PCreg[9] .power_up = "low";
// synopsys translate_on

// Location: FF_X54_Y33_N31
dffeas \PCreg[8] (
	.clk(CLK),
	.d(\PCregN~17_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\pcif.rambusy ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(PCreg_8),
	.prn(vcc));
// synopsys translate_off
defparam \PCreg[8] .is_wysiwyg = "true";
defparam \PCreg[8] .power_up = "low";
// synopsys translate_on

// Location: FF_X55_Y34_N15
dffeas \PCreg[11] (
	.clk(CLK),
	.d(\PCregN~19_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\pcif.rambusy ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(PCreg_11),
	.prn(vcc));
// synopsys translate_off
defparam \PCreg[11] .is_wysiwyg = "true";
defparam \PCreg[11] .power_up = "low";
// synopsys translate_on

// Location: FF_X55_Y34_N1
dffeas \PCreg[10] (
	.clk(CLK),
	.d(\PCregN~21_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\pcif.rambusy ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(PCreg_10),
	.prn(vcc));
// synopsys translate_off
defparam \PCreg[10] .is_wysiwyg = "true";
defparam \PCreg[10] .power_up = "low";
// synopsys translate_on

// Location: FF_X54_Y32_N9
dffeas \PCreg[13] (
	.clk(CLK),
	.d(\PCregN~23_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\pcif.rambusy ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(PCreg_13),
	.prn(vcc));
// synopsys translate_off
defparam \PCreg[13] .is_wysiwyg = "true";
defparam \PCreg[13] .power_up = "low";
// synopsys translate_on

// Location: FF_X54_Y32_N19
dffeas \PCreg[12] (
	.clk(CLK),
	.d(\PCregN~25_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\pcif.rambusy ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(PCreg_12),
	.prn(vcc));
// synopsys translate_off
defparam \PCreg[12] .is_wysiwyg = "true";
defparam \PCreg[12] .power_up = "low";
// synopsys translate_on

// Location: FF_X52_Y34_N5
dffeas \PCreg[15] (
	.clk(CLK),
	.d(\PCregN~27_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\pcif.rambusy ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(PCreg_15),
	.prn(vcc));
// synopsys translate_off
defparam \PCreg[15] .is_wysiwyg = "true";
defparam \PCreg[15] .power_up = "low";
// synopsys translate_on

// Location: FF_X52_Y34_N31
dffeas \PCreg[14] (
	.clk(CLK),
	.d(\PCreg[14]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\pcif.rambusy ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(PCreg_14),
	.prn(vcc));
// synopsys translate_off
defparam \PCreg[14] .is_wysiwyg = "true";
defparam \PCreg[14] .power_up = "low";
// synopsys translate_on

// Location: FF_X50_Y34_N5
dffeas \PCreg[17] (
	.clk(CLK),
	.d(\PCregN~31_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\pcif.rambusy ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(PCreg_17),
	.prn(vcc));
// synopsys translate_off
defparam \PCreg[17] .is_wysiwyg = "true";
defparam \PCreg[17] .power_up = "low";
// synopsys translate_on

// Location: FF_X50_Y34_N1
dffeas \PCreg[16] (
	.clk(CLK),
	.d(\PCregN~33_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\pcif.rambusy ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(PCreg_16),
	.prn(vcc));
// synopsys translate_off
defparam \PCreg[16] .is_wysiwyg = "true";
defparam \PCreg[16] .power_up = "low";
// synopsys translate_on

// Location: FF_X54_Y33_N1
dffeas \PCreg[19] (
	.clk(CLK),
	.d(\PCregN~35_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\pcif.rambusy ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(PCreg_19),
	.prn(vcc));
// synopsys translate_off
defparam \PCreg[19] .is_wysiwyg = "true";
defparam \PCreg[19] .power_up = "low";
// synopsys translate_on

// Location: FF_X54_Y33_N5
dffeas \PCreg[18] (
	.clk(CLK),
	.d(\PCregN~37_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\pcif.rambusy ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(PCreg_18),
	.prn(vcc));
// synopsys translate_off
defparam \PCreg[18] .is_wysiwyg = "true";
defparam \PCreg[18] .power_up = "low";
// synopsys translate_on

// Location: FF_X52_Y34_N17
dffeas \PCreg[21] (
	.clk(CLK),
	.d(\PCregN~39_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\pcif.rambusy ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(PCreg_21),
	.prn(vcc));
// synopsys translate_off
defparam \PCreg[21] .is_wysiwyg = "true";
defparam \PCreg[21] .power_up = "low";
// synopsys translate_on

// Location: FF_X56_Y34_N13
dffeas \PCreg[20] (
	.clk(CLK),
	.d(\PCregN~41_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\pcif.rambusy ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(PCreg_20),
	.prn(vcc));
// synopsys translate_off
defparam \PCreg[20] .is_wysiwyg = "true";
defparam \PCreg[20] .power_up = "low";
// synopsys translate_on

// Location: FF_X52_Y32_N31
dffeas \PCreg[23] (
	.clk(CLK),
	.d(\PCregN~43_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\pcif.rambusy ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(PCreg_23),
	.prn(vcc));
// synopsys translate_off
defparam \PCreg[23] .is_wysiwyg = "true";
defparam \PCreg[23] .power_up = "low";
// synopsys translate_on

// Location: FF_X52_Y34_N15
dffeas \PCreg[22] (
	.clk(CLK),
	.d(\PCregN~45_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\pcif.rambusy ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(PCreg_22),
	.prn(vcc));
// synopsys translate_off
defparam \PCreg[22] .is_wysiwyg = "true";
defparam \PCreg[22] .power_up = "low";
// synopsys translate_on

// Location: FF_X54_Y35_N19
dffeas \PCreg[25] (
	.clk(CLK),
	.d(\PCregN~47_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\pcif.rambusy ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(PCreg_25),
	.prn(vcc));
// synopsys translate_off
defparam \PCreg[25] .is_wysiwyg = "true";
defparam \PCreg[25] .power_up = "low";
// synopsys translate_on

// Location: FF_X53_Y33_N7
dffeas \PCreg[24] (
	.clk(CLK),
	.d(\PCregN~49_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\pcif.rambusy ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(PCreg_24),
	.prn(vcc));
// synopsys translate_off
defparam \PCreg[24] .is_wysiwyg = "true";
defparam \PCreg[24] .power_up = "low";
// synopsys translate_on

// Location: FF_X53_Y33_N29
dffeas \PCreg[27] (
	.clk(CLK),
	.d(\PCregN~51_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\pcif.rambusy ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(PCreg_27),
	.prn(vcc));
// synopsys translate_off
defparam \PCreg[27] .is_wysiwyg = "true";
defparam \PCreg[27] .power_up = "low";
// synopsys translate_on

// Location: FF_X55_Y33_N13
dffeas \PCreg[26] (
	.clk(CLK),
	.d(\PCregN~53_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\pcif.rambusy ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(PCreg_26),
	.prn(vcc));
// synopsys translate_off
defparam \PCreg[26] .is_wysiwyg = "true";
defparam \PCreg[26] .power_up = "low";
// synopsys translate_on

// Location: FF_X50_Y34_N7
dffeas \PCreg[29] (
	.clk(CLK),
	.d(\PCregN~55_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\pcif.rambusy ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(PCreg_29),
	.prn(vcc));
// synopsys translate_off
defparam \PCreg[29] .is_wysiwyg = "true";
defparam \PCreg[29] .power_up = "low";
// synopsys translate_on

// Location: FF_X50_Y34_N15
dffeas \PCreg[28] (
	.clk(CLK),
	.d(\PCregN~57_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\pcif.rambusy ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(PCreg_28),
	.prn(vcc));
// synopsys translate_off
defparam \PCreg[28] .is_wysiwyg = "true";
defparam \PCreg[28] .power_up = "low";
// synopsys translate_on

// Location: FF_X52_Y34_N21
dffeas \PCreg[31] (
	.clk(CLK),
	.d(\PCregN~59_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\pcif.rambusy ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(PCreg_31),
	.prn(vcc));
// synopsys translate_off
defparam \PCreg[31] .is_wysiwyg = "true";
defparam \PCreg[31] .power_up = "low";
// synopsys translate_on

// Location: FF_X56_Y34_N27
dffeas \PCreg[30] (
	.clk(CLK),
	.d(\PCregN~61_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\pcif.rambusy ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(PCreg_30),
	.prn(vcc));
// synopsys translate_off
defparam \PCreg[30] .is_wysiwyg = "true";
defparam \PCreg[30] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X53_Y31_N0
cycloneive_lcell_comb \PCregN~0 (
// Equation(s):
// \PCregN~0_combout  = (plif_memwbporto_l_1 & \pcsrc~0_combout )

	.dataa(gnd),
	.datab(plif_memwbporto_l_1),
	.datac(pcsrc),
	.datad(gnd),
	.cin(gnd),
	.combout(\PCregN~0_combout ),
	.cout());
// synopsys translate_off
defparam \PCregN~0 .lut_mask = 16'hC0C0;
defparam \PCregN~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X50_Y32_N24
cycloneive_lcell_comb \PCreg[1]~feeder (
// Equation(s):
// \PCreg[1]~feeder_combout  = \PCregN~0_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(\PCregN~0_combout ),
	.cin(gnd),
	.combout(\PCreg[1]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \PCreg[1]~feeder .lut_mask = 16'hFF00;
defparam \PCreg[1]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X50_Y32_N0
cycloneive_lcell_comb \PCreg[1]~0 (
// Equation(s):
// \PCreg[1]~0_combout  = (!always0 & (ifid_en & ((\pcsrc~0_combout ) # (plif_memwbpcsrc_l_1))))

	.dataa(pcsrc),
	.datab(always0),
	.datac(plif_memwbpcsrc_l_1),
	.datad(ifid_en),
	.cin(gnd),
	.combout(\PCreg[1]~0_combout ),
	.cout());
// synopsys translate_off
defparam \PCreg[1]~0 .lut_mask = 16'h3200;
defparam \PCreg[1]~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y31_N2
cycloneive_lcell_comb \PCregN~1 (
// Equation(s):
// \PCregN~1_combout  = (\pcsrc~0_combout  & plif_memwbporto_l_0)

	.dataa(gnd),
	.datab(gnd),
	.datac(pcsrc),
	.datad(plif_memwbporto_l_0),
	.cin(gnd),
	.combout(\PCregN~1_combout ),
	.cout());
// synopsys translate_off
defparam \PCregN~1 .lut_mask = 16'hF000;
defparam \PCregN~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X50_Y32_N10
cycloneive_lcell_comb \PCreg[0]~feeder (
// Equation(s):
// \PCreg[0]~feeder_combout  = \PCregN~1_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(\PCregN~1_combout ),
	.cin(gnd),
	.combout(\PCreg[0]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \PCreg[0]~feeder .lut_mask = 16'hFF00;
defparam \PCreg[0]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y32_N2
cycloneive_lcell_comb \Add1~0 (
// Equation(s):
// \Add1~0_combout  = (plif_memwbrtnaddr_l_2 & (plif_memwbextimm_l_0 $ (VCC))) # (!plif_memwbrtnaddr_l_2 & (plif_memwbextimm_l_0 & VCC))
// \Add1~1  = CARRY((plif_memwbrtnaddr_l_2 & plif_memwbextimm_l_0))

	.dataa(plif_memwbrtnaddr_l_2),
	.datab(plif_memwbextimm_l_0),
	.datac(gnd),
	.datad(vcc),
	.cin(gnd),
	.combout(\Add1~0_combout ),
	.cout(\Add1~1 ));
// synopsys translate_off
defparam \Add1~0 .lut_mask = 16'h6688;
defparam \Add1~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y32_N4
cycloneive_lcell_comb \Add1~2 (
// Equation(s):
// \Add1~2_combout  = (plif_memwbrtnaddr_l_3 & ((plif_memwbextimm_l_1 & (\Add1~1  & VCC)) # (!plif_memwbextimm_l_1 & (!\Add1~1 )))) # (!plif_memwbrtnaddr_l_3 & ((plif_memwbextimm_l_1 & (!\Add1~1 )) # (!plif_memwbextimm_l_1 & ((\Add1~1 ) # (GND)))))
// \Add1~3  = CARRY((plif_memwbrtnaddr_l_3 & (!plif_memwbextimm_l_1 & !\Add1~1 )) # (!plif_memwbrtnaddr_l_3 & ((!\Add1~1 ) # (!plif_memwbextimm_l_1))))

	.dataa(plif_memwbrtnaddr_l_3),
	.datab(plif_memwbextimm_l_1),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add1~1 ),
	.combout(\Add1~2_combout ),
	.cout(\Add1~3 ));
// synopsys translate_off
defparam \Add1~2 .lut_mask = 16'h9617;
defparam \Add1~2 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X53_Y35_N26
cycloneive_lcell_comb \PCregN~2 (
// Equation(s):
// \PCregN~2_combout  = (\pcsrc~0_combout  & ((\Add1~2_combout ) # ((plif_memwbpcsrc_l_1)))) # (!\pcsrc~0_combout  & (((!plif_memwbpcsrc_l_1 & pcifrtnaddr_3))))

	.dataa(pcsrc),
	.datab(\Add1~2_combout ),
	.datac(plif_memwbpcsrc_l_1),
	.datad(pcifrtnaddr_3),
	.cin(gnd),
	.combout(\PCregN~2_combout ),
	.cout());
// synopsys translate_off
defparam \PCregN~2 .lut_mask = 16'hADA8;
defparam \PCregN~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y35_N0
cycloneive_lcell_comb \PCregN~3 (
// Equation(s):
// \PCregN~3_combout  = (plif_memwbpcsrc_l_1 & ((\PCregN~2_combout  & (plif_memwbporto_l_3)) # (!\PCregN~2_combout  & ((plif_memwbjaddr_l_1))))) # (!plif_memwbpcsrc_l_1 & (((\PCregN~2_combout ))))

	.dataa(plif_memwbporto_l_3),
	.datab(plif_memwbpcsrc_l_1),
	.datac(\PCregN~2_combout ),
	.datad(plif_memwbjaddr_l_1),
	.cin(gnd),
	.combout(\PCregN~3_combout ),
	.cout());
// synopsys translate_off
defparam \PCregN~3 .lut_mask = 16'hBCB0;
defparam \PCregN~3 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X52_Y33_N0
cycloneive_lcell_comb \PCregN~4 (
// Equation(s):
// \PCregN~4_combout  = (\pcsrc~0_combout  & (plif_memwbpcsrc_l_1)) # (!\pcsrc~0_combout  & ((plif_memwbpcsrc_l_1 & (plif_memwbjaddr_l_0)) # (!plif_memwbpcsrc_l_1 & ((pcifrtnaddr_2)))))

	.dataa(pcsrc),
	.datab(plif_memwbpcsrc_l_1),
	.datac(plif_memwbjaddr_l_0),
	.datad(pcifrtnaddr_2),
	.cin(gnd),
	.combout(\PCregN~4_combout ),
	.cout());
// synopsys translate_off
defparam \PCregN~4 .lut_mask = 16'hD9C8;
defparam \PCregN~4 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y35_N2
cycloneive_lcell_comb \PCregN~5 (
// Equation(s):
// \PCregN~5_combout  = (\PCregN~4_combout  & (((plif_memwbporto_l_2)) # (!\pcsrc~0_combout ))) # (!\PCregN~4_combout  & (\pcsrc~0_combout  & (\Add1~0_combout )))

	.dataa(\PCregN~4_combout ),
	.datab(pcsrc),
	.datac(\Add1~0_combout ),
	.datad(plif_memwbporto_l_2),
	.cin(gnd),
	.combout(\PCregN~5_combout ),
	.cout());
// synopsys translate_off
defparam \PCregN~5 .lut_mask = 16'hEA62;
defparam \PCregN~5 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y32_N6
cycloneive_lcell_comb \Add1~4 (
// Equation(s):
// \Add1~4_combout  = ((plif_memwbextimm_l_2 $ (plif_memwbrtnaddr_l_4 $ (!\Add1~3 )))) # (GND)
// \Add1~5  = CARRY((plif_memwbextimm_l_2 & ((plif_memwbrtnaddr_l_4) # (!\Add1~3 ))) # (!plif_memwbextimm_l_2 & (plif_memwbrtnaddr_l_4 & !\Add1~3 )))

	.dataa(plif_memwbextimm_l_2),
	.datab(plif_memwbrtnaddr_l_4),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add1~3 ),
	.combout(\Add1~4_combout ),
	.cout(\Add1~5 ));
// synopsys translate_off
defparam \Add1~4 .lut_mask = 16'h698E;
defparam \Add1~4 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X56_Y32_N8
cycloneive_lcell_comb \Add1~6 (
// Equation(s):
// \Add1~6_combout  = (plif_memwbrtnaddr_l_5 & ((plif_memwbextimm_l_3 & (\Add1~5  & VCC)) # (!plif_memwbextimm_l_3 & (!\Add1~5 )))) # (!plif_memwbrtnaddr_l_5 & ((plif_memwbextimm_l_3 & (!\Add1~5 )) # (!plif_memwbextimm_l_3 & ((\Add1~5 ) # (GND)))))
// \Add1~7  = CARRY((plif_memwbrtnaddr_l_5 & (!plif_memwbextimm_l_3 & !\Add1~5 )) # (!plif_memwbrtnaddr_l_5 & ((!\Add1~5 ) # (!plif_memwbextimm_l_3))))

	.dataa(plif_memwbrtnaddr_l_5),
	.datab(plif_memwbextimm_l_3),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add1~5 ),
	.combout(\Add1~6_combout ),
	.cout(\Add1~7 ));
// synopsys translate_off
defparam \Add1~6 .lut_mask = 16'h9617;
defparam \Add1~6 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X53_Y33_N16
cycloneive_lcell_comb \PCregN~6 (
// Equation(s):
// \PCregN~6_combout  = (\pcsrc~0_combout  & ((plif_memwbpcsrc_l_1) # ((\Add1~6_combout )))) # (!\pcsrc~0_combout  & (!plif_memwbpcsrc_l_1 & ((pcifrtnaddr_5))))

	.dataa(pcsrc),
	.datab(plif_memwbpcsrc_l_1),
	.datac(\Add1~6_combout ),
	.datad(pcifrtnaddr_5),
	.cin(gnd),
	.combout(\PCregN~6_combout ),
	.cout());
// synopsys translate_off
defparam \PCregN~6 .lut_mask = 16'hB9A8;
defparam \PCregN~6 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X49_Y34_N30
cycloneive_lcell_comb \PCregN~7 (
// Equation(s):
// \PCregN~7_combout  = (plif_memwbpcsrc_l_1 & ((\PCregN~6_combout  & ((plif_memwbporto_l_5))) # (!\PCregN~6_combout  & (plif_memwbjaddr_l_3)))) # (!plif_memwbpcsrc_l_1 & (((\PCregN~6_combout ))))

	.dataa(plif_memwbpcsrc_l_1),
	.datab(plif_memwbjaddr_l_3),
	.datac(\PCregN~6_combout ),
	.datad(plif_memwbporto_l_5),
	.cin(gnd),
	.combout(\PCregN~7_combout ),
	.cout());
// synopsys translate_off
defparam \PCregN~7 .lut_mask = 16'hF858;
defparam \PCregN~7 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X50_Y33_N24
cycloneive_lcell_comb \PCregN~8 (
// Equation(s):
// \PCregN~8_combout  = (plif_memwbpcsrc_l_1 & (((plif_memwbjaddr_l_2) # (\pcsrc~0_combout )))) # (!plif_memwbpcsrc_l_1 & (pcifrtnaddr_4 & ((!\pcsrc~0_combout ))))

	.dataa(pcifrtnaddr_4),
	.datab(plif_memwbpcsrc_l_1),
	.datac(plif_memwbjaddr_l_2),
	.datad(pcsrc),
	.cin(gnd),
	.combout(\PCregN~8_combout ),
	.cout());
// synopsys translate_off
defparam \PCregN~8 .lut_mask = 16'hCCE2;
defparam \PCregN~8 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X49_Y34_N28
cycloneive_lcell_comb \PCregN~9 (
// Equation(s):
// \PCregN~9_combout  = (\pcsrc~0_combout  & ((\PCregN~8_combout  & ((plif_memwbporto_l_4))) # (!\PCregN~8_combout  & (\Add1~4_combout )))) # (!\pcsrc~0_combout  & (((\PCregN~8_combout ))))

	.dataa(\Add1~4_combout ),
	.datab(pcsrc),
	.datac(\PCregN~8_combout ),
	.datad(plif_memwbporto_l_4),
	.cin(gnd),
	.combout(\PCregN~9_combout ),
	.cout());
// synopsys translate_off
defparam \PCregN~9 .lut_mask = 16'hF838;
defparam \PCregN~9 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y32_N10
cycloneive_lcell_comb \Add1~8 (
// Equation(s):
// \Add1~8_combout  = ((plif_memwbextimm_l_4 $ (plif_memwbrtnaddr_l_6 $ (!\Add1~7 )))) # (GND)
// \Add1~9  = CARRY((plif_memwbextimm_l_4 & ((plif_memwbrtnaddr_l_6) # (!\Add1~7 ))) # (!plif_memwbextimm_l_4 & (plif_memwbrtnaddr_l_6 & !\Add1~7 )))

	.dataa(plif_memwbextimm_l_4),
	.datab(plif_memwbrtnaddr_l_6),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add1~7 ),
	.combout(\Add1~8_combout ),
	.cout(\Add1~9 ));
// synopsys translate_off
defparam \Add1~8 .lut_mask = 16'h698E;
defparam \Add1~8 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X56_Y32_N12
cycloneive_lcell_comb \Add1~10 (
// Equation(s):
// \Add1~10_combout  = (plif_memwbrtnaddr_l_7 & ((plif_memwbextimm_l_5 & (\Add1~9  & VCC)) # (!plif_memwbextimm_l_5 & (!\Add1~9 )))) # (!plif_memwbrtnaddr_l_7 & ((plif_memwbextimm_l_5 & (!\Add1~9 )) # (!plif_memwbextimm_l_5 & ((\Add1~9 ) # (GND)))))
// \Add1~11  = CARRY((plif_memwbrtnaddr_l_7 & (!plif_memwbextimm_l_5 & !\Add1~9 )) # (!plif_memwbrtnaddr_l_7 & ((!\Add1~9 ) # (!plif_memwbextimm_l_5))))

	.dataa(plif_memwbrtnaddr_l_7),
	.datab(plif_memwbextimm_l_5),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add1~9 ),
	.combout(\Add1~10_combout ),
	.cout(\Add1~11 ));
// synopsys translate_off
defparam \Add1~10 .lut_mask = 16'h9617;
defparam \Add1~10 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X55_Y34_N22
cycloneive_lcell_comb \PCregN~10 (
// Equation(s):
// \PCregN~10_combout  = (\pcsrc~0_combout  & (((\Add1~10_combout ) # (plif_memwbpcsrc_l_1)))) # (!\pcsrc~0_combout  & (pcifrtnaddr_7 & ((!plif_memwbpcsrc_l_1))))

	.dataa(pcifrtnaddr_7),
	.datab(\Add1~10_combout ),
	.datac(pcsrc),
	.datad(plif_memwbpcsrc_l_1),
	.cin(gnd),
	.combout(\PCregN~10_combout ),
	.cout());
// synopsys translate_off
defparam \PCregN~10 .lut_mask = 16'hF0CA;
defparam \PCregN~10 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y34_N20
cycloneive_lcell_comb \PCregN~11 (
// Equation(s):
// \PCregN~11_combout  = (\PCregN~10_combout  & (((plif_memwbporto_l_7) # (!plif_memwbpcsrc_l_1)))) # (!\PCregN~10_combout  & (plif_memwbjaddr_l_5 & ((plif_memwbpcsrc_l_1))))

	.dataa(\PCregN~10_combout ),
	.datab(plif_memwbjaddr_l_5),
	.datac(plif_memwbporto_l_7),
	.datad(plif_memwbpcsrc_l_1),
	.cin(gnd),
	.combout(\PCregN~11_combout ),
	.cout());
// synopsys translate_off
defparam \PCregN~11 .lut_mask = 16'hE4AA;
defparam \PCregN~11 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X50_Y33_N10
cycloneive_lcell_comb \PCregN~12 (
// Equation(s):
// \PCregN~12_combout  = (plif_memwbpcsrc_l_1 & (((plif_memwbjaddr_l_4) # (\pcsrc~0_combout )))) # (!plif_memwbpcsrc_l_1 & (pcifrtnaddr_6 & ((!\pcsrc~0_combout ))))

	.dataa(pcifrtnaddr_6),
	.datab(plif_memwbpcsrc_l_1),
	.datac(plif_memwbjaddr_l_4),
	.datad(pcsrc),
	.cin(gnd),
	.combout(\PCregN~12_combout ),
	.cout());
// synopsys translate_off
defparam \PCregN~12 .lut_mask = 16'hCCE2;
defparam \PCregN~12 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y34_N30
cycloneive_lcell_comb \PCregN~13 (
// Equation(s):
// \PCregN~13_combout  = (\PCregN~12_combout  & (((plif_memwbporto_l_6) # (!\pcsrc~0_combout )))) # (!\PCregN~12_combout  & (\Add1~8_combout  & (\pcsrc~0_combout )))

	.dataa(\Add1~8_combout ),
	.datab(\PCregN~12_combout ),
	.datac(pcsrc),
	.datad(plif_memwbporto_l_6),
	.cin(gnd),
	.combout(\PCregN~13_combout ),
	.cout());
// synopsys translate_off
defparam \PCregN~13 .lut_mask = 16'hEC2C;
defparam \PCregN~13 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y32_N26
cycloneive_lcell_comb \PCregN~14 (
// Equation(s):
// \PCregN~14_combout  = (plif_memwbpcsrc_l_1 & (((\pcsrc~0_combout )))) # (!plif_memwbpcsrc_l_1 & ((\pcsrc~0_combout  & (\Add1~14_combout )) # (!\pcsrc~0_combout  & ((pcifrtnaddr_9)))))

	.dataa(\Add1~14_combout ),
	.datab(plif_memwbpcsrc_l_1),
	.datac(pcifrtnaddr_9),
	.datad(pcsrc),
	.cin(gnd),
	.combout(\PCregN~14_combout ),
	.cout());
// synopsys translate_off
defparam \PCregN~14 .lut_mask = 16'hEE30;
defparam \PCregN~14 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y33_N12
cycloneive_lcell_comb \PCregN~15 (
// Equation(s):
// \PCregN~15_combout  = (plif_memwbpcsrc_l_1 & ((\PCregN~14_combout  & (plif_memwbporto_l_9)) # (!\PCregN~14_combout  & ((plif_memwbjaddr_l_7))))) # (!plif_memwbpcsrc_l_1 & (((\PCregN~14_combout ))))

	.dataa(plif_memwbporto_l_9),
	.datab(plif_memwbpcsrc_l_1),
	.datac(plif_memwbjaddr_l_7),
	.datad(\PCregN~14_combout ),
	.cin(gnd),
	.combout(\PCregN~15_combout ),
	.cout());
// synopsys translate_off
defparam \PCregN~15 .lut_mask = 16'hBBC0;
defparam \PCregN~15 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y33_N4
cycloneive_lcell_comb \PCregN~16 (
// Equation(s):
// \PCregN~16_combout  = (plif_memwbpcsrc_l_1 & (((plif_memwbjaddr_l_6) # (\pcsrc~0_combout )))) # (!plif_memwbpcsrc_l_1 & (pcifrtnaddr_8 & ((!\pcsrc~0_combout ))))

	.dataa(pcifrtnaddr_8),
	.datab(plif_memwbpcsrc_l_1),
	.datac(plif_memwbjaddr_l_6),
	.datad(pcsrc),
	.cin(gnd),
	.combout(\PCregN~16_combout ),
	.cout());
// synopsys translate_off
defparam \PCregN~16 .lut_mask = 16'hCCE2;
defparam \PCregN~16 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y32_N14
cycloneive_lcell_comb \Add1~12 (
// Equation(s):
// \Add1~12_combout  = ((plif_memwbrtnaddr_l_8 $ (plif_memwbextimm_l_6 $ (!\Add1~11 )))) # (GND)
// \Add1~13  = CARRY((plif_memwbrtnaddr_l_8 & ((plif_memwbextimm_l_6) # (!\Add1~11 ))) # (!plif_memwbrtnaddr_l_8 & (plif_memwbextimm_l_6 & !\Add1~11 )))

	.dataa(plif_memwbrtnaddr_l_8),
	.datab(plif_memwbextimm_l_6),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add1~11 ),
	.combout(\Add1~12_combout ),
	.cout(\Add1~13 ));
// synopsys translate_off
defparam \Add1~12 .lut_mask = 16'h698E;
defparam \Add1~12 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X54_Y33_N30
cycloneive_lcell_comb \PCregN~17 (
// Equation(s):
// \PCregN~17_combout  = (\PCregN~16_combout  & ((plif_memwbporto_l_8) # ((!\pcsrc~0_combout )))) # (!\PCregN~16_combout  & (((\pcsrc~0_combout  & \Add1~12_combout ))))

	.dataa(\PCregN~16_combout ),
	.datab(plif_memwbporto_l_8),
	.datac(pcsrc),
	.datad(\Add1~12_combout ),
	.cin(gnd),
	.combout(\PCregN~17_combout ),
	.cout());
// synopsys translate_off
defparam \PCregN~17 .lut_mask = 16'hDA8A;
defparam \PCregN~17 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y32_N18
cycloneive_lcell_comb \Add1~16 (
// Equation(s):
// \Add1~16_combout  = ((plif_memwbrtnaddr_l_10 $ (plif_memwbextimm_l_8 $ (!\Add1~15 )))) # (GND)
// \Add1~17  = CARRY((plif_memwbrtnaddr_l_10 & ((plif_memwbextimm_l_8) # (!\Add1~15 ))) # (!plif_memwbrtnaddr_l_10 & (plif_memwbextimm_l_8 & !\Add1~15 )))

	.dataa(plif_memwbrtnaddr_l_10),
	.datab(plif_memwbextimm_l_8),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add1~15 ),
	.combout(\Add1~16_combout ),
	.cout(\Add1~17 ));
// synopsys translate_off
defparam \Add1~16 .lut_mask = 16'h698E;
defparam \Add1~16 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X56_Y32_N20
cycloneive_lcell_comb \Add1~18 (
// Equation(s):
// \Add1~18_combout  = (plif_memwbextimm_l_9 & ((plif_memwbrtnaddr_l_11 & (\Add1~17  & VCC)) # (!plif_memwbrtnaddr_l_11 & (!\Add1~17 )))) # (!plif_memwbextimm_l_9 & ((plif_memwbrtnaddr_l_11 & (!\Add1~17 )) # (!plif_memwbrtnaddr_l_11 & ((\Add1~17 ) # 
// (GND)))))
// \Add1~19  = CARRY((plif_memwbextimm_l_9 & (!plif_memwbrtnaddr_l_11 & !\Add1~17 )) # (!plif_memwbextimm_l_9 & ((!\Add1~17 ) # (!plif_memwbrtnaddr_l_11))))

	.dataa(plif_memwbextimm_l_9),
	.datab(plif_memwbrtnaddr_l_11),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add1~17 ),
	.combout(\Add1~18_combout ),
	.cout(\Add1~19 ));
// synopsys translate_off
defparam \Add1~18 .lut_mask = 16'h9617;
defparam \Add1~18 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X53_Y33_N0
cycloneive_lcell_comb \PCregN~18 (
// Equation(s):
// \PCregN~18_combout  = (\pcsrc~0_combout  & ((\Add1~18_combout ) # ((plif_memwbpcsrc_l_1)))) # (!\pcsrc~0_combout  & (((!plif_memwbpcsrc_l_1 & pcifrtnaddr_11))))

	.dataa(pcsrc),
	.datab(\Add1~18_combout ),
	.datac(plif_memwbpcsrc_l_1),
	.datad(pcifrtnaddr_11),
	.cin(gnd),
	.combout(\PCregN~18_combout ),
	.cout());
// synopsys translate_off
defparam \PCregN~18 .lut_mask = 16'hADA8;
defparam \PCregN~18 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y34_N14
cycloneive_lcell_comb \PCregN~19 (
// Equation(s):
// \PCregN~19_combout  = (\PCregN~18_combout  & (((plif_memwbporto_l_11) # (!plif_memwbpcsrc_l_1)))) # (!\PCregN~18_combout  & (plif_memwbjaddr_l_9 & ((plif_memwbpcsrc_l_1))))

	.dataa(plif_memwbjaddr_l_9),
	.datab(plif_memwbporto_l_11),
	.datac(\PCregN~18_combout ),
	.datad(plif_memwbpcsrc_l_1),
	.cin(gnd),
	.combout(\PCregN~19_combout ),
	.cout());
// synopsys translate_off
defparam \PCregN~19 .lut_mask = 16'hCAF0;
defparam \PCregN~19 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y34_N4
cycloneive_lcell_comb \PCregN~20 (
// Equation(s):
// \PCregN~20_combout  = (\pcsrc~0_combout  & (plif_memwbpcsrc_l_1)) # (!\pcsrc~0_combout  & ((plif_memwbpcsrc_l_1 & (plif_memwbjaddr_l_8)) # (!plif_memwbpcsrc_l_1 & ((pcifrtnaddr_10)))))

	.dataa(pcsrc),
	.datab(plif_memwbpcsrc_l_1),
	.datac(plif_memwbjaddr_l_8),
	.datad(pcifrtnaddr_10),
	.cin(gnd),
	.combout(\PCregN~20_combout ),
	.cout());
// synopsys translate_off
defparam \PCregN~20 .lut_mask = 16'hD9C8;
defparam \PCregN~20 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y34_N0
cycloneive_lcell_comb \PCregN~21 (
// Equation(s):
// \PCregN~21_combout  = (\pcsrc~0_combout  & ((\PCregN~20_combout  & (plif_memwbporto_l_10)) # (!\PCregN~20_combout  & ((\Add1~16_combout ))))) # (!\pcsrc~0_combout  & (((\PCregN~20_combout ))))

	.dataa(plif_memwbporto_l_10),
	.datab(pcsrc),
	.datac(\Add1~16_combout ),
	.datad(\PCregN~20_combout ),
	.cin(gnd),
	.combout(\PCregN~21_combout ),
	.cout());
// synopsys translate_off
defparam \PCregN~21 .lut_mask = 16'hBBC0;
defparam \PCregN~21 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y32_N22
cycloneive_lcell_comb \Add1~20 (
// Equation(s):
// \Add1~20_combout  = ((plif_memwbrtnaddr_l_12 $ (plif_memwbextimm_l_10 $ (!\Add1~19 )))) # (GND)
// \Add1~21  = CARRY((plif_memwbrtnaddr_l_12 & ((plif_memwbextimm_l_10) # (!\Add1~19 ))) # (!plif_memwbrtnaddr_l_12 & (plif_memwbextimm_l_10 & !\Add1~19 )))

	.dataa(plif_memwbrtnaddr_l_12),
	.datab(plif_memwbextimm_l_10),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add1~19 ),
	.combout(\Add1~20_combout ),
	.cout(\Add1~21 ));
// synopsys translate_off
defparam \Add1~20 .lut_mask = 16'h698E;
defparam \Add1~20 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X56_Y32_N24
cycloneive_lcell_comb \Add1~22 (
// Equation(s):
// \Add1~22_combout  = (plif_memwbextimm_l_11 & ((plif_memwbrtnaddr_l_13 & (\Add1~21  & VCC)) # (!plif_memwbrtnaddr_l_13 & (!\Add1~21 )))) # (!plif_memwbextimm_l_11 & ((plif_memwbrtnaddr_l_13 & (!\Add1~21 )) # (!plif_memwbrtnaddr_l_13 & ((\Add1~21 ) # 
// (GND)))))
// \Add1~23  = CARRY((plif_memwbextimm_l_11 & (!plif_memwbrtnaddr_l_13 & !\Add1~21 )) # (!plif_memwbextimm_l_11 & ((!\Add1~21 ) # (!plif_memwbrtnaddr_l_13))))

	.dataa(plif_memwbextimm_l_11),
	.datab(plif_memwbrtnaddr_l_13),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add1~21 ),
	.combout(\Add1~22_combout ),
	.cout(\Add1~23 ));
// synopsys translate_off
defparam \Add1~22 .lut_mask = 16'h9617;
defparam \Add1~22 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X54_Y32_N12
cycloneive_lcell_comb \PCregN~22 (
// Equation(s):
// \PCregN~22_combout  = (plif_memwbpcsrc_l_1 & (((\pcsrc~0_combout )))) # (!plif_memwbpcsrc_l_1 & ((\pcsrc~0_combout  & ((\Add1~22_combout ))) # (!\pcsrc~0_combout  & (pcifrtnaddr_13))))

	.dataa(pcifrtnaddr_13),
	.datab(plif_memwbpcsrc_l_1),
	.datac(\Add1~22_combout ),
	.datad(pcsrc),
	.cin(gnd),
	.combout(\PCregN~22_combout ),
	.cout());
// synopsys translate_off
defparam \PCregN~22 .lut_mask = 16'hFC22;
defparam \PCregN~22 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y32_N8
cycloneive_lcell_comb \PCregN~23 (
// Equation(s):
// \PCregN~23_combout  = (plif_memwbpcsrc_l_1 & ((\PCregN~22_combout  & ((plif_memwbporto_l_13))) # (!\PCregN~22_combout  & (plif_memwbjaddr_l_11)))) # (!plif_memwbpcsrc_l_1 & (((\PCregN~22_combout ))))

	.dataa(plif_memwbjaddr_l_11),
	.datab(plif_memwbpcsrc_l_1),
	.datac(plif_memwbporto_l_13),
	.datad(\PCregN~22_combout ),
	.cin(gnd),
	.combout(\PCregN~23_combout ),
	.cout());
// synopsys translate_off
defparam \PCregN~23 .lut_mask = 16'hF388;
defparam \PCregN~23 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X50_Y33_N14
cycloneive_lcell_comb \PCregN~24 (
// Equation(s):
// \PCregN~24_combout  = (plif_memwbpcsrc_l_1 & (((plif_memwbjaddr_l_10) # (\pcsrc~0_combout )))) # (!plif_memwbpcsrc_l_1 & (pcifrtnaddr_12 & ((!\pcsrc~0_combout ))))

	.dataa(pcifrtnaddr_12),
	.datab(plif_memwbpcsrc_l_1),
	.datac(plif_memwbjaddr_l_10),
	.datad(pcsrc),
	.cin(gnd),
	.combout(\PCregN~24_combout ),
	.cout());
// synopsys translate_off
defparam \PCregN~24 .lut_mask = 16'hCCE2;
defparam \PCregN~24 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y32_N18
cycloneive_lcell_comb \PCregN~25 (
// Equation(s):
// \PCregN~25_combout  = (\pcsrc~0_combout  & ((\PCregN~24_combout  & (plif_memwbporto_l_12)) # (!\PCregN~24_combout  & ((\Add1~20_combout ))))) # (!\pcsrc~0_combout  & (((\PCregN~24_combout ))))

	.dataa(plif_memwbporto_l_12),
	.datab(pcsrc),
	.datac(\PCregN~24_combout ),
	.datad(\Add1~20_combout ),
	.cin(gnd),
	.combout(\PCregN~25_combout ),
	.cout());
// synopsys translate_off
defparam \PCregN~25 .lut_mask = 16'hBCB0;
defparam \PCregN~25 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y32_N28
cycloneive_lcell_comb \Add1~26 (
// Equation(s):
// \Add1~26_combout  = (plif_memwbrtnaddr_l_15 & ((plif_memwbextimm_l_13 & (\Add1~25  & VCC)) # (!plif_memwbextimm_l_13 & (!\Add1~25 )))) # (!plif_memwbrtnaddr_l_15 & ((plif_memwbextimm_l_13 & (!\Add1~25 )) # (!plif_memwbextimm_l_13 & ((\Add1~25 ) # 
// (GND)))))
// \Add1~27  = CARRY((plif_memwbrtnaddr_l_15 & (!plif_memwbextimm_l_13 & !\Add1~25 )) # (!plif_memwbrtnaddr_l_15 & ((!\Add1~25 ) # (!plif_memwbextimm_l_13))))

	.dataa(plif_memwbrtnaddr_l_15),
	.datab(plif_memwbextimm_l_13),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add1~25 ),
	.combout(\Add1~26_combout ),
	.cout(\Add1~27 ));
// synopsys translate_off
defparam \Add1~26 .lut_mask = 16'h9617;
defparam \Add1~26 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X52_Y34_N10
cycloneive_lcell_comb \PCregN~26 (
// Equation(s):
// \PCregN~26_combout  = (plif_memwbpcsrc_l_1 & (((\pcsrc~0_combout )))) # (!plif_memwbpcsrc_l_1 & ((\pcsrc~0_combout  & ((\Add1~26_combout ))) # (!\pcsrc~0_combout  & (pcifrtnaddr_15))))

	.dataa(pcifrtnaddr_15),
	.datab(plif_memwbpcsrc_l_1),
	.datac(pcsrc),
	.datad(\Add1~26_combout ),
	.cin(gnd),
	.combout(\PCregN~26_combout ),
	.cout());
// synopsys translate_off
defparam \PCregN~26 .lut_mask = 16'hF2C2;
defparam \PCregN~26 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X52_Y34_N4
cycloneive_lcell_comb \PCregN~27 (
// Equation(s):
// \PCregN~27_combout  = (plif_memwbpcsrc_l_1 & ((\PCregN~26_combout  & ((plif_memwbporto_l_15))) # (!\PCregN~26_combout  & (plif_memwbjaddr_l_13)))) # (!plif_memwbpcsrc_l_1 & (((\PCregN~26_combout ))))

	.dataa(plif_memwbjaddr_l_13),
	.datab(plif_memwbpcsrc_l_1),
	.datac(plif_memwbporto_l_15),
	.datad(\PCregN~26_combout ),
	.cin(gnd),
	.combout(\PCregN~27_combout ),
	.cout());
// synopsys translate_off
defparam \PCregN~27 .lut_mask = 16'hF388;
defparam \PCregN~27 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X50_Y33_N2
cycloneive_lcell_comb \PCregN~28 (
// Equation(s):
// \PCregN~28_combout  = (plif_memwbpcsrc_l_1 & (((plif_memwbjaddr_l_12) # (\pcsrc~0_combout )))) # (!plif_memwbpcsrc_l_1 & (pcifrtnaddr_14 & ((!\pcsrc~0_combout ))))

	.dataa(pcifrtnaddr_14),
	.datab(plif_memwbpcsrc_l_1),
	.datac(plif_memwbjaddr_l_12),
	.datad(pcsrc),
	.cin(gnd),
	.combout(\PCregN~28_combout ),
	.cout());
// synopsys translate_off
defparam \PCregN~28 .lut_mask = 16'hCCE2;
defparam \PCregN~28 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y34_N28
cycloneive_lcell_comb \PCregN~29 (
// Equation(s):
// \PCregN~29_combout  = (\pcsrc~0_combout  & ((\PCregN~28_combout  & ((plif_memwbporto_l_14))) # (!\PCregN~28_combout  & (\Add1~24_combout )))) # (!\pcsrc~0_combout  & (((\PCregN~28_combout ))))

	.dataa(\Add1~24_combout ),
	.datab(plif_memwbporto_l_14),
	.datac(pcsrc),
	.datad(\PCregN~28_combout ),
	.cin(gnd),
	.combout(\PCregN~29_combout ),
	.cout());
// synopsys translate_off
defparam \PCregN~29 .lut_mask = 16'hCFA0;
defparam \PCregN~29 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X52_Y34_N30
cycloneive_lcell_comb \PCreg[14]~feeder (
// Equation(s):
// \PCreg[14]~feeder_combout  = \PCregN~29_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(\PCregN~29_combout ),
	.cin(gnd),
	.combout(\PCreg[14]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \PCreg[14]~feeder .lut_mask = 16'hFF00;
defparam \PCreg[14]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y32_N30
cycloneive_lcell_comb \Add1~28 (
// Equation(s):
// \Add1~28_combout  = ((plif_memwbextimm_l_14 $ (plif_memwbrtnaddr_l_16 $ (!\Add1~27 )))) # (GND)
// \Add1~29  = CARRY((plif_memwbextimm_l_14 & ((plif_memwbrtnaddr_l_16) # (!\Add1~27 ))) # (!plif_memwbextimm_l_14 & (plif_memwbrtnaddr_l_16 & !\Add1~27 )))

	.dataa(plif_memwbextimm_l_14),
	.datab(plif_memwbrtnaddr_l_16),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add1~27 ),
	.combout(\Add1~28_combout ),
	.cout(\Add1~29 ));
// synopsys translate_off
defparam \Add1~28 .lut_mask = 16'h698E;
defparam \Add1~28 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X56_Y31_N0
cycloneive_lcell_comb \Add1~30 (
// Equation(s):
// \Add1~30_combout  = (plif_memwbextimm_l_15 & ((plif_memwbrtnaddr_l_17 & (\Add1~29  & VCC)) # (!plif_memwbrtnaddr_l_17 & (!\Add1~29 )))) # (!plif_memwbextimm_l_15 & ((plif_memwbrtnaddr_l_17 & (!\Add1~29 )) # (!plif_memwbrtnaddr_l_17 & ((\Add1~29 ) # 
// (GND)))))
// \Add1~31  = CARRY((plif_memwbextimm_l_15 & (!plif_memwbrtnaddr_l_17 & !\Add1~29 )) # (!plif_memwbextimm_l_15 & ((!\Add1~29 ) # (!plif_memwbrtnaddr_l_17))))

	.dataa(plif_memwbextimm_l_15),
	.datab(plif_memwbrtnaddr_l_17),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add1~29 ),
	.combout(\Add1~30_combout ),
	.cout(\Add1~31 ));
// synopsys translate_off
defparam \Add1~30 .lut_mask = 16'h9617;
defparam \Add1~30 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X50_Y34_N30
cycloneive_lcell_comb \PCregN~30 (
// Equation(s):
// \PCregN~30_combout  = (plif_memwbpcsrc_l_1 & (\pcsrc~0_combout )) # (!plif_memwbpcsrc_l_1 & ((\pcsrc~0_combout  & (\Add1~30_combout )) # (!\pcsrc~0_combout  & ((pcifrtnaddr_17)))))

	.dataa(plif_memwbpcsrc_l_1),
	.datab(pcsrc),
	.datac(\Add1~30_combout ),
	.datad(pcifrtnaddr_17),
	.cin(gnd),
	.combout(\PCregN~30_combout ),
	.cout());
// synopsys translate_off
defparam \PCregN~30 .lut_mask = 16'hD9C8;
defparam \PCregN~30 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X50_Y34_N4
cycloneive_lcell_comb \PCregN~31 (
// Equation(s):
// \PCregN~31_combout  = (plif_memwbpcsrc_l_1 & ((\PCregN~30_combout  & ((plif_memwbporto_l_17))) # (!\PCregN~30_combout  & (plif_memwbjaddr_l_15)))) # (!plif_memwbpcsrc_l_1 & (((\PCregN~30_combout ))))

	.dataa(plif_memwbpcsrc_l_1),
	.datab(plif_memwbjaddr_l_15),
	.datac(\PCregN~30_combout ),
	.datad(plif_memwbporto_l_17),
	.cin(gnd),
	.combout(\PCregN~31_combout ),
	.cout());
// synopsys translate_off
defparam \PCregN~31 .lut_mask = 16'hF858;
defparam \PCregN~31 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X50_Y33_N0
cycloneive_lcell_comb \PCregN~32 (
// Equation(s):
// \PCregN~32_combout  = (plif_memwbpcsrc_l_1 & (((plif_memwbjaddr_l_14) # (\pcsrc~0_combout )))) # (!plif_memwbpcsrc_l_1 & (pcifrtnaddr_16 & ((!\pcsrc~0_combout ))))

	.dataa(pcifrtnaddr_16),
	.datab(plif_memwbpcsrc_l_1),
	.datac(plif_memwbjaddr_l_14),
	.datad(pcsrc),
	.cin(gnd),
	.combout(\PCregN~32_combout ),
	.cout());
// synopsys translate_off
defparam \PCregN~32 .lut_mask = 16'hCCE2;
defparam \PCregN~32 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X50_Y34_N0
cycloneive_lcell_comb \PCregN~33 (
// Equation(s):
// \PCregN~33_combout  = (\pcsrc~0_combout  & ((\PCregN~32_combout  & (plif_memwbporto_l_16)) # (!\PCregN~32_combout  & ((\Add1~28_combout ))))) # (!\pcsrc~0_combout  & (((\PCregN~32_combout ))))

	.dataa(plif_memwbporto_l_16),
	.datab(\Add1~28_combout ),
	.datac(pcsrc),
	.datad(\PCregN~32_combout ),
	.cin(gnd),
	.combout(\PCregN~33_combout ),
	.cout());
// synopsys translate_off
defparam \PCregN~33 .lut_mask = 16'hAFC0;
defparam \PCregN~33 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y31_N2
cycloneive_lcell_comb \Add1~32 (
// Equation(s):
// \Add1~32_combout  = ((plif_memwbrtnaddr_l_18 $ (plif_memwbextimm_l_16 $ (!\Add1~31 )))) # (GND)
// \Add1~33  = CARRY((plif_memwbrtnaddr_l_18 & ((plif_memwbextimm_l_16) # (!\Add1~31 ))) # (!plif_memwbrtnaddr_l_18 & (plif_memwbextimm_l_16 & !\Add1~31 )))

	.dataa(plif_memwbrtnaddr_l_18),
	.datab(plif_memwbextimm_l_16),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add1~31 ),
	.combout(\Add1~32_combout ),
	.cout(\Add1~33 ));
// synopsys translate_off
defparam \Add1~32 .lut_mask = 16'h698E;
defparam \Add1~32 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X56_Y31_N4
cycloneive_lcell_comb \Add1~34 (
// Equation(s):
// \Add1~34_combout  = (plif_memwbrtnaddr_l_19 & ((plif_memwbextimm_l_17 & (\Add1~33  & VCC)) # (!plif_memwbextimm_l_17 & (!\Add1~33 )))) # (!plif_memwbrtnaddr_l_19 & ((plif_memwbextimm_l_17 & (!\Add1~33 )) # (!plif_memwbextimm_l_17 & ((\Add1~33 ) # 
// (GND)))))
// \Add1~35  = CARRY((plif_memwbrtnaddr_l_19 & (!plif_memwbextimm_l_17 & !\Add1~33 )) # (!plif_memwbrtnaddr_l_19 & ((!\Add1~33 ) # (!plif_memwbextimm_l_17))))

	.dataa(plif_memwbrtnaddr_l_19),
	.datab(plif_memwbextimm_l_17),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add1~33 ),
	.combout(\Add1~34_combout ),
	.cout(\Add1~35 ));
// synopsys translate_off
defparam \Add1~34 .lut_mask = 16'h9617;
defparam \Add1~34 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X54_Y33_N28
cycloneive_lcell_comb \PCregN~34 (
// Equation(s):
// \PCregN~34_combout  = (plif_memwbpcsrc_l_1 & (((\pcsrc~0_combout )))) # (!plif_memwbpcsrc_l_1 & ((\pcsrc~0_combout  & ((\Add1~34_combout ))) # (!\pcsrc~0_combout  & (pcifrtnaddr_19))))

	.dataa(pcifrtnaddr_19),
	.datab(plif_memwbpcsrc_l_1),
	.datac(pcsrc),
	.datad(\Add1~34_combout ),
	.cin(gnd),
	.combout(\PCregN~34_combout ),
	.cout());
// synopsys translate_off
defparam \PCregN~34 .lut_mask = 16'hF2C2;
defparam \PCregN~34 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y33_N0
cycloneive_lcell_comb \PCregN~35 (
// Equation(s):
// \PCregN~35_combout  = (plif_memwbpcsrc_l_1 & ((\PCregN~34_combout  & (plif_memwbporto_l_19)) # (!\PCregN~34_combout  & ((plif_memwbjaddr_l_17))))) # (!plif_memwbpcsrc_l_1 & (((\PCregN~34_combout ))))

	.dataa(plif_memwbporto_l_19),
	.datab(plif_memwbpcsrc_l_1),
	.datac(plif_memwbjaddr_l_17),
	.datad(\PCregN~34_combout ),
	.cin(gnd),
	.combout(\PCregN~35_combout ),
	.cout());
// synopsys translate_off
defparam \PCregN~35 .lut_mask = 16'hBBC0;
defparam \PCregN~35 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y33_N2
cycloneive_lcell_comb \PCregN~36 (
// Equation(s):
// \PCregN~36_combout  = (\pcsrc~0_combout  & (plif_memwbpcsrc_l_1)) # (!\pcsrc~0_combout  & ((plif_memwbpcsrc_l_1 & (plif_memwbjaddr_l_16)) # (!plif_memwbpcsrc_l_1 & ((pcifrtnaddr_18)))))

	.dataa(pcsrc),
	.datab(plif_memwbpcsrc_l_1),
	.datac(plif_memwbjaddr_l_16),
	.datad(pcifrtnaddr_18),
	.cin(gnd),
	.combout(\PCregN~36_combout ),
	.cout());
// synopsys translate_off
defparam \PCregN~36 .lut_mask = 16'hD9C8;
defparam \PCregN~36 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y33_N4
cycloneive_lcell_comb \PCregN~37 (
// Equation(s):
// \PCregN~37_combout  = (\PCregN~36_combout  & ((plif_memwbporto_l_18) # ((!\pcsrc~0_combout )))) # (!\PCregN~36_combout  & (((\pcsrc~0_combout  & \Add1~32_combout ))))

	.dataa(\PCregN~36_combout ),
	.datab(plif_memwbporto_l_18),
	.datac(pcsrc),
	.datad(\Add1~32_combout ),
	.cin(gnd),
	.combout(\PCregN~37_combout ),
	.cout());
// synopsys translate_off
defparam \PCregN~37 .lut_mask = 16'hDA8A;
defparam \PCregN~37 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y31_N6
cycloneive_lcell_comb \Add1~36 (
// Equation(s):
// \Add1~36_combout  = ((plif_memwbextimm_l_18 $ (plif_memwbrtnaddr_l_20 $ (!\Add1~35 )))) # (GND)
// \Add1~37  = CARRY((plif_memwbextimm_l_18 & ((plif_memwbrtnaddr_l_20) # (!\Add1~35 ))) # (!plif_memwbextimm_l_18 & (plif_memwbrtnaddr_l_20 & !\Add1~35 )))

	.dataa(plif_memwbextimm_l_18),
	.datab(plif_memwbrtnaddr_l_20),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add1~35 ),
	.combout(\Add1~36_combout ),
	.cout(\Add1~37 ));
// synopsys translate_off
defparam \Add1~36 .lut_mask = 16'h698E;
defparam \Add1~36 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X56_Y31_N8
cycloneive_lcell_comb \Add1~38 (
// Equation(s):
// \Add1~38_combout  = (plif_memwbrtnaddr_l_21 & ((plif_memwbextimm_l_19 & (\Add1~37  & VCC)) # (!plif_memwbextimm_l_19 & (!\Add1~37 )))) # (!plif_memwbrtnaddr_l_21 & ((plif_memwbextimm_l_19 & (!\Add1~37 )) # (!plif_memwbextimm_l_19 & ((\Add1~37 ) # 
// (GND)))))
// \Add1~39  = CARRY((plif_memwbrtnaddr_l_21 & (!plif_memwbextimm_l_19 & !\Add1~37 )) # (!plif_memwbrtnaddr_l_21 & ((!\Add1~37 ) # (!plif_memwbextimm_l_19))))

	.dataa(plif_memwbrtnaddr_l_21),
	.datab(plif_memwbextimm_l_19),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add1~37 ),
	.combout(\Add1~38_combout ),
	.cout(\Add1~39 ));
// synopsys translate_off
defparam \Add1~38 .lut_mask = 16'h9617;
defparam \Add1~38 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X53_Y31_N4
cycloneive_lcell_comb \PCregN~38 (
// Equation(s):
// \PCregN~38_combout  = (plif_memwbpcsrc_l_1 & (\pcsrc~0_combout )) # (!plif_memwbpcsrc_l_1 & ((\pcsrc~0_combout  & ((\Add1~38_combout ))) # (!\pcsrc~0_combout  & (pcifrtnaddr_21))))

	.dataa(plif_memwbpcsrc_l_1),
	.datab(pcsrc),
	.datac(pcifrtnaddr_21),
	.datad(\Add1~38_combout ),
	.cin(gnd),
	.combout(\PCregN~38_combout ),
	.cout());
// synopsys translate_off
defparam \PCregN~38 .lut_mask = 16'hDC98;
defparam \PCregN~38 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X52_Y34_N16
cycloneive_lcell_comb \PCregN~39 (
// Equation(s):
// \PCregN~39_combout  = (\PCregN~38_combout  & (((plif_memwbporto_l_21) # (!plif_memwbpcsrc_l_1)))) # (!\PCregN~38_combout  & (plif_memwbjaddr_l_19 & ((plif_memwbpcsrc_l_1))))

	.dataa(\PCregN~38_combout ),
	.datab(plif_memwbjaddr_l_19),
	.datac(plif_memwbporto_l_21),
	.datad(plif_memwbpcsrc_l_1),
	.cin(gnd),
	.combout(\PCregN~39_combout ),
	.cout());
// synopsys translate_off
defparam \PCregN~39 .lut_mask = 16'hE4AA;
defparam \PCregN~39 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y33_N14
cycloneive_lcell_comb \PCregN~40 (
// Equation(s):
// \PCregN~40_combout  = (\pcsrc~0_combout  & (plif_memwbpcsrc_l_1)) # (!\pcsrc~0_combout  & ((plif_memwbpcsrc_l_1 & (plif_memwbjaddr_l_18)) # (!plif_memwbpcsrc_l_1 & ((pcifrtnaddr_20)))))

	.dataa(pcsrc),
	.datab(plif_memwbpcsrc_l_1),
	.datac(plif_memwbjaddr_l_18),
	.datad(pcifrtnaddr_20),
	.cin(gnd),
	.combout(\PCregN~40_combout ),
	.cout());
// synopsys translate_off
defparam \PCregN~40 .lut_mask = 16'hD9C8;
defparam \PCregN~40 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y34_N12
cycloneive_lcell_comb \PCregN~41 (
// Equation(s):
// \PCregN~41_combout  = (\pcsrc~0_combout  & ((\PCregN~40_combout  & (plif_memwbporto_l_20)) # (!\PCregN~40_combout  & ((\Add1~36_combout ))))) # (!\pcsrc~0_combout  & (((\PCregN~40_combout ))))

	.dataa(pcsrc),
	.datab(plif_memwbporto_l_20),
	.datac(\PCregN~40_combout ),
	.datad(\Add1~36_combout ),
	.cin(gnd),
	.combout(\PCregN~41_combout ),
	.cout());
// synopsys translate_off
defparam \PCregN~41 .lut_mask = 16'hDAD0;
defparam \PCregN~41 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y31_N10
cycloneive_lcell_comb \Add1~40 (
// Equation(s):
// \Add1~40_combout  = ((plif_memwbrtnaddr_l_22 $ (plif_memwbextimm_l_20 $ (!\Add1~39 )))) # (GND)
// \Add1~41  = CARRY((plif_memwbrtnaddr_l_22 & ((plif_memwbextimm_l_20) # (!\Add1~39 ))) # (!plif_memwbrtnaddr_l_22 & (plif_memwbextimm_l_20 & !\Add1~39 )))

	.dataa(plif_memwbrtnaddr_l_22),
	.datab(plif_memwbextimm_l_20),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add1~39 ),
	.combout(\Add1~40_combout ),
	.cout(\Add1~41 ));
// synopsys translate_off
defparam \Add1~40 .lut_mask = 16'h698E;
defparam \Add1~40 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X56_Y31_N12
cycloneive_lcell_comb \Add1~42 (
// Equation(s):
// \Add1~42_combout  = (plif_memwbrtnaddr_l_23 & ((plif_memwbextimm_l_21 & (\Add1~41  & VCC)) # (!plif_memwbextimm_l_21 & (!\Add1~41 )))) # (!plif_memwbrtnaddr_l_23 & ((plif_memwbextimm_l_21 & (!\Add1~41 )) # (!plif_memwbextimm_l_21 & ((\Add1~41 ) # 
// (GND)))))
// \Add1~43  = CARRY((plif_memwbrtnaddr_l_23 & (!plif_memwbextimm_l_21 & !\Add1~41 )) # (!plif_memwbrtnaddr_l_23 & ((!\Add1~41 ) # (!plif_memwbextimm_l_21))))

	.dataa(plif_memwbrtnaddr_l_23),
	.datab(plif_memwbextimm_l_21),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add1~41 ),
	.combout(\Add1~42_combout ),
	.cout(\Add1~43 ));
// synopsys translate_off
defparam \Add1~42 .lut_mask = 16'h9617;
defparam \Add1~42 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X52_Y31_N0
cycloneive_lcell_comb \PCregN~42 (
// Equation(s):
// \PCregN~42_combout  = (\pcsrc~0_combout  & (((\Add1~42_combout ) # (plif_memwbpcsrc_l_1)))) # (!\pcsrc~0_combout  & (pcifrtnaddr_23 & ((!plif_memwbpcsrc_l_1))))

	.dataa(pcifrtnaddr_23),
	.datab(\Add1~42_combout ),
	.datac(pcsrc),
	.datad(plif_memwbpcsrc_l_1),
	.cin(gnd),
	.combout(\PCregN~42_combout ),
	.cout());
// synopsys translate_off
defparam \PCregN~42 .lut_mask = 16'hF0CA;
defparam \PCregN~42 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X52_Y32_N30
cycloneive_lcell_comb \PCregN~43 (
// Equation(s):
// \PCregN~43_combout  = (plif_memwbpcsrc_l_1 & ((\PCregN~42_combout  & (plif_memwbporto_l_23)) # (!\PCregN~42_combout  & ((plif_memwbjaddr_l_21))))) # (!plif_memwbpcsrc_l_1 & (((\PCregN~42_combout ))))

	.dataa(plif_memwbporto_l_23),
	.datab(plif_memwbpcsrc_l_1),
	.datac(plif_memwbjaddr_l_21),
	.datad(\PCregN~42_combout ),
	.cin(gnd),
	.combout(\PCregN~43_combout ),
	.cout());
// synopsys translate_off
defparam \PCregN~43 .lut_mask = 16'hBBC0;
defparam \PCregN~43 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y33_N4
cycloneive_lcell_comb \PCregN~44 (
// Equation(s):
// \PCregN~44_combout  = (\pcsrc~0_combout  & (plif_memwbpcsrc_l_1)) # (!\pcsrc~0_combout  & ((plif_memwbpcsrc_l_1 & (plif_memwbjaddr_l_20)) # (!plif_memwbpcsrc_l_1 & ((pcifrtnaddr_22)))))

	.dataa(pcsrc),
	.datab(plif_memwbpcsrc_l_1),
	.datac(plif_memwbjaddr_l_20),
	.datad(pcifrtnaddr_22),
	.cin(gnd),
	.combout(\PCregN~44_combout ),
	.cout());
// synopsys translate_off
defparam \PCregN~44 .lut_mask = 16'hD9C8;
defparam \PCregN~44 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X52_Y34_N14
cycloneive_lcell_comb \PCregN~45 (
// Equation(s):
// \PCregN~45_combout  = (\pcsrc~0_combout  & ((\PCregN~44_combout  & (plif_memwbporto_l_22)) # (!\PCregN~44_combout  & ((\Add1~40_combout ))))) # (!\pcsrc~0_combout  & (((\PCregN~44_combout ))))

	.dataa(plif_memwbporto_l_22),
	.datab(pcsrc),
	.datac(\PCregN~44_combout ),
	.datad(\Add1~40_combout ),
	.cin(gnd),
	.combout(\PCregN~45_combout ),
	.cout());
// synopsys translate_off
defparam \PCregN~45 .lut_mask = 16'hBCB0;
defparam \PCregN~45 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y31_N14
cycloneive_lcell_comb \Add1~44 (
// Equation(s):
// \Add1~44_combout  = ((plif_memwbextimm_l_22 $ (plif_memwbrtnaddr_l_24 $ (!\Add1~43 )))) # (GND)
// \Add1~45  = CARRY((plif_memwbextimm_l_22 & ((plif_memwbrtnaddr_l_24) # (!\Add1~43 ))) # (!plif_memwbextimm_l_22 & (plif_memwbrtnaddr_l_24 & !\Add1~43 )))

	.dataa(plif_memwbextimm_l_22),
	.datab(plif_memwbrtnaddr_l_24),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add1~43 ),
	.combout(\Add1~44_combout ),
	.cout(\Add1~45 ));
// synopsys translate_off
defparam \Add1~44 .lut_mask = 16'h698E;
defparam \Add1~44 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X56_Y31_N16
cycloneive_lcell_comb \Add1~46 (
// Equation(s):
// \Add1~46_combout  = (plif_memwbrtnaddr_l_25 & ((plif_memwbextimm_l_23 & (\Add1~45  & VCC)) # (!plif_memwbextimm_l_23 & (!\Add1~45 )))) # (!plif_memwbrtnaddr_l_25 & ((plif_memwbextimm_l_23 & (!\Add1~45 )) # (!plif_memwbextimm_l_23 & ((\Add1~45 ) # 
// (GND)))))
// \Add1~47  = CARRY((plif_memwbrtnaddr_l_25 & (!plif_memwbextimm_l_23 & !\Add1~45 )) # (!plif_memwbrtnaddr_l_25 & ((!\Add1~45 ) # (!plif_memwbextimm_l_23))))

	.dataa(plif_memwbrtnaddr_l_25),
	.datab(plif_memwbextimm_l_23),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add1~45 ),
	.combout(\Add1~46_combout ),
	.cout(\Add1~47 ));
// synopsys translate_off
defparam \Add1~46 .lut_mask = 16'h9617;
defparam \Add1~46 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X52_Y31_N14
cycloneive_lcell_comb \PCregN~46 (
// Equation(s):
// \PCregN~46_combout  = (plif_memwbpcsrc_l_1 & (((\pcsrc~0_combout )))) # (!plif_memwbpcsrc_l_1 & ((\pcsrc~0_combout  & (\Add1~46_combout )) # (!\pcsrc~0_combout  & ((pcifrtnaddr_25)))))

	.dataa(plif_memwbpcsrc_l_1),
	.datab(\Add1~46_combout ),
	.datac(pcsrc),
	.datad(pcifrtnaddr_25),
	.cin(gnd),
	.combout(\PCregN~46_combout ),
	.cout());
// synopsys translate_off
defparam \PCregN~46 .lut_mask = 16'hE5E0;
defparam \PCregN~46 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y35_N18
cycloneive_lcell_comb \PCregN~47 (
// Equation(s):
// \PCregN~47_combout  = (\PCregN~46_combout  & (((plif_memwbporto_l_25) # (!plif_memwbpcsrc_l_1)))) # (!\PCregN~46_combout  & (plif_memwbjaddr_l_23 & ((plif_memwbpcsrc_l_1))))

	.dataa(plif_memwbjaddr_l_23),
	.datab(plif_memwbporto_l_25),
	.datac(\PCregN~46_combout ),
	.datad(plif_memwbpcsrc_l_1),
	.cin(gnd),
	.combout(\PCregN~47_combout ),
	.cout());
// synopsys translate_off
defparam \PCregN~47 .lut_mask = 16'hCAF0;
defparam \PCregN~47 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y33_N18
cycloneive_lcell_comb \PCregN~48 (
// Equation(s):
// \PCregN~48_combout  = (\pcsrc~0_combout  & (plif_memwbpcsrc_l_1)) # (!\pcsrc~0_combout  & ((plif_memwbpcsrc_l_1 & (plif_memwbjaddr_l_22)) # (!plif_memwbpcsrc_l_1 & ((pcifrtnaddr_24)))))

	.dataa(pcsrc),
	.datab(plif_memwbpcsrc_l_1),
	.datac(plif_memwbjaddr_l_22),
	.datad(pcifrtnaddr_24),
	.cin(gnd),
	.combout(\PCregN~48_combout ),
	.cout());
// synopsys translate_off
defparam \PCregN~48 .lut_mask = 16'hD9C8;
defparam \PCregN~48 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y33_N6
cycloneive_lcell_comb \PCregN~49 (
// Equation(s):
// \PCregN~49_combout  = (\pcsrc~0_combout  & ((\PCregN~48_combout  & (plif_memwbporto_l_24)) # (!\PCregN~48_combout  & ((\Add1~44_combout ))))) # (!\pcsrc~0_combout  & (\PCregN~48_combout ))

	.dataa(pcsrc),
	.datab(\PCregN~48_combout ),
	.datac(plif_memwbporto_l_24),
	.datad(\Add1~44_combout ),
	.cin(gnd),
	.combout(\PCregN~49_combout ),
	.cout());
// synopsys translate_off
defparam \PCregN~49 .lut_mask = 16'hE6C4;
defparam \PCregN~49 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y31_N18
cycloneive_lcell_comb \Add1~48 (
// Equation(s):
// \Add1~48_combout  = ((plif_memwbextimm_l_24 $ (plif_memwbrtnaddr_l_26 $ (!\Add1~47 )))) # (GND)
// \Add1~49  = CARRY((plif_memwbextimm_l_24 & ((plif_memwbrtnaddr_l_26) # (!\Add1~47 ))) # (!plif_memwbextimm_l_24 & (plif_memwbrtnaddr_l_26 & !\Add1~47 )))

	.dataa(plif_memwbextimm_l_24),
	.datab(plif_memwbrtnaddr_l_26),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add1~47 ),
	.combout(\Add1~48_combout ),
	.cout(\Add1~49 ));
// synopsys translate_off
defparam \Add1~48 .lut_mask = 16'h698E;
defparam \Add1~48 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X56_Y31_N20
cycloneive_lcell_comb \Add1~50 (
// Equation(s):
// \Add1~50_combout  = (plif_memwbrtnaddr_l_27 & ((plif_memwbextimm_l_25 & (\Add1~49  & VCC)) # (!plif_memwbextimm_l_25 & (!\Add1~49 )))) # (!plif_memwbrtnaddr_l_27 & ((plif_memwbextimm_l_25 & (!\Add1~49 )) # (!plif_memwbextimm_l_25 & ((\Add1~49 ) # 
// (GND)))))
// \Add1~51  = CARRY((plif_memwbrtnaddr_l_27 & (!plif_memwbextimm_l_25 & !\Add1~49 )) # (!plif_memwbrtnaddr_l_27 & ((!\Add1~49 ) # (!plif_memwbextimm_l_25))))

	.dataa(plif_memwbrtnaddr_l_27),
	.datab(plif_memwbextimm_l_25),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add1~49 ),
	.combout(\Add1~50_combout ),
	.cout(\Add1~51 ));
// synopsys translate_off
defparam \Add1~50 .lut_mask = 16'h9617;
defparam \Add1~50 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X53_Y31_N18
cycloneive_lcell_comb \PCregN~50 (
// Equation(s):
// \PCregN~50_combout  = (plif_memwbpcsrc_l_1 & (\pcsrc~0_combout )) # (!plif_memwbpcsrc_l_1 & ((\pcsrc~0_combout  & (\Add1~50_combout )) # (!\pcsrc~0_combout  & ((pcifrtnaddr_27)))))

	.dataa(plif_memwbpcsrc_l_1),
	.datab(pcsrc),
	.datac(\Add1~50_combout ),
	.datad(pcifrtnaddr_27),
	.cin(gnd),
	.combout(\PCregN~50_combout ),
	.cout());
// synopsys translate_off
defparam \PCregN~50 .lut_mask = 16'hD9C8;
defparam \PCregN~50 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y33_N28
cycloneive_lcell_comb \PCregN~51 (
// Equation(s):
// \PCregN~51_combout  = (plif_memwbpcsrc_l_1 & ((\PCregN~50_combout  & ((plif_memwbporto_l_27))) # (!\PCregN~50_combout  & (plif_memwbjaddr_l_25)))) # (!plif_memwbpcsrc_l_1 & (((\PCregN~50_combout ))))

	.dataa(plif_memwbjaddr_l_25),
	.datab(plif_memwbporto_l_27),
	.datac(plif_memwbpcsrc_l_1),
	.datad(\PCregN~50_combout ),
	.cin(gnd),
	.combout(\PCregN~51_combout ),
	.cout());
// synopsys translate_off
defparam \PCregN~51 .lut_mask = 16'hCFA0;
defparam \PCregN~51 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y33_N14
cycloneive_lcell_comb \PCregN~52 (
// Equation(s):
// \PCregN~52_combout  = (\pcsrc~0_combout  & (plif_memwbpcsrc_l_1)) # (!\pcsrc~0_combout  & ((plif_memwbpcsrc_l_1 & (plif_memwbjaddr_l_24)) # (!plif_memwbpcsrc_l_1 & ((pcifrtnaddr_26)))))

	.dataa(pcsrc),
	.datab(plif_memwbpcsrc_l_1),
	.datac(plif_memwbjaddr_l_24),
	.datad(pcifrtnaddr_26),
	.cin(gnd),
	.combout(\PCregN~52_combout ),
	.cout());
// synopsys translate_off
defparam \PCregN~52 .lut_mask = 16'hD9C8;
defparam \PCregN~52 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y33_N12
cycloneive_lcell_comb \PCregN~53 (
// Equation(s):
// \PCregN~53_combout  = (\pcsrc~0_combout  & ((\PCregN~52_combout  & ((plif_memwbporto_l_26))) # (!\PCregN~52_combout  & (\Add1~48_combout )))) # (!\pcsrc~0_combout  & (\PCregN~52_combout ))

	.dataa(pcsrc),
	.datab(\PCregN~52_combout ),
	.datac(\Add1~48_combout ),
	.datad(plif_memwbporto_l_26),
	.cin(gnd),
	.combout(\PCregN~53_combout ),
	.cout());
// synopsys translate_off
defparam \PCregN~53 .lut_mask = 16'hEC64;
defparam \PCregN~53 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y31_N8
cycloneive_lcell_comb \PCregN~54 (
// Equation(s):
// \PCregN~54_combout  = (\pcsrc~0_combout  & ((\Add1~54_combout ) # ((plif_memwbpcsrc_l_1)))) # (!\pcsrc~0_combout  & (((pcifrtnaddr_29 & !plif_memwbpcsrc_l_1))))

	.dataa(\Add1~54_combout ),
	.datab(pcifrtnaddr_29),
	.datac(pcsrc),
	.datad(plif_memwbpcsrc_l_1),
	.cin(gnd),
	.combout(\PCregN~54_combout ),
	.cout());
// synopsys translate_off
defparam \PCregN~54 .lut_mask = 16'hF0AC;
defparam \PCregN~54 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X50_Y34_N6
cycloneive_lcell_comb \PCregN~55 (
// Equation(s):
// \PCregN~55_combout  = (plif_memwbpcsrc_l_1 & ((\PCregN~54_combout  & ((plif_memwbporto_l_29))) # (!\PCregN~54_combout  & (plif_memwbrtnaddr_l_29)))) # (!plif_memwbpcsrc_l_1 & (((\PCregN~54_combout ))))

	.dataa(plif_memwbpcsrc_l_1),
	.datab(plif_memwbrtnaddr_l_29),
	.datac(plif_memwbporto_l_29),
	.datad(\PCregN~54_combout ),
	.cin(gnd),
	.combout(\PCregN~55_combout ),
	.cout());
// synopsys translate_off
defparam \PCregN~55 .lut_mask = 16'hF588;
defparam \PCregN~55 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X52_Y30_N12
cycloneive_lcell_comb \PCregN~56 (
// Equation(s):
// \PCregN~56_combout  = (\pcsrc~0_combout  & (plif_memwbpcsrc_l_1)) # (!\pcsrc~0_combout  & ((plif_memwbpcsrc_l_1 & (plif_memwbrtnaddr_l_28)) # (!plif_memwbpcsrc_l_1 & ((pcifrtnaddr_28)))))

	.dataa(pcsrc),
	.datab(plif_memwbpcsrc_l_1),
	.datac(plif_memwbrtnaddr_l_28),
	.datad(pcifrtnaddr_28),
	.cin(gnd),
	.combout(\PCregN~56_combout ),
	.cout());
// synopsys translate_off
defparam \PCregN~56 .lut_mask = 16'hD9C8;
defparam \PCregN~56 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y31_N22
cycloneive_lcell_comb \Add1~52 (
// Equation(s):
// \Add1~52_combout  = ((plif_memwbrtnaddr_l_28 $ (plif_memwbextimm_l_26 $ (!\Add1~51 )))) # (GND)
// \Add1~53  = CARRY((plif_memwbrtnaddr_l_28 & ((plif_memwbextimm_l_26) # (!\Add1~51 ))) # (!plif_memwbrtnaddr_l_28 & (plif_memwbextimm_l_26 & !\Add1~51 )))

	.dataa(plif_memwbrtnaddr_l_28),
	.datab(plif_memwbextimm_l_26),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add1~51 ),
	.combout(\Add1~52_combout ),
	.cout(\Add1~53 ));
// synopsys translate_off
defparam \Add1~52 .lut_mask = 16'h698E;
defparam \Add1~52 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X50_Y34_N14
cycloneive_lcell_comb \PCregN~57 (
// Equation(s):
// \PCregN~57_combout  = (\pcsrc~0_combout  & ((\PCregN~56_combout  & (plif_memwbporto_l_28)) # (!\PCregN~56_combout  & ((\Add1~52_combout ))))) # (!\pcsrc~0_combout  & (((\PCregN~56_combout ))))

	.dataa(plif_memwbporto_l_28),
	.datab(pcsrc),
	.datac(\PCregN~56_combout ),
	.datad(\Add1~52_combout ),
	.cin(gnd),
	.combout(\PCregN~57_combout ),
	.cout());
// synopsys translate_off
defparam \PCregN~57 .lut_mask = 16'hBCB0;
defparam \PCregN~57 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y31_N26
cycloneive_lcell_comb \Add1~56 (
// Equation(s):
// \Add1~56_combout  = ((plif_memwbextimm_l_28 $ (plif_memwbrtnaddr_l_30 $ (!\Add1~55 )))) # (GND)
// \Add1~57  = CARRY((plif_memwbextimm_l_28 & ((plif_memwbrtnaddr_l_30) # (!\Add1~55 ))) # (!plif_memwbextimm_l_28 & (plif_memwbrtnaddr_l_30 & !\Add1~55 )))

	.dataa(plif_memwbextimm_l_28),
	.datab(plif_memwbrtnaddr_l_30),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add1~55 ),
	.combout(\Add1~56_combout ),
	.cout(\Add1~57 ));
// synopsys translate_off
defparam \Add1~56 .lut_mask = 16'h698E;
defparam \Add1~56 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X56_Y31_N28
cycloneive_lcell_comb \Add1~58 (
// Equation(s):
// \Add1~58_combout  = plif_memwbextimm_l_29 $ (\Add1~57  $ (plif_memwbrtnaddr_l_31))

	.dataa(gnd),
	.datab(plif_memwbextimm_l_29),
	.datac(gnd),
	.datad(plif_memwbrtnaddr_l_31),
	.cin(\Add1~57 ),
	.combout(\Add1~58_combout ),
	.cout());
// synopsys translate_off
defparam \Add1~58 .lut_mask = 16'hC33C;
defparam \Add1~58 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X52_Y30_N18
cycloneive_lcell_comb \PCregN~58 (
// Equation(s):
// \PCregN~58_combout  = (\pcsrc~0_combout  & ((plif_memwbpcsrc_l_1) # ((\Add1~58_combout )))) # (!\pcsrc~0_combout  & (!plif_memwbpcsrc_l_1 & (pcifrtnaddr_31)))

	.dataa(pcsrc),
	.datab(plif_memwbpcsrc_l_1),
	.datac(pcifrtnaddr_31),
	.datad(\Add1~58_combout ),
	.cin(gnd),
	.combout(\PCregN~58_combout ),
	.cout());
// synopsys translate_off
defparam \PCregN~58 .lut_mask = 16'hBA98;
defparam \PCregN~58 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X52_Y34_N20
cycloneive_lcell_comb \PCregN~59 (
// Equation(s):
// \PCregN~59_combout  = (plif_memwbpcsrc_l_1 & ((\PCregN~58_combout  & ((plif_memwbporto_l_31))) # (!\PCregN~58_combout  & (plif_memwbrtnaddr_l_31)))) # (!plif_memwbpcsrc_l_1 & (((\PCregN~58_combout ))))

	.dataa(plif_memwbrtnaddr_l_31),
	.datab(plif_memwbpcsrc_l_1),
	.datac(plif_memwbporto_l_31),
	.datad(\PCregN~58_combout ),
	.cin(gnd),
	.combout(\PCregN~59_combout ),
	.cout());
// synopsys translate_off
defparam \PCregN~59 .lut_mask = 16'hF388;
defparam \PCregN~59 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y42_N2
cycloneive_lcell_comb \PCregN~60 (
// Equation(s):
// \PCregN~60_combout  = (plif_memwbpcsrc_l_1 & ((\pcsrc~0_combout  & ((plif_memwbporto_l_30))) # (!\pcsrc~0_combout  & (plif_memwbrtnaddr_l_30)))) # (!plif_memwbpcsrc_l_1 & (((\pcsrc~0_combout ))))

	.dataa(plif_memwbpcsrc_l_1),
	.datab(plif_memwbrtnaddr_l_30),
	.datac(plif_memwbporto_l_30),
	.datad(pcsrc),
	.cin(gnd),
	.combout(\PCregN~60_combout ),
	.cout());
// synopsys translate_off
defparam \PCregN~60 .lut_mask = 16'hF588;
defparam \PCregN~60 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y34_N26
cycloneive_lcell_comb \PCregN~61 (
// Equation(s):
// \PCregN~61_combout  = (\PCregN~60_combout  & ((plif_memwbpcsrc_l_1) # ((\Add1~56_combout )))) # (!\PCregN~60_combout  & (!plif_memwbpcsrc_l_1 & (pcifrtnaddr_30)))

	.dataa(\PCregN~60_combout ),
	.datab(plif_memwbpcsrc_l_1),
	.datac(pcifrtnaddr_30),
	.datad(\Add1~56_combout ),
	.cin(gnd),
	.combout(\PCregN~61_combout ),
	.cout());
// synopsys translate_off
defparam \PCregN~61 .lut_mask = 16'hBA98;
defparam \PCregN~61 .sum_lutc_input = "datac";
// synopsys translate_on

endmodule

module pipeline_exmem (
	plif_exmemhlt_l,
	plif_exmemporto_l_1,
	plif_exmemdmemWEN_l,
	plif_exmemdmemREN_l,
	plif_exmemporto_l_0,
	plif_exmemporto_l_3,
	plif_exmemporto_l_2,
	plif_exmemporto_l_5,
	plif_exmemporto_l_4,
	plif_exmemporto_l_7,
	plif_exmemporto_l_6,
	plif_exmemporto_l_9,
	plif_exmemporto_l_8,
	plif_exmemporto_l_11,
	plif_exmemporto_l_10,
	plif_exmemporto_l_13,
	plif_exmemporto_l_12,
	plif_exmemporto_l_15,
	plif_exmemporto_l_14,
	plif_exmemporto_l_17,
	plif_exmemporto_l_16,
	plif_exmemporto_l_19,
	plif_exmemporto_l_18,
	plif_exmemporto_l_21,
	plif_exmemporto_l_20,
	plif_exmemporto_l_23,
	plif_exmemporto_l_22,
	plif_exmemporto_l_25,
	plif_exmemporto_l_24,
	plif_exmemporto_l_27,
	plif_exmemporto_l_26,
	plif_exmemporto_l_29,
	plif_exmemporto_l_28,
	plif_exmemporto_l_31,
	plif_exmemporto_l_30,
	plif_idexhlt_l,
	plif_idexpcsrc_l_1,
	plif_idexpcsrc_l_0,
	plif_exmempcsrc_l_1,
	plif_exmempcsrc_l_0,
	exmem_en,
	plif_exmemrdat2_l_0,
	plif_exmemregen_l,
	plif_exmemwsel_l_0,
	plif_exmemwsel_l_1,
	plif_exmemwsel_l_4,
	plif_exmemwsel_l_3,
	plif_exmemwsel_l_2,
	plif_idexextimm_l_29,
	plif_idexextimm_l_28,
	plif_idexextimm_l_27,
	plif_idexextimm_l_26,
	plif_idexextimm_l_25,
	plif_idexextimm_l_24,
	plif_idexextimm_l_23,
	plif_idexextimm_l_22,
	plif_idexextimm_l_21,
	plif_idexextimm_l_20,
	plif_idexextimm_l_19,
	plif_idexextimm_l_18,
	plif_idexextimm_l_17,
	plif_idexextimm_l_16,
	plif_idexextimm_l_15,
	plif_idexextimm_l_14,
	plif_idexextimm_l_13,
	plif_idexextimm_l_12,
	plif_idexextimm_l_11,
	plif_idexextimm_l_10,
	plif_idexextimm_l_9,
	plif_idexextimm_l_8,
	plif_idexextimm_l_7,
	plif_idexextimm_l_6,
	plif_idexextimm_l_5,
	plif_idexextimm_l_0,
	plif_idexextimm_l_1,
	plif_idexextimm_l_2,
	plif_idexextimm_l_3,
	plif_idexextimm_l_4,
	Selector30,
	plif_idexdmemREN_l,
	plif_idexwsel_l_0,
	plif_idexwsel_l_1,
	plif_idexwsel_l_2,
	plif_idexwsel_l_3,
	plif_idexwsel_l_4,
	plif_idexdmemWEN_l,
	Selector31,
	Selector28,
	Selector29,
	Selector26,
	Selector27,
	Selector24,
	Selector25,
	Selector22,
	Selector23,
	Selector20,
	Selector21,
	Selector18,
	Selector19,
	Selector16,
	Selector17,
	Selector14,
	Selector15,
	Selector12,
	Selector13,
	Selector10,
	Selector11,
	Selector8,
	Selector9,
	Selector6,
	Selector7,
	Selector4,
	Selector5,
	Selector2,
	Selector3,
	Selector0,
	Selector1,
	plif_exmemrdat2_l_1,
	plif_exmemrdat2_l_2,
	plif_exmemrdat2_l_3,
	plif_exmemrdat2_l_4,
	plif_exmemrdat2_l_5,
	plif_exmemrdat2_l_6,
	plif_exmemrdat2_l_7,
	plif_exmemrdat2_l_8,
	plif_exmemrdat2_l_9,
	plif_exmemrdat2_l_10,
	plif_exmemrdat2_l_11,
	plif_exmemrdat2_l_12,
	plif_exmemrdat2_l_13,
	plif_exmemrdat2_l_14,
	plif_exmemrdat2_l_15,
	plif_exmemrdat2_l_16,
	plif_exmemrdat2_l_17,
	plif_exmemrdat2_l_18,
	plif_exmemrdat2_l_19,
	plif_exmemrdat2_l_20,
	plif_exmemrdat2_l_21,
	plif_exmemrdat2_l_22,
	plif_exmemrdat2_l_23,
	plif_exmemrdat2_l_24,
	plif_exmemrdat2_l_25,
	plif_exmemrdat2_l_26,
	plif_exmemrdat2_l_27,
	plif_exmemrdat2_l_28,
	plif_exmemrdat2_l_29,
	plif_exmemrdat2_l_30,
	plif_exmemrdat2_l_31,
	plif_idexregen_l,
	plif_exmemregsrc_l_0,
	plif_exmemregsrc_l_1,
	plif_exmemrtnaddr_l_31,
	plif_exmemrtnaddr_l_30,
	plif_exmemrtnaddr_l_29,
	plif_exmemrtnaddr_l_28,
	plif_exmemrtnaddr_l_27,
	plif_exmemrtnaddr_l_26,
	plif_exmemrtnaddr_l_25,
	plif_exmemrtnaddr_l_24,
	plif_exmemrtnaddr_l_23,
	plif_exmemrtnaddr_l_22,
	plif_exmemrtnaddr_l_21,
	plif_exmemrtnaddr_l_20,
	plif_exmemrtnaddr_l_19,
	plif_exmemrtnaddr_l_18,
	plif_exmemrtnaddr_l_17,
	plif_exmemrtnaddr_l_16,
	plif_exmemrtnaddr_l_15,
	plif_exmemrtnaddr_l_14,
	plif_exmemrtnaddr_l_13,
	plif_exmemrtnaddr_l_12,
	plif_exmemrtnaddr_l_11,
	plif_exmemrtnaddr_l_10,
	plif_exmemrtnaddr_l_9,
	plif_exmemrtnaddr_l_8,
	plif_exmemrtnaddr_l_7,
	plif_exmemrtnaddr_l_6,
	plif_exmemrtnaddr_l_5,
	plif_exmemrtnaddr_l_2,
	plif_exmemrtnaddr_l_1,
	plif_exmemrtnaddr_l_0,
	plif_exmemrtnaddr_l_4,
	plif_exmemrtnaddr_l_3,
	plif_exmembtype_l,
	plif_exmemzero_l,
	plif_exmemjaddr_l_1,
	plif_exmemextimm_l_1,
	plif_exmemextimm_l_0,
	plif_exmemjaddr_l_0,
	plif_exmemjaddr_l_3,
	plif_exmemextimm_l_3,
	plif_exmemextimm_l_2,
	plif_exmemjaddr_l_2,
	plif_exmemjaddr_l_5,
	plif_exmemextimm_l_5,
	plif_exmemextimm_l_4,
	plif_exmemjaddr_l_4,
	plif_exmemjaddr_l_7,
	plif_exmemextimm_l_7,
	plif_exmemextimm_l_6,
	plif_exmemjaddr_l_6,
	plif_exmemjaddr_l_9,
	plif_exmemextimm_l_9,
	plif_exmemextimm_l_8,
	plif_exmemjaddr_l_8,
	plif_exmemjaddr_l_11,
	plif_exmemextimm_l_11,
	plif_exmemextimm_l_10,
	plif_exmemjaddr_l_10,
	plif_exmemjaddr_l_13,
	plif_exmemextimm_l_13,
	plif_exmemextimm_l_12,
	plif_exmemjaddr_l_12,
	plif_exmemjaddr_l_15,
	plif_exmemextimm_l_15,
	plif_exmemextimm_l_14,
	plif_exmemjaddr_l_14,
	plif_exmemjaddr_l_17,
	plif_exmemextimm_l_17,
	plif_exmemextimm_l_16,
	plif_exmemjaddr_l_16,
	plif_exmemjaddr_l_19,
	plif_exmemextimm_l_19,
	plif_exmemextimm_l_18,
	plif_exmemjaddr_l_18,
	plif_exmemjaddr_l_21,
	plif_exmemextimm_l_21,
	plif_exmemextimm_l_20,
	plif_exmemjaddr_l_20,
	plif_exmemjaddr_l_23,
	plif_exmemextimm_l_23,
	plif_exmemextimm_l_22,
	plif_exmemjaddr_l_22,
	plif_exmemjaddr_l_25,
	plif_exmemextimm_l_25,
	plif_exmemextimm_l_24,
	plif_exmemjaddr_l_24,
	plif_exmemextimm_l_27,
	plif_exmemextimm_l_26,
	plif_exmemextimm_l_29,
	plif_exmemextimm_l_28,
	plif_idexregsrc_l_0,
	plif_idexregsrc_l_1,
	plif_idexrtnaddr_l_31,
	plif_idexrtnaddr_l_30,
	plif_idexrtnaddr_l_29,
	plif_idexrtnaddr_l_28,
	plif_idexrtnaddr_l_27,
	plif_idexrtnaddr_l_26,
	plif_idexrtnaddr_l_25,
	plif_idexrtnaddr_l_24,
	plif_idexrtnaddr_l_23,
	plif_idexrtnaddr_l_22,
	plif_idexrtnaddr_l_21,
	plif_idexrtnaddr_l_20,
	plif_idexrtnaddr_l_19,
	plif_idexrtnaddr_l_18,
	plif_idexrtnaddr_l_17,
	plif_idexrtnaddr_l_16,
	plif_idexrtnaddr_l_15,
	plif_idexrtnaddr_l_14,
	plif_idexrtnaddr_l_13,
	plif_idexrtnaddr_l_12,
	plif_idexrtnaddr_l_11,
	plif_idexrtnaddr_l_10,
	plif_idexrtnaddr_l_9,
	plif_idexrtnaddr_l_8,
	plif_idexrtnaddr_l_7,
	plif_idexrtnaddr_l_6,
	plif_idexrtnaddr_l_5,
	plif_idexrtnaddr_l_2,
	plif_idexrtnaddr_l_1,
	plif_idexrtnaddr_l_0,
	plif_idexrtnaddr_l_4,
	plif_idexrtnaddr_l_3,
	plif_idexbtype_l,
	WideOr1,
	plif_idexjaddr_l_1,
	plif_idexjaddr_l_0,
	plif_idexjaddr_l_3,
	plif_idexjaddr_l_2,
	plif_idexjaddr_l_5,
	plif_idexjaddr_l_4,
	plif_idexjaddr_l_7,
	plif_idexjaddr_l_6,
	plif_idexjaddr_l_9,
	plif_idexjaddr_l_8,
	plif_idexjaddr_l_11,
	plif_idexjaddr_l_10,
	plif_idexjaddr_l_13,
	plif_idexjaddr_l_12,
	plif_idexjaddr_l_15,
	plif_idexjaddr_l_14,
	plif_idexjaddr_l_17,
	plif_idexjaddr_l_16,
	plif_idexjaddr_l_19,
	plif_idexjaddr_l_18,
	plif_idexjaddr_l_21,
	plif_idexjaddr_l_20,
	plif_idexjaddr_l_23,
	plif_idexjaddr_l_22,
	plif_idexjaddr_l_25,
	plif_idexjaddr_l_24,
	rdat2,
	rdat21,
	rdat22,
	rdat23,
	rdat24,
	rdat25,
	rdat26,
	rdat27,
	rdat28,
	rdat29,
	rdat210,
	rdat211,
	rdat212,
	rdat213,
	rdat214,
	rdat215,
	rdat216,
	rdat217,
	rdat218,
	rdat219,
	rdat220,
	rdat221,
	rdat222,
	rdat223,
	rdat224,
	rdat225,
	rdat226,
	rdat227,
	rdat228,
	rdat229,
	rdat230,
	rdat231,
	CPUCLK,
	nRST,
	devpor,
	devclrn,
	devoe);
output 	plif_exmemhlt_l;
output 	plif_exmemporto_l_1;
output 	plif_exmemdmemWEN_l;
output 	plif_exmemdmemREN_l;
output 	plif_exmemporto_l_0;
output 	plif_exmemporto_l_3;
output 	plif_exmemporto_l_2;
output 	plif_exmemporto_l_5;
output 	plif_exmemporto_l_4;
output 	plif_exmemporto_l_7;
output 	plif_exmemporto_l_6;
output 	plif_exmemporto_l_9;
output 	plif_exmemporto_l_8;
output 	plif_exmemporto_l_11;
output 	plif_exmemporto_l_10;
output 	plif_exmemporto_l_13;
output 	plif_exmemporto_l_12;
output 	plif_exmemporto_l_15;
output 	plif_exmemporto_l_14;
output 	plif_exmemporto_l_17;
output 	plif_exmemporto_l_16;
output 	plif_exmemporto_l_19;
output 	plif_exmemporto_l_18;
output 	plif_exmemporto_l_21;
output 	plif_exmemporto_l_20;
output 	plif_exmemporto_l_23;
output 	plif_exmemporto_l_22;
output 	plif_exmemporto_l_25;
output 	plif_exmemporto_l_24;
output 	plif_exmemporto_l_27;
output 	plif_exmemporto_l_26;
output 	plif_exmemporto_l_29;
output 	plif_exmemporto_l_28;
output 	plif_exmemporto_l_31;
output 	plif_exmemporto_l_30;
input 	plif_idexhlt_l;
input 	plif_idexpcsrc_l_1;
input 	plif_idexpcsrc_l_0;
output 	plif_exmempcsrc_l_1;
output 	plif_exmempcsrc_l_0;
input 	exmem_en;
output 	plif_exmemrdat2_l_0;
output 	plif_exmemregen_l;
output 	plif_exmemwsel_l_0;
output 	plif_exmemwsel_l_1;
output 	plif_exmemwsel_l_4;
output 	plif_exmemwsel_l_3;
output 	plif_exmemwsel_l_2;
input 	plif_idexextimm_l_29;
input 	plif_idexextimm_l_28;
input 	plif_idexextimm_l_27;
input 	plif_idexextimm_l_26;
input 	plif_idexextimm_l_25;
input 	plif_idexextimm_l_24;
input 	plif_idexextimm_l_23;
input 	plif_idexextimm_l_22;
input 	plif_idexextimm_l_21;
input 	plif_idexextimm_l_20;
input 	plif_idexextimm_l_19;
input 	plif_idexextimm_l_18;
input 	plif_idexextimm_l_17;
input 	plif_idexextimm_l_16;
input 	plif_idexextimm_l_15;
input 	plif_idexextimm_l_14;
input 	plif_idexextimm_l_13;
input 	plif_idexextimm_l_12;
input 	plif_idexextimm_l_11;
input 	plif_idexextimm_l_10;
input 	plif_idexextimm_l_9;
input 	plif_idexextimm_l_8;
input 	plif_idexextimm_l_7;
input 	plif_idexextimm_l_6;
input 	plif_idexextimm_l_5;
input 	plif_idexextimm_l_0;
input 	plif_idexextimm_l_1;
input 	plif_idexextimm_l_2;
input 	plif_idexextimm_l_3;
input 	plif_idexextimm_l_4;
input 	Selector30;
input 	plif_idexdmemREN_l;
input 	plif_idexwsel_l_0;
input 	plif_idexwsel_l_1;
input 	plif_idexwsel_l_2;
input 	plif_idexwsel_l_3;
input 	plif_idexwsel_l_4;
input 	plif_idexdmemWEN_l;
input 	Selector31;
input 	Selector28;
input 	Selector29;
input 	Selector26;
input 	Selector27;
input 	Selector24;
input 	Selector25;
input 	Selector22;
input 	Selector23;
input 	Selector20;
input 	Selector21;
input 	Selector18;
input 	Selector19;
input 	Selector16;
input 	Selector17;
input 	Selector14;
input 	Selector15;
input 	Selector12;
input 	Selector13;
input 	Selector10;
input 	Selector11;
input 	Selector8;
input 	Selector9;
input 	Selector6;
input 	Selector7;
input 	Selector4;
input 	Selector5;
input 	Selector2;
input 	Selector3;
input 	Selector0;
input 	Selector1;
output 	plif_exmemrdat2_l_1;
output 	plif_exmemrdat2_l_2;
output 	plif_exmemrdat2_l_3;
output 	plif_exmemrdat2_l_4;
output 	plif_exmemrdat2_l_5;
output 	plif_exmemrdat2_l_6;
output 	plif_exmemrdat2_l_7;
output 	plif_exmemrdat2_l_8;
output 	plif_exmemrdat2_l_9;
output 	plif_exmemrdat2_l_10;
output 	plif_exmemrdat2_l_11;
output 	plif_exmemrdat2_l_12;
output 	plif_exmemrdat2_l_13;
output 	plif_exmemrdat2_l_14;
output 	plif_exmemrdat2_l_15;
output 	plif_exmemrdat2_l_16;
output 	plif_exmemrdat2_l_17;
output 	plif_exmemrdat2_l_18;
output 	plif_exmemrdat2_l_19;
output 	plif_exmemrdat2_l_20;
output 	plif_exmemrdat2_l_21;
output 	plif_exmemrdat2_l_22;
output 	plif_exmemrdat2_l_23;
output 	plif_exmemrdat2_l_24;
output 	plif_exmemrdat2_l_25;
output 	plif_exmemrdat2_l_26;
output 	plif_exmemrdat2_l_27;
output 	plif_exmemrdat2_l_28;
output 	plif_exmemrdat2_l_29;
output 	plif_exmemrdat2_l_30;
output 	plif_exmemrdat2_l_31;
input 	plif_idexregen_l;
output 	plif_exmemregsrc_l_0;
output 	plif_exmemregsrc_l_1;
output 	plif_exmemrtnaddr_l_31;
output 	plif_exmemrtnaddr_l_30;
output 	plif_exmemrtnaddr_l_29;
output 	plif_exmemrtnaddr_l_28;
output 	plif_exmemrtnaddr_l_27;
output 	plif_exmemrtnaddr_l_26;
output 	plif_exmemrtnaddr_l_25;
output 	plif_exmemrtnaddr_l_24;
output 	plif_exmemrtnaddr_l_23;
output 	plif_exmemrtnaddr_l_22;
output 	plif_exmemrtnaddr_l_21;
output 	plif_exmemrtnaddr_l_20;
output 	plif_exmemrtnaddr_l_19;
output 	plif_exmemrtnaddr_l_18;
output 	plif_exmemrtnaddr_l_17;
output 	plif_exmemrtnaddr_l_16;
output 	plif_exmemrtnaddr_l_15;
output 	plif_exmemrtnaddr_l_14;
output 	plif_exmemrtnaddr_l_13;
output 	plif_exmemrtnaddr_l_12;
output 	plif_exmemrtnaddr_l_11;
output 	plif_exmemrtnaddr_l_10;
output 	plif_exmemrtnaddr_l_9;
output 	plif_exmemrtnaddr_l_8;
output 	plif_exmemrtnaddr_l_7;
output 	plif_exmemrtnaddr_l_6;
output 	plif_exmemrtnaddr_l_5;
output 	plif_exmemrtnaddr_l_2;
output 	plif_exmemrtnaddr_l_1;
output 	plif_exmemrtnaddr_l_0;
output 	plif_exmemrtnaddr_l_4;
output 	plif_exmemrtnaddr_l_3;
output 	plif_exmembtype_l;
output 	plif_exmemzero_l;
output 	plif_exmemjaddr_l_1;
output 	plif_exmemextimm_l_1;
output 	plif_exmemextimm_l_0;
output 	plif_exmemjaddr_l_0;
output 	plif_exmemjaddr_l_3;
output 	plif_exmemextimm_l_3;
output 	plif_exmemextimm_l_2;
output 	plif_exmemjaddr_l_2;
output 	plif_exmemjaddr_l_5;
output 	plif_exmemextimm_l_5;
output 	plif_exmemextimm_l_4;
output 	plif_exmemjaddr_l_4;
output 	plif_exmemjaddr_l_7;
output 	plif_exmemextimm_l_7;
output 	plif_exmemextimm_l_6;
output 	plif_exmemjaddr_l_6;
output 	plif_exmemjaddr_l_9;
output 	plif_exmemextimm_l_9;
output 	plif_exmemextimm_l_8;
output 	plif_exmemjaddr_l_8;
output 	plif_exmemjaddr_l_11;
output 	plif_exmemextimm_l_11;
output 	plif_exmemextimm_l_10;
output 	plif_exmemjaddr_l_10;
output 	plif_exmemjaddr_l_13;
output 	plif_exmemextimm_l_13;
output 	plif_exmemextimm_l_12;
output 	plif_exmemjaddr_l_12;
output 	plif_exmemjaddr_l_15;
output 	plif_exmemextimm_l_15;
output 	plif_exmemextimm_l_14;
output 	plif_exmemjaddr_l_14;
output 	plif_exmemjaddr_l_17;
output 	plif_exmemextimm_l_17;
output 	plif_exmemextimm_l_16;
output 	plif_exmemjaddr_l_16;
output 	plif_exmemjaddr_l_19;
output 	plif_exmemextimm_l_19;
output 	plif_exmemextimm_l_18;
output 	plif_exmemjaddr_l_18;
output 	plif_exmemjaddr_l_21;
output 	plif_exmemextimm_l_21;
output 	plif_exmemextimm_l_20;
output 	plif_exmemjaddr_l_20;
output 	plif_exmemjaddr_l_23;
output 	plif_exmemextimm_l_23;
output 	plif_exmemextimm_l_22;
output 	plif_exmemjaddr_l_22;
output 	plif_exmemjaddr_l_25;
output 	plif_exmemextimm_l_25;
output 	plif_exmemextimm_l_24;
output 	plif_exmemjaddr_l_24;
output 	plif_exmemextimm_l_27;
output 	plif_exmemextimm_l_26;
output 	plif_exmemextimm_l_29;
output 	plif_exmemextimm_l_28;
input 	plif_idexregsrc_l_0;
input 	plif_idexregsrc_l_1;
input 	plif_idexrtnaddr_l_31;
input 	plif_idexrtnaddr_l_30;
input 	plif_idexrtnaddr_l_29;
input 	plif_idexrtnaddr_l_28;
input 	plif_idexrtnaddr_l_27;
input 	plif_idexrtnaddr_l_26;
input 	plif_idexrtnaddr_l_25;
input 	plif_idexrtnaddr_l_24;
input 	plif_idexrtnaddr_l_23;
input 	plif_idexrtnaddr_l_22;
input 	plif_idexrtnaddr_l_21;
input 	plif_idexrtnaddr_l_20;
input 	plif_idexrtnaddr_l_19;
input 	plif_idexrtnaddr_l_18;
input 	plif_idexrtnaddr_l_17;
input 	plif_idexrtnaddr_l_16;
input 	plif_idexrtnaddr_l_15;
input 	plif_idexrtnaddr_l_14;
input 	plif_idexrtnaddr_l_13;
input 	plif_idexrtnaddr_l_12;
input 	plif_idexrtnaddr_l_11;
input 	plif_idexrtnaddr_l_10;
input 	plif_idexrtnaddr_l_9;
input 	plif_idexrtnaddr_l_8;
input 	plif_idexrtnaddr_l_7;
input 	plif_idexrtnaddr_l_6;
input 	plif_idexrtnaddr_l_5;
input 	plif_idexrtnaddr_l_2;
input 	plif_idexrtnaddr_l_1;
input 	plif_idexrtnaddr_l_0;
input 	plif_idexrtnaddr_l_4;
input 	plif_idexrtnaddr_l_3;
input 	plif_idexbtype_l;
input 	WideOr1;
input 	plif_idexjaddr_l_1;
input 	plif_idexjaddr_l_0;
input 	plif_idexjaddr_l_3;
input 	plif_idexjaddr_l_2;
input 	plif_idexjaddr_l_5;
input 	plif_idexjaddr_l_4;
input 	plif_idexjaddr_l_7;
input 	plif_idexjaddr_l_6;
input 	plif_idexjaddr_l_9;
input 	plif_idexjaddr_l_8;
input 	plif_idexjaddr_l_11;
input 	plif_idexjaddr_l_10;
input 	plif_idexjaddr_l_13;
input 	plif_idexjaddr_l_12;
input 	plif_idexjaddr_l_15;
input 	plif_idexjaddr_l_14;
input 	plif_idexjaddr_l_17;
input 	plif_idexjaddr_l_16;
input 	plif_idexjaddr_l_19;
input 	plif_idexjaddr_l_18;
input 	plif_idexjaddr_l_21;
input 	plif_idexjaddr_l_20;
input 	plif_idexjaddr_l_23;
input 	plif_idexjaddr_l_22;
input 	plif_idexjaddr_l_25;
input 	plif_idexjaddr_l_24;
input 	rdat2;
input 	rdat21;
input 	rdat22;
input 	rdat23;
input 	rdat24;
input 	rdat25;
input 	rdat26;
input 	rdat27;
input 	rdat28;
input 	rdat29;
input 	rdat210;
input 	rdat211;
input 	rdat212;
input 	rdat213;
input 	rdat214;
input 	rdat215;
input 	rdat216;
input 	rdat217;
input 	rdat218;
input 	rdat219;
input 	rdat220;
input 	rdat221;
input 	rdat222;
input 	rdat223;
input 	rdat224;
input 	rdat225;
input 	rdat226;
input 	rdat227;
input 	rdat228;
input 	rdat229;
input 	rdat230;
input 	rdat231;
input 	CPUCLK;
input 	nRST;

// Design Ports Information

input 	devpor;
input 	devclrn;
input 	devoe;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
assign unknown = 1'bx;

wire \plif_exmem.porto_l[1]~feeder_combout ;
wire \plif_exmem.porto_l[5]~feeder_combout ;
wire \plif_exmem.porto_l[7]~feeder_combout ;
wire \plif_exmem.porto_l[8]~feeder_combout ;
wire \plif_exmem.porto_l[11]~feeder_combout ;
wire \plif_exmem.porto_l[12]~feeder_combout ;
wire \plif_exmem.porto_l[14]~feeder_combout ;
wire \plif_exmem.porto_l[16]~feeder_combout ;
wire \plif_exmem.porto_l[21]~feeder_combout ;
wire \plif_exmem.porto_l[20]~feeder_combout ;
wire \plif_exmem.pcsrc_l[1]~feeder_combout ;
wire \plif_exmem.pcsrc_l[0]~feeder_combout ;
wire \plif_exmem.regsrc_l[0]~feeder_combout ;
wire \plif_exmem.rtnaddr_l[31]~feeder_combout ;
wire \plif_exmem.rtnaddr_l[27]~feeder_combout ;
wire \plif_exmem.rtnaddr_l[24]~feeder_combout ;
wire \plif_exmem.rtnaddr_l[23]~feeder_combout ;
wire \plif_exmem.rtnaddr_l[21]~feeder_combout ;
wire \plif_exmem.rtnaddr_l[20]~feeder_combout ;
wire \plif_exmem.rtnaddr_l[19]~feeder_combout ;
wire \plif_exmem.rtnaddr_l[17]~feeder_combout ;
wire \plif_exmem.rtnaddr_l[15]~feeder_combout ;
wire \plif_exmem.rtnaddr_l[13]~feeder_combout ;
wire \plif_exmem.rtnaddr_l[12]~feeder_combout ;
wire \plif_exmem.rtnaddr_l[11]~feeder_combout ;
wire \plif_exmem.rtnaddr_l[9]~feeder_combout ;
wire \plif_exmem.rtnaddr_l[8]~feeder_combout ;
wire \plif_exmem.rtnaddr_l[7]~feeder_combout ;
wire \plif_exmem.rtnaddr_l[2]~feeder_combout ;
wire \plif_exmem.rtnaddr_l[4]~feeder_combout ;
wire \plif_exmem.rtnaddr_l[3]~feeder_combout ;
wire \plif_exmem.extimm_l[3]~feeder_combout ;
wire \plif_exmem.jaddr_l[2]~feeder_combout ;
wire \plif_exmem.extimm_l[4]~feeder_combout ;
wire \plif_exmem.jaddr_l[7]~feeder_combout ;
wire \plif_exmem.jaddr_l[9]~feeder_combout ;
wire \plif_exmem.jaddr_l[8]~feeder_combout ;
wire \plif_exmem.jaddr_l[11]~feeder_combout ;
wire \plif_exmem.extimm_l[10]~feeder_combout ;
wire \plif_exmem.jaddr_l[13]~feeder_combout ;
wire \plif_exmem.extimm_l[12]~feeder_combout ;
wire \plif_exmem.jaddr_l[12]~feeder_combout ;
wire \plif_exmem.jaddr_l[15]~feeder_combout ;
wire \plif_exmem.extimm_l[15]~feeder_combout ;
wire \plif_exmem.extimm_l[14]~feeder_combout ;
wire \plif_exmem.jaddr_l[14]~feeder_combout ;
wire \plif_exmem.jaddr_l[17]~feeder_combout ;
wire \plif_exmem.extimm_l[16]~feeder_combout ;
wire \plif_exmem.jaddr_l[16]~feeder_combout ;
wire \plif_exmem.jaddr_l[19]~feeder_combout ;
wire \plif_exmem.extimm_l[18]~feeder_combout ;
wire \plif_exmem.jaddr_l[21]~feeder_combout ;
wire \plif_exmem.extimm_l[21]~feeder_combout ;
wire \plif_exmem.jaddr_l[20]~feeder_combout ;
wire \plif_exmem.jaddr_l[23]~feeder_combout ;
wire \plif_exmem.extimm_l[22]~feeder_combout ;
wire \plif_exmem.jaddr_l[22]~feeder_combout ;
wire \plif_exmem.jaddr_l[25]~feeder_combout ;
wire \plif_exmem.jaddr_l[24]~feeder_combout ;


// Location: DDIOOUTCELL_X49_Y0_N4
dffeas \plif_exmem.hlt_l (
	.clk(CPUCLK),
	.d(plif_idexhlt_l),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(exmem_en),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(plif_exmemhlt_l),
	.prn(vcc));
// synopsys translate_off
defparam \plif_exmem.hlt_l .is_wysiwyg = "true";
defparam \plif_exmem.hlt_l .power_up = "low";
// synopsys translate_on

// Location: FF_X53_Y39_N17
dffeas \plif_exmem.porto_l[1] (
	.clk(CPUCLK),
	.d(\plif_exmem.porto_l[1]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(exmem_en),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(plif_exmemporto_l_1),
	.prn(vcc));
// synopsys translate_off
defparam \plif_exmem.porto_l[1] .is_wysiwyg = "true";
defparam \plif_exmem.porto_l[1] .power_up = "low";
// synopsys translate_on

// Location: FF_X53_Y34_N21
dffeas \plif_exmem.dmemWEN_l (
	.clk(CPUCLK),
	.d(gnd),
	.asdata(plif_idexdmemWEN_l),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(exmem_en),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(plif_exmemdmemWEN_l),
	.prn(vcc));
// synopsys translate_off
defparam \plif_exmem.dmemWEN_l .is_wysiwyg = "true";
defparam \plif_exmem.dmemWEN_l .power_up = "low";
// synopsys translate_on

// Location: FF_X53_Y34_N7
dffeas \plif_exmem.dmemREN_l (
	.clk(CPUCLK),
	.d(gnd),
	.asdata(plif_idexdmemREN_l),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(exmem_en),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(plif_exmemdmemREN_l),
	.prn(vcc));
// synopsys translate_off
defparam \plif_exmem.dmemREN_l .is_wysiwyg = "true";
defparam \plif_exmem.dmemREN_l .power_up = "low";
// synopsys translate_on

// Location: FF_X50_Y39_N1
dffeas \plif_exmem.porto_l[0] (
	.clk(CPUCLK),
	.d(Selector31),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(exmem_en),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(plif_exmemporto_l_0),
	.prn(vcc));
// synopsys translate_off
defparam \plif_exmem.porto_l[0] .is_wysiwyg = "true";
defparam \plif_exmem.porto_l[0] .power_up = "low";
// synopsys translate_on

// Location: FF_X52_Y40_N21
dffeas \plif_exmem.porto_l[3] (
	.clk(CPUCLK),
	.d(Selector28),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(exmem_en),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(plif_exmemporto_l_3),
	.prn(vcc));
// synopsys translate_off
defparam \plif_exmem.porto_l[3] .is_wysiwyg = "true";
defparam \plif_exmem.porto_l[3] .power_up = "low";
// synopsys translate_on

// Location: FF_X52_Y40_N31
dffeas \plif_exmem.porto_l[2] (
	.clk(CPUCLK),
	.d(Selector29),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(exmem_en),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(plif_exmemporto_l_2),
	.prn(vcc));
// synopsys translate_off
defparam \plif_exmem.porto_l[2] .is_wysiwyg = "true";
defparam \plif_exmem.porto_l[2] .power_up = "low";
// synopsys translate_on

// Location: FF_X50_Y41_N17
dffeas \plif_exmem.porto_l[5] (
	.clk(CPUCLK),
	.d(\plif_exmem.porto_l[5]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(exmem_en),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(plif_exmemporto_l_5),
	.prn(vcc));
// synopsys translate_off
defparam \plif_exmem.porto_l[5] .is_wysiwyg = "true";
defparam \plif_exmem.porto_l[5] .power_up = "low";
// synopsys translate_on

// Location: FF_X50_Y38_N29
dffeas \plif_exmem.porto_l[4] (
	.clk(CPUCLK),
	.d(gnd),
	.asdata(Selector27),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(exmem_en),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(plif_exmemporto_l_4),
	.prn(vcc));
// synopsys translate_off
defparam \plif_exmem.porto_l[4] .is_wysiwyg = "true";
defparam \plif_exmem.porto_l[4] .power_up = "low";
// synopsys translate_on

// Location: FF_X53_Y42_N1
dffeas \plif_exmem.porto_l[7] (
	.clk(CPUCLK),
	.d(\plif_exmem.porto_l[7]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(exmem_en),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(plif_exmemporto_l_7),
	.prn(vcc));
// synopsys translate_off
defparam \plif_exmem.porto_l[7] .is_wysiwyg = "true";
defparam \plif_exmem.porto_l[7] .power_up = "low";
// synopsys translate_on

// Location: FF_X55_Y39_N21
dffeas \plif_exmem.porto_l[6] (
	.clk(CPUCLK),
	.d(gnd),
	.asdata(Selector25),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(exmem_en),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(plif_exmemporto_l_6),
	.prn(vcc));
// synopsys translate_off
defparam \plif_exmem.porto_l[6] .is_wysiwyg = "true";
defparam \plif_exmem.porto_l[6] .power_up = "low";
// synopsys translate_on

// Location: FF_X53_Y41_N17
dffeas \plif_exmem.porto_l[9] (
	.clk(CPUCLK),
	.d(gnd),
	.asdata(Selector22),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(exmem_en),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(plif_exmemporto_l_9),
	.prn(vcc));
// synopsys translate_off
defparam \plif_exmem.porto_l[9] .is_wysiwyg = "true";
defparam \plif_exmem.porto_l[9] .power_up = "low";
// synopsys translate_on

// Location: FF_X53_Y40_N29
dffeas \plif_exmem.porto_l[8] (
	.clk(CPUCLK),
	.d(\plif_exmem.porto_l[8]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(exmem_en),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(plif_exmemporto_l_8),
	.prn(vcc));
// synopsys translate_off
defparam \plif_exmem.porto_l[8] .is_wysiwyg = "true";
defparam \plif_exmem.porto_l[8] .power_up = "low";
// synopsys translate_on

// Location: FF_X54_Y37_N17
dffeas \plif_exmem.porto_l[11] (
	.clk(CPUCLK),
	.d(\plif_exmem.porto_l[11]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(exmem_en),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(plif_exmemporto_l_11),
	.prn(vcc));
// synopsys translate_off
defparam \plif_exmem.porto_l[11] .is_wysiwyg = "true";
defparam \plif_exmem.porto_l[11] .power_up = "low";
// synopsys translate_on

// Location: FF_X54_Y37_N1
dffeas \plif_exmem.porto_l[10] (
	.clk(CPUCLK),
	.d(Selector21),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(exmem_en),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(plif_exmemporto_l_10),
	.prn(vcc));
// synopsys translate_off
defparam \plif_exmem.porto_l[10] .is_wysiwyg = "true";
defparam \plif_exmem.porto_l[10] .power_up = "low";
// synopsys translate_on

// Location: FF_X53_Y38_N29
dffeas \plif_exmem.porto_l[13] (
	.clk(CPUCLK),
	.d(gnd),
	.asdata(Selector18),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(exmem_en),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(plif_exmemporto_l_13),
	.prn(vcc));
// synopsys translate_off
defparam \plif_exmem.porto_l[13] .is_wysiwyg = "true";
defparam \plif_exmem.porto_l[13] .power_up = "low";
// synopsys translate_on

// Location: FF_X53_Y40_N3
dffeas \plif_exmem.porto_l[12] (
	.clk(CPUCLK),
	.d(\plif_exmem.porto_l[12]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(exmem_en),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(plif_exmemporto_l_12),
	.prn(vcc));
// synopsys translate_off
defparam \plif_exmem.porto_l[12] .is_wysiwyg = "true";
defparam \plif_exmem.porto_l[12] .power_up = "low";
// synopsys translate_on

// Location: FF_X52_Y36_N1
dffeas \plif_exmem.porto_l[15] (
	.clk(CPUCLK),
	.d(gnd),
	.asdata(Selector16),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(exmem_en),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(plif_exmemporto_l_15),
	.prn(vcc));
// synopsys translate_off
defparam \plif_exmem.porto_l[15] .is_wysiwyg = "true";
defparam \plif_exmem.porto_l[15] .power_up = "low";
// synopsys translate_on

// Location: FF_X53_Y39_N31
dffeas \plif_exmem.porto_l[14] (
	.clk(CPUCLK),
	.d(\plif_exmem.porto_l[14]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(exmem_en),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(plif_exmemporto_l_14),
	.prn(vcc));
// synopsys translate_off
defparam \plif_exmem.porto_l[14] .is_wysiwyg = "true";
defparam \plif_exmem.porto_l[14] .power_up = "low";
// synopsys translate_on

// Location: FF_X54_Y41_N5
dffeas \plif_exmem.porto_l[17] (
	.clk(CPUCLK),
	.d(gnd),
	.asdata(Selector14),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(exmem_en),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(plif_exmemporto_l_17),
	.prn(vcc));
// synopsys translate_off
defparam \plif_exmem.porto_l[17] .is_wysiwyg = "true";
defparam \plif_exmem.porto_l[17] .power_up = "low";
// synopsys translate_on

// Location: FF_X52_Y35_N25
dffeas \plif_exmem.porto_l[16] (
	.clk(CPUCLK),
	.d(\plif_exmem.porto_l[16]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(exmem_en),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(plif_exmemporto_l_16),
	.prn(vcc));
// synopsys translate_off
defparam \plif_exmem.porto_l[16] .is_wysiwyg = "true";
defparam \plif_exmem.porto_l[16] .power_up = "low";
// synopsys translate_on

// Location: FF_X53_Y37_N9
dffeas \plif_exmem.porto_l[19] (
	.clk(CPUCLK),
	.d(gnd),
	.asdata(Selector12),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(exmem_en),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(plif_exmemporto_l_19),
	.prn(vcc));
// synopsys translate_off
defparam \plif_exmem.porto_l[19] .is_wysiwyg = "true";
defparam \plif_exmem.porto_l[19] .power_up = "low";
// synopsys translate_on

// Location: FF_X55_Y37_N9
dffeas \plif_exmem.porto_l[18] (
	.clk(CPUCLK),
	.d(Selector13),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(exmem_en),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(plif_exmemporto_l_18),
	.prn(vcc));
// synopsys translate_off
defparam \plif_exmem.porto_l[18] .is_wysiwyg = "true";
defparam \plif_exmem.porto_l[18] .power_up = "low";
// synopsys translate_on

// Location: FF_X54_Y42_N21
dffeas \plif_exmem.porto_l[21] (
	.clk(CPUCLK),
	.d(\plif_exmem.porto_l[21]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(exmem_en),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(plif_exmemporto_l_21),
	.prn(vcc));
// synopsys translate_off
defparam \plif_exmem.porto_l[21] .is_wysiwyg = "true";
defparam \plif_exmem.porto_l[21] .power_up = "low";
// synopsys translate_on

// Location: FF_X54_Y39_N23
dffeas \plif_exmem.porto_l[20] (
	.clk(CPUCLK),
	.d(\plif_exmem.porto_l[20]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(exmem_en),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(plif_exmemporto_l_20),
	.prn(vcc));
// synopsys translate_off
defparam \plif_exmem.porto_l[20] .is_wysiwyg = "true";
defparam \plif_exmem.porto_l[20] .power_up = "low";
// synopsys translate_on

// Location: FF_X52_Y39_N5
dffeas \plif_exmem.porto_l[23] (
	.clk(CPUCLK),
	.d(gnd),
	.asdata(Selector8),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(exmem_en),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(plif_exmemporto_l_23),
	.prn(vcc));
// synopsys translate_off
defparam \plif_exmem.porto_l[23] .is_wysiwyg = "true";
defparam \plif_exmem.porto_l[23] .power_up = "low";
// synopsys translate_on

// Location: FF_X52_Y39_N11
dffeas \plif_exmem.porto_l[22] (
	.clk(CPUCLK),
	.d(gnd),
	.asdata(Selector9),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(exmem_en),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(plif_exmemporto_l_22),
	.prn(vcc));
// synopsys translate_off
defparam \plif_exmem.porto_l[22] .is_wysiwyg = "true";
defparam \plif_exmem.porto_l[22] .power_up = "low";
// synopsys translate_on

// Location: FF_X54_Y36_N29
dffeas \plif_exmem.porto_l[25] (
	.clk(CPUCLK),
	.d(gnd),
	.asdata(Selector6),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(exmem_en),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(plif_exmemporto_l_25),
	.prn(vcc));
// synopsys translate_off
defparam \plif_exmem.porto_l[25] .is_wysiwyg = "true";
defparam \plif_exmem.porto_l[25] .power_up = "low";
// synopsys translate_on

// Location: FF_X53_Y35_N13
dffeas \plif_exmem.porto_l[24] (
	.clk(CPUCLK),
	.d(Selector7),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(exmem_en),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(plif_exmemporto_l_24),
	.prn(vcc));
// synopsys translate_off
defparam \plif_exmem.porto_l[24] .is_wysiwyg = "true";
defparam \plif_exmem.porto_l[24] .power_up = "low";
// synopsys translate_on

// Location: FF_X54_Y36_N23
dffeas \plif_exmem.porto_l[27] (
	.clk(CPUCLK),
	.d(gnd),
	.asdata(Selector4),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(exmem_en),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(plif_exmemporto_l_27),
	.prn(vcc));
// synopsys translate_off
defparam \plif_exmem.porto_l[27] .is_wysiwyg = "true";
defparam \plif_exmem.porto_l[27] .power_up = "low";
// synopsys translate_on

// Location: FF_X54_Y36_N9
dffeas \plif_exmem.porto_l[26] (
	.clk(CPUCLK),
	.d(gnd),
	.asdata(Selector5),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(exmem_en),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(plif_exmemporto_l_26),
	.prn(vcc));
// synopsys translate_off
defparam \plif_exmem.porto_l[26] .is_wysiwyg = "true";
defparam \plif_exmem.porto_l[26] .power_up = "low";
// synopsys translate_on

// Location: FF_X50_Y39_N23
dffeas \plif_exmem.porto_l[29] (
	.clk(CPUCLK),
	.d(gnd),
	.asdata(Selector2),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(exmem_en),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(plif_exmemporto_l_29),
	.prn(vcc));
// synopsys translate_off
defparam \plif_exmem.porto_l[29] .is_wysiwyg = "true";
defparam \plif_exmem.porto_l[29] .power_up = "low";
// synopsys translate_on

// Location: FF_X50_Y39_N13
dffeas \plif_exmem.porto_l[28] (
	.clk(CPUCLK),
	.d(gnd),
	.asdata(Selector3),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(exmem_en),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(plif_exmemporto_l_28),
	.prn(vcc));
// synopsys translate_off
defparam \plif_exmem.porto_l[28] .is_wysiwyg = "true";
defparam \plif_exmem.porto_l[28] .power_up = "low";
// synopsys translate_on

// Location: FF_X52_Y42_N29
dffeas \plif_exmem.porto_l[31] (
	.clk(CPUCLK),
	.d(gnd),
	.asdata(Selector0),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(exmem_en),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(plif_exmemporto_l_31),
	.prn(vcc));
// synopsys translate_off
defparam \plif_exmem.porto_l[31] .is_wysiwyg = "true";
defparam \plif_exmem.porto_l[31] .power_up = "low";
// synopsys translate_on

// Location: FF_X55_Y42_N15
dffeas \plif_exmem.porto_l[30] (
	.clk(CPUCLK),
	.d(Selector1),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(exmem_en),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(plif_exmemporto_l_30),
	.prn(vcc));
// synopsys translate_off
defparam \plif_exmem.porto_l[30] .is_wysiwyg = "true";
defparam \plif_exmem.porto_l[30] .power_up = "low";
// synopsys translate_on

// Location: FF_X55_Y32_N31
dffeas \plif_exmem.pcsrc_l[1] (
	.clk(CPUCLK),
	.d(\plif_exmem.pcsrc_l[1]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(exmem_en),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(plif_exmempcsrc_l_1),
	.prn(vcc));
// synopsys translate_off
defparam \plif_exmem.pcsrc_l[1] .is_wysiwyg = "true";
defparam \plif_exmem.pcsrc_l[1] .power_up = "low";
// synopsys translate_on

// Location: FF_X55_Y32_N23
dffeas \plif_exmem.pcsrc_l[0] (
	.clk(CPUCLK),
	.d(\plif_exmem.pcsrc_l[0]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(exmem_en),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(plif_exmempcsrc_l_0),
	.prn(vcc));
// synopsys translate_off
defparam \plif_exmem.pcsrc_l[0] .is_wysiwyg = "true";
defparam \plif_exmem.pcsrc_l[0] .power_up = "low";
// synopsys translate_on

// Location: FF_X59_Y39_N1
dffeas \plif_exmem.rdat2_l[0] (
	.clk(CPUCLK),
	.d(rdat2),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(exmem_en),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(plif_exmemrdat2_l_0),
	.prn(vcc));
// synopsys translate_off
defparam \plif_exmem.rdat2_l[0] .is_wysiwyg = "true";
defparam \plif_exmem.rdat2_l[0] .power_up = "low";
// synopsys translate_on

// Location: FF_X57_Y37_N15
dffeas \plif_exmem.regen_l (
	.clk(CPUCLK),
	.d(gnd),
	.asdata(plif_idexregen_l),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(exmem_en),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(plif_exmemregen_l),
	.prn(vcc));
// synopsys translate_off
defparam \plif_exmem.regen_l .is_wysiwyg = "true";
defparam \plif_exmem.regen_l .power_up = "low";
// synopsys translate_on

// Location: FF_X57_Y37_N27
dffeas \plif_exmem.wsel_l[0] (
	.clk(CPUCLK),
	.d(gnd),
	.asdata(plif_idexwsel_l_0),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(exmem_en),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(plif_exmemwsel_l_0),
	.prn(vcc));
// synopsys translate_off
defparam \plif_exmem.wsel_l[0] .is_wysiwyg = "true";
defparam \plif_exmem.wsel_l[0] .power_up = "low";
// synopsys translate_on

// Location: FF_X57_Y37_N11
dffeas \plif_exmem.wsel_l[1] (
	.clk(CPUCLK),
	.d(gnd),
	.asdata(plif_idexwsel_l_1),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(exmem_en),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(plif_exmemwsel_l_1),
	.prn(vcc));
// synopsys translate_off
defparam \plif_exmem.wsel_l[1] .is_wysiwyg = "true";
defparam \plif_exmem.wsel_l[1] .power_up = "low";
// synopsys translate_on

// Location: FF_X57_Y37_N31
dffeas \plif_exmem.wsel_l[4] (
	.clk(CPUCLK),
	.d(gnd),
	.asdata(plif_idexwsel_l_4),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(exmem_en),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(plif_exmemwsel_l_4),
	.prn(vcc));
// synopsys translate_off
defparam \plif_exmem.wsel_l[4] .is_wysiwyg = "true";
defparam \plif_exmem.wsel_l[4] .power_up = "low";
// synopsys translate_on

// Location: FF_X57_Y37_N23
dffeas \plif_exmem.wsel_l[3] (
	.clk(CPUCLK),
	.d(gnd),
	.asdata(plif_idexwsel_l_3),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(exmem_en),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(plif_exmemwsel_l_3),
	.prn(vcc));
// synopsys translate_off
defparam \plif_exmem.wsel_l[3] .is_wysiwyg = "true";
defparam \plif_exmem.wsel_l[3] .power_up = "low";
// synopsys translate_on

// Location: FF_X57_Y37_N1
dffeas \plif_exmem.wsel_l[2] (
	.clk(CPUCLK),
	.d(gnd),
	.asdata(plif_idexwsel_l_2),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(exmem_en),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(plif_exmemwsel_l_2),
	.prn(vcc));
// synopsys translate_off
defparam \plif_exmem.wsel_l[2] .is_wysiwyg = "true";
defparam \plif_exmem.wsel_l[2] .power_up = "low";
// synopsys translate_on

// Location: FF_X57_Y35_N3
dffeas \plif_exmem.rdat2_l[1] (
	.clk(CPUCLK),
	.d(rdat21),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(exmem_en),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(plif_exmemrdat2_l_1),
	.prn(vcc));
// synopsys translate_off
defparam \plif_exmem.rdat2_l[1] .is_wysiwyg = "true";
defparam \plif_exmem.rdat2_l[1] .power_up = "low";
// synopsys translate_on

// Location: FF_X56_Y39_N23
dffeas \plif_exmem.rdat2_l[2] (
	.clk(CPUCLK),
	.d(rdat22),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(exmem_en),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(plif_exmemrdat2_l_2),
	.prn(vcc));
// synopsys translate_off
defparam \plif_exmem.rdat2_l[2] .is_wysiwyg = "true";
defparam \plif_exmem.rdat2_l[2] .power_up = "low";
// synopsys translate_on

// Location: FF_X58_Y34_N29
dffeas \plif_exmem.rdat2_l[3] (
	.clk(CPUCLK),
	.d(rdat23),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(exmem_en),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(plif_exmemrdat2_l_3),
	.prn(vcc));
// synopsys translate_off
defparam \plif_exmem.rdat2_l[3] .is_wysiwyg = "true";
defparam \plif_exmem.rdat2_l[3] .power_up = "low";
// synopsys translate_on

// Location: FF_X58_Y41_N19
dffeas \plif_exmem.rdat2_l[4] (
	.clk(CPUCLK),
	.d(rdat24),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(exmem_en),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(plif_exmemrdat2_l_4),
	.prn(vcc));
// synopsys translate_off
defparam \plif_exmem.rdat2_l[4] .is_wysiwyg = "true";
defparam \plif_exmem.rdat2_l[4] .power_up = "low";
// synopsys translate_on

// Location: FF_X59_Y39_N3
dffeas \plif_exmem.rdat2_l[5] (
	.clk(CPUCLK),
	.d(rdat25),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(exmem_en),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(plif_exmemrdat2_l_5),
	.prn(vcc));
// synopsys translate_off
defparam \plif_exmem.rdat2_l[5] .is_wysiwyg = "true";
defparam \plif_exmem.rdat2_l[5] .power_up = "low";
// synopsys translate_on

// Location: FF_X55_Y35_N7
dffeas \plif_exmem.rdat2_l[6] (
	.clk(CPUCLK),
	.d(rdat26),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(exmem_en),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(plif_exmemrdat2_l_6),
	.prn(vcc));
// synopsys translate_off
defparam \plif_exmem.rdat2_l[6] .is_wysiwyg = "true";
defparam \plif_exmem.rdat2_l[6] .power_up = "low";
// synopsys translate_on

// Location: FF_X58_Y34_N13
dffeas \plif_exmem.rdat2_l[7] (
	.clk(CPUCLK),
	.d(rdat27),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(exmem_en),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(plif_exmemrdat2_l_7),
	.prn(vcc));
// synopsys translate_off
defparam \plif_exmem.rdat2_l[7] .is_wysiwyg = "true";
defparam \plif_exmem.rdat2_l[7] .power_up = "low";
// synopsys translate_on

// Location: FF_X58_Y34_N21
dffeas \plif_exmem.rdat2_l[8] (
	.clk(CPUCLK),
	.d(rdat28),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(exmem_en),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(plif_exmemrdat2_l_8),
	.prn(vcc));
// synopsys translate_off
defparam \plif_exmem.rdat2_l[8] .is_wysiwyg = "true";
defparam \plif_exmem.rdat2_l[8] .power_up = "low";
// synopsys translate_on

// Location: FF_X58_Y35_N19
dffeas \plif_exmem.rdat2_l[9] (
	.clk(CPUCLK),
	.d(rdat29),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(exmem_en),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(plif_exmemrdat2_l_9),
	.prn(vcc));
// synopsys translate_off
defparam \plif_exmem.rdat2_l[9] .is_wysiwyg = "true";
defparam \plif_exmem.rdat2_l[9] .power_up = "low";
// synopsys translate_on

// Location: FF_X57_Y34_N15
dffeas \plif_exmem.rdat2_l[10] (
	.clk(CPUCLK),
	.d(rdat210),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(exmem_en),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(plif_exmemrdat2_l_10),
	.prn(vcc));
// synopsys translate_off
defparam \plif_exmem.rdat2_l[10] .is_wysiwyg = "true";
defparam \plif_exmem.rdat2_l[10] .power_up = "low";
// synopsys translate_on

// Location: FF_X58_Y35_N25
dffeas \plif_exmem.rdat2_l[11] (
	.clk(CPUCLK),
	.d(rdat211),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(exmem_en),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(plif_exmemrdat2_l_11),
	.prn(vcc));
// synopsys translate_off
defparam \plif_exmem.rdat2_l[11] .is_wysiwyg = "true";
defparam \plif_exmem.rdat2_l[11] .power_up = "low";
// synopsys translate_on

// Location: FF_X58_Y34_N3
dffeas \plif_exmem.rdat2_l[12] (
	.clk(CPUCLK),
	.d(rdat212),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(exmem_en),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(plif_exmemrdat2_l_12),
	.prn(vcc));
// synopsys translate_off
defparam \plif_exmem.rdat2_l[12] .is_wysiwyg = "true";
defparam \plif_exmem.rdat2_l[12] .power_up = "low";
// synopsys translate_on

// Location: FF_X59_Y39_N27
dffeas \plif_exmem.rdat2_l[13] (
	.clk(CPUCLK),
	.d(rdat213),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(exmem_en),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(plif_exmemrdat2_l_13),
	.prn(vcc));
// synopsys translate_off
defparam \plif_exmem.rdat2_l[13] .is_wysiwyg = "true";
defparam \plif_exmem.rdat2_l[13] .power_up = "low";
// synopsys translate_on

// Location: FF_X58_Y35_N15
dffeas \plif_exmem.rdat2_l[14] (
	.clk(CPUCLK),
	.d(rdat214),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(exmem_en),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(plif_exmemrdat2_l_14),
	.prn(vcc));
// synopsys translate_off
defparam \plif_exmem.rdat2_l[14] .is_wysiwyg = "true";
defparam \plif_exmem.rdat2_l[14] .power_up = "low";
// synopsys translate_on

// Location: FF_X57_Y35_N29
dffeas \plif_exmem.rdat2_l[15] (
	.clk(CPUCLK),
	.d(rdat215),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(exmem_en),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(plif_exmemrdat2_l_15),
	.prn(vcc));
// synopsys translate_off
defparam \plif_exmem.rdat2_l[15] .is_wysiwyg = "true";
defparam \plif_exmem.rdat2_l[15] .power_up = "low";
// synopsys translate_on

// Location: FF_X55_Y35_N13
dffeas \plif_exmem.rdat2_l[16] (
	.clk(CPUCLK),
	.d(rdat216),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(exmem_en),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(plif_exmemrdat2_l_16),
	.prn(vcc));
// synopsys translate_off
defparam \plif_exmem.rdat2_l[16] .is_wysiwyg = "true";
defparam \plif_exmem.rdat2_l[16] .power_up = "low";
// synopsys translate_on

// Location: FF_X59_Y39_N7
dffeas \plif_exmem.rdat2_l[17] (
	.clk(CPUCLK),
	.d(rdat217),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(exmem_en),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(plif_exmemrdat2_l_17),
	.prn(vcc));
// synopsys translate_off
defparam \plif_exmem.rdat2_l[17] .is_wysiwyg = "true";
defparam \plif_exmem.rdat2_l[17] .power_up = "low";
// synopsys translate_on

// Location: FF_X55_Y37_N23
dffeas \plif_exmem.rdat2_l[18] (
	.clk(CPUCLK),
	.d(rdat218),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(exmem_en),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(plif_exmemrdat2_l_18),
	.prn(vcc));
// synopsys translate_off
defparam \plif_exmem.rdat2_l[18] .is_wysiwyg = "true";
defparam \plif_exmem.rdat2_l[18] .power_up = "low";
// synopsys translate_on

// Location: FF_X57_Y34_N9
dffeas \plif_exmem.rdat2_l[19] (
	.clk(CPUCLK),
	.d(rdat219),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(exmem_en),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(plif_exmemrdat2_l_19),
	.prn(vcc));
// synopsys translate_off
defparam \plif_exmem.rdat2_l[19] .is_wysiwyg = "true";
defparam \plif_exmem.rdat2_l[19] .power_up = "low";
// synopsys translate_on

// Location: FF_X54_Y39_N15
dffeas \plif_exmem.rdat2_l[20] (
	.clk(CPUCLK),
	.d(rdat220),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(exmem_en),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(plif_exmemrdat2_l_20),
	.prn(vcc));
// synopsys translate_off
defparam \plif_exmem.rdat2_l[20] .is_wysiwyg = "true";
defparam \plif_exmem.rdat2_l[20] .power_up = "low";
// synopsys translate_on

// Location: FF_X58_Y34_N1
dffeas \plif_exmem.rdat2_l[21] (
	.clk(CPUCLK),
	.d(rdat221),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(exmem_en),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(plif_exmemrdat2_l_21),
	.prn(vcc));
// synopsys translate_off
defparam \plif_exmem.rdat2_l[21] .is_wysiwyg = "true";
defparam \plif_exmem.rdat2_l[21] .power_up = "low";
// synopsys translate_on

// Location: FF_X58_Y39_N13
dffeas \plif_exmem.rdat2_l[22] (
	.clk(CPUCLK),
	.d(rdat222),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(exmem_en),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(plif_exmemrdat2_l_22),
	.prn(vcc));
// synopsys translate_off
defparam \plif_exmem.rdat2_l[22] .is_wysiwyg = "true";
defparam \plif_exmem.rdat2_l[22] .power_up = "low";
// synopsys translate_on

// Location: FF_X52_Y39_N27
dffeas \plif_exmem.rdat2_l[23] (
	.clk(CPUCLK),
	.d(rdat223),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(exmem_en),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(plif_exmemrdat2_l_23),
	.prn(vcc));
// synopsys translate_off
defparam \plif_exmem.rdat2_l[23] .is_wysiwyg = "true";
defparam \plif_exmem.rdat2_l[23] .power_up = "low";
// synopsys translate_on

// Location: FF_X53_Y35_N19
dffeas \plif_exmem.rdat2_l[24] (
	.clk(CPUCLK),
	.d(rdat224),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(exmem_en),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(plif_exmemrdat2_l_24),
	.prn(vcc));
// synopsys translate_off
defparam \plif_exmem.rdat2_l[24] .is_wysiwyg = "true";
defparam \plif_exmem.rdat2_l[24] .power_up = "low";
// synopsys translate_on

// Location: FF_X54_Y36_N21
dffeas \plif_exmem.rdat2_l[25] (
	.clk(CPUCLK),
	.d(rdat225),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(exmem_en),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(plif_exmemrdat2_l_25),
	.prn(vcc));
// synopsys translate_off
defparam \plif_exmem.rdat2_l[25] .is_wysiwyg = "true";
defparam \plif_exmem.rdat2_l[25] .power_up = "low";
// synopsys translate_on

// Location: FF_X54_Y36_N3
dffeas \plif_exmem.rdat2_l[26] (
	.clk(CPUCLK),
	.d(rdat226),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(exmem_en),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(plif_exmemrdat2_l_26),
	.prn(vcc));
// synopsys translate_off
defparam \plif_exmem.rdat2_l[26] .is_wysiwyg = "true";
defparam \plif_exmem.rdat2_l[26] .power_up = "low";
// synopsys translate_on

// Location: FF_X54_Y36_N5
dffeas \plif_exmem.rdat2_l[27] (
	.clk(CPUCLK),
	.d(rdat227),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(exmem_en),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(plif_exmemrdat2_l_27),
	.prn(vcc));
// synopsys translate_off
defparam \plif_exmem.rdat2_l[27] .is_wysiwyg = "true";
defparam \plif_exmem.rdat2_l[27] .power_up = "low";
// synopsys translate_on

// Location: FF_X57_Y35_N31
dffeas \plif_exmem.rdat2_l[28] (
	.clk(CPUCLK),
	.d(rdat228),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(exmem_en),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(plif_exmemrdat2_l_28),
	.prn(vcc));
// synopsys translate_off
defparam \plif_exmem.rdat2_l[28] .is_wysiwyg = "true";
defparam \plif_exmem.rdat2_l[28] .power_up = "low";
// synopsys translate_on

// Location: FF_X58_Y34_N11
dffeas \plif_exmem.rdat2_l[29] (
	.clk(CPUCLK),
	.d(rdat229),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(exmem_en),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(plif_exmemrdat2_l_29),
	.prn(vcc));
// synopsys translate_off
defparam \plif_exmem.rdat2_l[29] .is_wysiwyg = "true";
defparam \plif_exmem.rdat2_l[29] .power_up = "low";
// synopsys translate_on

// Location: FF_X55_Y42_N27
dffeas \plif_exmem.rdat2_l[30] (
	.clk(CPUCLK),
	.d(rdat230),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(exmem_en),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(plif_exmemrdat2_l_30),
	.prn(vcc));
// synopsys translate_off
defparam \plif_exmem.rdat2_l[30] .is_wysiwyg = "true";
defparam \plif_exmem.rdat2_l[30] .power_up = "low";
// synopsys translate_on

// Location: FF_X55_Y41_N25
dffeas \plif_exmem.rdat2_l[31] (
	.clk(CPUCLK),
	.d(rdat231),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(exmem_en),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(plif_exmemrdat2_l_31),
	.prn(vcc));
// synopsys translate_off
defparam \plif_exmem.rdat2_l[31] .is_wysiwyg = "true";
defparam \plif_exmem.rdat2_l[31] .power_up = "low";
// synopsys translate_on

// Location: FF_X57_Y32_N17
dffeas \plif_exmem.regsrc_l[0] (
	.clk(CPUCLK),
	.d(\plif_exmem.regsrc_l[0]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(exmem_en),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(plif_exmemregsrc_l_0),
	.prn(vcc));
// synopsys translate_off
defparam \plif_exmem.regsrc_l[0] .is_wysiwyg = "true";
defparam \plif_exmem.regsrc_l[0] .power_up = "low";
// synopsys translate_on

// Location: FF_X57_Y35_N7
dffeas \plif_exmem.regsrc_l[1] (
	.clk(CPUCLK),
	.d(gnd),
	.asdata(plif_idexregsrc_l_1),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(exmem_en),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(plif_exmemregsrc_l_1),
	.prn(vcc));
// synopsys translate_off
defparam \plif_exmem.regsrc_l[1] .is_wysiwyg = "true";
defparam \plif_exmem.regsrc_l[1] .power_up = "low";
// synopsys translate_on

// Location: FF_X55_Y31_N27
dffeas \plif_exmem.rtnaddr_l[31] (
	.clk(CPUCLK),
	.d(\plif_exmem.rtnaddr_l[31]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(exmem_en),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(plif_exmemrtnaddr_l_31),
	.prn(vcc));
// synopsys translate_off
defparam \plif_exmem.rtnaddr_l[31] .is_wysiwyg = "true";
defparam \plif_exmem.rtnaddr_l[31] .power_up = "low";
// synopsys translate_on

// Location: FF_X55_Y42_N23
dffeas \plif_exmem.rtnaddr_l[30] (
	.clk(CPUCLK),
	.d(gnd),
	.asdata(plif_idexrtnaddr_l_30),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(exmem_en),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(plif_exmemrtnaddr_l_30),
	.prn(vcc));
// synopsys translate_off
defparam \plif_exmem.rtnaddr_l[30] .is_wysiwyg = "true";
defparam \plif_exmem.rtnaddr_l[30] .power_up = "low";
// synopsys translate_on

// Location: FF_X58_Y31_N5
dffeas \plif_exmem.rtnaddr_l[29] (
	.clk(CPUCLK),
	.d(gnd),
	.asdata(plif_idexrtnaddr_l_29),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(exmem_en),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(plif_exmemrtnaddr_l_29),
	.prn(vcc));
// synopsys translate_off
defparam \plif_exmem.rtnaddr_l[29] .is_wysiwyg = "true";
defparam \plif_exmem.rtnaddr_l[29] .power_up = "low";
// synopsys translate_on

// Location: FF_X58_Y35_N5
dffeas \plif_exmem.rtnaddr_l[28] (
	.clk(CPUCLK),
	.d(gnd),
	.asdata(plif_idexrtnaddr_l_28),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(exmem_en),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(plif_exmemrtnaddr_l_28),
	.prn(vcc));
// synopsys translate_off
defparam \plif_exmem.rtnaddr_l[28] .is_wysiwyg = "true";
defparam \plif_exmem.rtnaddr_l[28] .power_up = "low";
// synopsys translate_on

// Location: FF_X55_Y32_N9
dffeas \plif_exmem.rtnaddr_l[27] (
	.clk(CPUCLK),
	.d(\plif_exmem.rtnaddr_l[27]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(exmem_en),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(plif_exmemrtnaddr_l_27),
	.prn(vcc));
// synopsys translate_off
defparam \plif_exmem.rtnaddr_l[27] .is_wysiwyg = "true";
defparam \plif_exmem.rtnaddr_l[27] .power_up = "low";
// synopsys translate_on

// Location: FF_X55_Y39_N3
dffeas \plif_exmem.rtnaddr_l[26] (
	.clk(CPUCLK),
	.d(gnd),
	.asdata(plif_idexrtnaddr_l_26),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(exmem_en),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(plif_exmemrtnaddr_l_26),
	.prn(vcc));
// synopsys translate_off
defparam \plif_exmem.rtnaddr_l[26] .is_wysiwyg = "true";
defparam \plif_exmem.rtnaddr_l[26] .power_up = "low";
// synopsys translate_on

// Location: FF_X57_Y35_N27
dffeas \plif_exmem.rtnaddr_l[25] (
	.clk(CPUCLK),
	.d(gnd),
	.asdata(plif_idexrtnaddr_l_25),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(exmem_en),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(plif_exmemrtnaddr_l_25),
	.prn(vcc));
// synopsys translate_off
defparam \plif_exmem.rtnaddr_l[25] .is_wysiwyg = "true";
defparam \plif_exmem.rtnaddr_l[25] .power_up = "low";
// synopsys translate_on

// Location: FF_X53_Y32_N15
dffeas \plif_exmem.rtnaddr_l[24] (
	.clk(CPUCLK),
	.d(\plif_exmem.rtnaddr_l[24]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(exmem_en),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(plif_exmemrtnaddr_l_24),
	.prn(vcc));
// synopsys translate_off
defparam \plif_exmem.rtnaddr_l[24] .is_wysiwyg = "true";
defparam \plif_exmem.rtnaddr_l[24] .power_up = "low";
// synopsys translate_on

// Location: FF_X52_Y39_N25
dffeas \plif_exmem.rtnaddr_l[23] (
	.clk(CPUCLK),
	.d(\plif_exmem.rtnaddr_l[23]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(exmem_en),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(plif_exmemrtnaddr_l_23),
	.prn(vcc));
// synopsys translate_off
defparam \plif_exmem.rtnaddr_l[23] .is_wysiwyg = "true";
defparam \plif_exmem.rtnaddr_l[23] .power_up = "low";
// synopsys translate_on

// Location: FF_X58_Y39_N15
dffeas \plif_exmem.rtnaddr_l[22] (
	.clk(CPUCLK),
	.d(gnd),
	.asdata(plif_idexrtnaddr_l_22),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(exmem_en),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(plif_exmemrtnaddr_l_22),
	.prn(vcc));
// synopsys translate_off
defparam \plif_exmem.rtnaddr_l[22] .is_wysiwyg = "true";
defparam \plif_exmem.rtnaddr_l[22] .power_up = "low";
// synopsys translate_on

// Location: FF_X55_Y31_N13
dffeas \plif_exmem.rtnaddr_l[21] (
	.clk(CPUCLK),
	.d(\plif_exmem.rtnaddr_l[21]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(exmem_en),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(plif_exmemrtnaddr_l_21),
	.prn(vcc));
// synopsys translate_off
defparam \plif_exmem.rtnaddr_l[21] .is_wysiwyg = "true";
defparam \plif_exmem.rtnaddr_l[21] .power_up = "low";
// synopsys translate_on

// Location: FF_X53_Y32_N17
dffeas \plif_exmem.rtnaddr_l[20] (
	.clk(CPUCLK),
	.d(\plif_exmem.rtnaddr_l[20]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(exmem_en),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(plif_exmemrtnaddr_l_20),
	.prn(vcc));
// synopsys translate_off
defparam \plif_exmem.rtnaddr_l[20] .is_wysiwyg = "true";
defparam \plif_exmem.rtnaddr_l[20] .power_up = "low";
// synopsys translate_on

// Location: FF_X53_Y30_N5
dffeas \plif_exmem.rtnaddr_l[19] (
	.clk(CPUCLK),
	.d(\plif_exmem.rtnaddr_l[19]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(exmem_en),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(plif_exmemrtnaddr_l_19),
	.prn(vcc));
// synopsys translate_off
defparam \plif_exmem.rtnaddr_l[19] .is_wysiwyg = "true";
defparam \plif_exmem.rtnaddr_l[19] .power_up = "low";
// synopsys translate_on

// Location: FF_X53_Y30_N15
dffeas \plif_exmem.rtnaddr_l[18] (
	.clk(CPUCLK),
	.d(gnd),
	.asdata(plif_idexrtnaddr_l_18),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(exmem_en),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(plif_exmemrtnaddr_l_18),
	.prn(vcc));
// synopsys translate_off
defparam \plif_exmem.rtnaddr_l[18] .is_wysiwyg = "true";
defparam \plif_exmem.rtnaddr_l[18] .power_up = "low";
// synopsys translate_on

// Location: FF_X53_Y30_N9
dffeas \plif_exmem.rtnaddr_l[17] (
	.clk(CPUCLK),
	.d(\plif_exmem.rtnaddr_l[17]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(exmem_en),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(plif_exmemrtnaddr_l_17),
	.prn(vcc));
// synopsys translate_off
defparam \plif_exmem.rtnaddr_l[17] .is_wysiwyg = "true";
defparam \plif_exmem.rtnaddr_l[17] .power_up = "low";
// synopsys translate_on

// Location: FF_X53_Y30_N11
dffeas \plif_exmem.rtnaddr_l[16] (
	.clk(CPUCLK),
	.d(gnd),
	.asdata(plif_idexrtnaddr_l_16),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(exmem_en),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(plif_exmemrtnaddr_l_16),
	.prn(vcc));
// synopsys translate_off
defparam \plif_exmem.rtnaddr_l[16] .is_wysiwyg = "true";
defparam \plif_exmem.rtnaddr_l[16] .power_up = "low";
// synopsys translate_on

// Location: FF_X53_Y30_N13
dffeas \plif_exmem.rtnaddr_l[15] (
	.clk(CPUCLK),
	.d(\plif_exmem.rtnaddr_l[15]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(exmem_en),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(plif_exmemrtnaddr_l_15),
	.prn(vcc));
// synopsys translate_off
defparam \plif_exmem.rtnaddr_l[15] .is_wysiwyg = "true";
defparam \plif_exmem.rtnaddr_l[15] .power_up = "low";
// synopsys translate_on

// Location: FF_X53_Y30_N19
dffeas \plif_exmem.rtnaddr_l[14] (
	.clk(CPUCLK),
	.d(gnd),
	.asdata(plif_idexrtnaddr_l_14),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(exmem_en),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(plif_exmemrtnaddr_l_14),
	.prn(vcc));
// synopsys translate_off
defparam \plif_exmem.rtnaddr_l[14] .is_wysiwyg = "true";
defparam \plif_exmem.rtnaddr_l[14] .power_up = "low";
// synopsys translate_on

// Location: FF_X54_Y31_N19
dffeas \plif_exmem.rtnaddr_l[13] (
	.clk(CPUCLK),
	.d(\plif_exmem.rtnaddr_l[13]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(exmem_en),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(plif_exmemrtnaddr_l_13),
	.prn(vcc));
// synopsys translate_off
defparam \plif_exmem.rtnaddr_l[13] .is_wysiwyg = "true";
defparam \plif_exmem.rtnaddr_l[13] .power_up = "low";
// synopsys translate_on

// Location: FF_X58_Y34_N31
dffeas \plif_exmem.rtnaddr_l[12] (
	.clk(CPUCLK),
	.d(\plif_exmem.rtnaddr_l[12]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(exmem_en),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(plif_exmemrtnaddr_l_12),
	.prn(vcc));
// synopsys translate_off
defparam \plif_exmem.rtnaddr_l[12] .is_wysiwyg = "true";
defparam \plif_exmem.rtnaddr_l[12] .power_up = "low";
// synopsys translate_on

// Location: FF_X54_Y31_N5
dffeas \plif_exmem.rtnaddr_l[11] (
	.clk(CPUCLK),
	.d(\plif_exmem.rtnaddr_l[11]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(exmem_en),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(plif_exmemrtnaddr_l_11),
	.prn(vcc));
// synopsys translate_off
defparam \plif_exmem.rtnaddr_l[11] .is_wysiwyg = "true";
defparam \plif_exmem.rtnaddr_l[11] .power_up = "low";
// synopsys translate_on

// Location: FF_X54_Y31_N23
dffeas \plif_exmem.rtnaddr_l[10] (
	.clk(CPUCLK),
	.d(gnd),
	.asdata(plif_idexrtnaddr_l_10),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(exmem_en),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(plif_exmemrtnaddr_l_10),
	.prn(vcc));
// synopsys translate_off
defparam \plif_exmem.rtnaddr_l[10] .is_wysiwyg = "true";
defparam \plif_exmem.rtnaddr_l[10] .power_up = "low";
// synopsys translate_on

// Location: FF_X54_Y31_N13
dffeas \plif_exmem.rtnaddr_l[9] (
	.clk(CPUCLK),
	.d(\plif_exmem.rtnaddr_l[9]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(exmem_en),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(plif_exmemrtnaddr_l_9),
	.prn(vcc));
// synopsys translate_off
defparam \plif_exmem.rtnaddr_l[9] .is_wysiwyg = "true";
defparam \plif_exmem.rtnaddr_l[9] .power_up = "low";
// synopsys translate_on

// Location: FF_X54_Y31_N27
dffeas \plif_exmem.rtnaddr_l[8] (
	.clk(CPUCLK),
	.d(\plif_exmem.rtnaddr_l[8]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(exmem_en),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(plif_exmemrtnaddr_l_8),
	.prn(vcc));
// synopsys translate_off
defparam \plif_exmem.rtnaddr_l[8] .is_wysiwyg = "true";
defparam \plif_exmem.rtnaddr_l[8] .power_up = "low";
// synopsys translate_on

// Location: FF_X54_Y31_N17
dffeas \plif_exmem.rtnaddr_l[7] (
	.clk(CPUCLK),
	.d(\plif_exmem.rtnaddr_l[7]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(exmem_en),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(plif_exmemrtnaddr_l_7),
	.prn(vcc));
// synopsys translate_off
defparam \plif_exmem.rtnaddr_l[7] .is_wysiwyg = "true";
defparam \plif_exmem.rtnaddr_l[7] .power_up = "low";
// synopsys translate_on

// Location: FF_X56_Y39_N9
dffeas \plif_exmem.rtnaddr_l[6] (
	.clk(CPUCLK),
	.d(gnd),
	.asdata(plif_idexrtnaddr_l_6),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(exmem_en),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(plif_exmemrtnaddr_l_6),
	.prn(vcc));
// synopsys translate_off
defparam \plif_exmem.rtnaddr_l[6] .is_wysiwyg = "true";
defparam \plif_exmem.rtnaddr_l[6] .power_up = "low";
// synopsys translate_on

// Location: FF_X55_Y31_N23
dffeas \plif_exmem.rtnaddr_l[5] (
	.clk(CPUCLK),
	.d(gnd),
	.asdata(plif_idexrtnaddr_l_5),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(exmem_en),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(plif_exmemrtnaddr_l_5),
	.prn(vcc));
// synopsys translate_off
defparam \plif_exmem.rtnaddr_l[5] .is_wysiwyg = "true";
defparam \plif_exmem.rtnaddr_l[5] .power_up = "low";
// synopsys translate_on

// Location: FF_X50_Y41_N5
dffeas \plif_exmem.rtnaddr_l[2] (
	.clk(CPUCLK),
	.d(\plif_exmem.rtnaddr_l[2]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(exmem_en),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(plif_exmemrtnaddr_l_2),
	.prn(vcc));
// synopsys translate_off
defparam \plif_exmem.rtnaddr_l[2] .is_wysiwyg = "true";
defparam \plif_exmem.rtnaddr_l[2] .power_up = "low";
// synopsys translate_on

// Location: FF_X58_Y34_N17
dffeas \plif_exmem.rtnaddr_l[1] (
	.clk(CPUCLK),
	.d(gnd),
	.asdata(plif_idexrtnaddr_l_1),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(exmem_en),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(plif_exmemrtnaddr_l_1),
	.prn(vcc));
// synopsys translate_off
defparam \plif_exmem.rtnaddr_l[1] .is_wysiwyg = "true";
defparam \plif_exmem.rtnaddr_l[1] .power_up = "low";
// synopsys translate_on

// Location: FF_X50_Y41_N3
dffeas \plif_exmem.rtnaddr_l[0] (
	.clk(CPUCLK),
	.d(gnd),
	.asdata(plif_idexrtnaddr_l_0),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(exmem_en),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(plif_exmemrtnaddr_l_0),
	.prn(vcc));
// synopsys translate_off
defparam \plif_exmem.rtnaddr_l[0] .is_wysiwyg = "true";
defparam \plif_exmem.rtnaddr_l[0] .power_up = "low";
// synopsys translate_on

// Location: FF_X50_Y41_N21
dffeas \plif_exmem.rtnaddr_l[4] (
	.clk(CPUCLK),
	.d(\plif_exmem.rtnaddr_l[4]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(exmem_en),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(plif_exmemrtnaddr_l_4),
	.prn(vcc));
// synopsys translate_off
defparam \plif_exmem.rtnaddr_l[4] .is_wysiwyg = "true";
defparam \plif_exmem.rtnaddr_l[4] .power_up = "low";
// synopsys translate_on

// Location: FF_X50_Y41_N31
dffeas \plif_exmem.rtnaddr_l[3] (
	.clk(CPUCLK),
	.d(\plif_exmem.rtnaddr_l[3]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(exmem_en),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(plif_exmemrtnaddr_l_3),
	.prn(vcc));
// synopsys translate_off
defparam \plif_exmem.rtnaddr_l[3] .is_wysiwyg = "true";
defparam \plif_exmem.rtnaddr_l[3] .power_up = "low";
// synopsys translate_on

// Location: FF_X55_Y32_N29
dffeas \plif_exmem.btype_l (
	.clk(CPUCLK),
	.d(gnd),
	.asdata(plif_idexbtype_l),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(exmem_en),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(plif_exmembtype_l),
	.prn(vcc));
// synopsys translate_off
defparam \plif_exmem.btype_l .is_wysiwyg = "true";
defparam \plif_exmem.btype_l .power_up = "low";
// synopsys translate_on

// Location: FF_X53_Y39_N7
dffeas \plif_exmem.zero_l (
	.clk(CPUCLK),
	.d(WideOr1),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(exmem_en),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(plif_exmemzero_l),
	.prn(vcc));
// synopsys translate_off
defparam \plif_exmem.zero_l .is_wysiwyg = "true";
defparam \plif_exmem.zero_l .power_up = "low";
// synopsys translate_on

// Location: FF_X54_Y29_N1
dffeas \plif_exmem.jaddr_l[1] (
	.clk(CPUCLK),
	.d(gnd),
	.asdata(plif_idexjaddr_l_1),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(exmem_en),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(plif_exmemjaddr_l_1),
	.prn(vcc));
// synopsys translate_off
defparam \plif_exmem.jaddr_l[1] .is_wysiwyg = "true";
defparam \plif_exmem.jaddr_l[1] .power_up = "low";
// synopsys translate_on

// Location: FF_X56_Y32_N19
dffeas \plif_exmem.extimm_l[1] (
	.clk(CPUCLK),
	.d(gnd),
	.asdata(plif_idexextimm_l_1),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(exmem_en),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(plif_exmemextimm_l_1),
	.prn(vcc));
// synopsys translate_off
defparam \plif_exmem.extimm_l[1] .is_wysiwyg = "true";
defparam \plif_exmem.extimm_l[1] .power_up = "low";
// synopsys translate_on

// Location: FF_X57_Y29_N27
dffeas \plif_exmem.extimm_l[0] (
	.clk(CPUCLK),
	.d(gnd),
	.asdata(plif_idexextimm_l_0),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(exmem_en),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(plif_exmemextimm_l_0),
	.prn(vcc));
// synopsys translate_off
defparam \plif_exmem.extimm_l[0] .is_wysiwyg = "true";
defparam \plif_exmem.extimm_l[0] .power_up = "low";
// synopsys translate_on

// Location: FF_X52_Y33_N21
dffeas \plif_exmem.jaddr_l[0] (
	.clk(CPUCLK),
	.d(gnd),
	.asdata(plif_idexjaddr_l_0),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(exmem_en),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(plif_exmemjaddr_l_0),
	.prn(vcc));
// synopsys translate_off
defparam \plif_exmem.jaddr_l[0] .is_wysiwyg = "true";
defparam \plif_exmem.jaddr_l[0] .power_up = "low";
// synopsys translate_on

// Location: FF_X59_Y39_N31
dffeas \plif_exmem.jaddr_l[3] (
	.clk(CPUCLK),
	.d(gnd),
	.asdata(plif_idexjaddr_l_3),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(exmem_en),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(plif_exmemjaddr_l_3),
	.prn(vcc));
// synopsys translate_off
defparam \plif_exmem.jaddr_l[3] .is_wysiwyg = "true";
defparam \plif_exmem.jaddr_l[3] .power_up = "low";
// synopsys translate_on

// Location: FF_X53_Y32_N7
dffeas \plif_exmem.extimm_l[3] (
	.clk(CPUCLK),
	.d(\plif_exmem.extimm_l[3]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(exmem_en),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(plif_exmemextimm_l_3),
	.prn(vcc));
// synopsys translate_off
defparam \plif_exmem.extimm_l[3] .is_wysiwyg = "true";
defparam \plif_exmem.extimm_l[3] .power_up = "low";
// synopsys translate_on

// Location: FF_X53_Y32_N9
dffeas \plif_exmem.extimm_l[2] (
	.clk(CPUCLK),
	.d(gnd),
	.asdata(plif_idexextimm_l_2),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(exmem_en),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(plif_exmemextimm_l_2),
	.prn(vcc));
// synopsys translate_off
defparam \plif_exmem.extimm_l[2] .is_wysiwyg = "true";
defparam \plif_exmem.extimm_l[2] .power_up = "low";
// synopsys translate_on

// Location: FF_X50_Y33_N9
dffeas \plif_exmem.jaddr_l[2] (
	.clk(CPUCLK),
	.d(\plif_exmem.jaddr_l[2]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(exmem_en),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(plif_exmemjaddr_l_2),
	.prn(vcc));
// synopsys translate_off
defparam \plif_exmem.jaddr_l[2] .is_wysiwyg = "true";
defparam \plif_exmem.jaddr_l[2] .power_up = "low";
// synopsys translate_on

// Location: FF_X57_Y29_N29
dffeas \plif_exmem.jaddr_l[5] (
	.clk(CPUCLK),
	.d(gnd),
	.asdata(plif_idexjaddr_l_5),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(exmem_en),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(plif_exmemjaddr_l_5),
	.prn(vcc));
// synopsys translate_off
defparam \plif_exmem.jaddr_l[5] .is_wysiwyg = "true";
defparam \plif_exmem.jaddr_l[5] .power_up = "low";
// synopsys translate_on

// Location: FF_X57_Y29_N31
dffeas \plif_exmem.extimm_l[5] (
	.clk(CPUCLK),
	.d(gnd),
	.asdata(plif_idexextimm_l_5),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(exmem_en),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(plif_exmemextimm_l_5),
	.prn(vcc));
// synopsys translate_off
defparam \plif_exmem.extimm_l[5] .is_wysiwyg = "true";
defparam \plif_exmem.extimm_l[5] .power_up = "low";
// synopsys translate_on

// Location: FF_X58_Y41_N31
dffeas \plif_exmem.extimm_l[4] (
	.clk(CPUCLK),
	.d(\plif_exmem.extimm_l[4]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(exmem_en),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(plif_exmemextimm_l_4),
	.prn(vcc));
// synopsys translate_off
defparam \plif_exmem.extimm_l[4] .is_wysiwyg = "true";
defparam \plif_exmem.extimm_l[4] .power_up = "low";
// synopsys translate_on

// Location: FF_X50_Y33_N31
dffeas \plif_exmem.jaddr_l[4] (
	.clk(CPUCLK),
	.d(gnd),
	.asdata(plif_idexjaddr_l_4),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(exmem_en),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(plif_exmemjaddr_l_4),
	.prn(vcc));
// synopsys translate_off
defparam \plif_exmem.jaddr_l[4] .is_wysiwyg = "true";
defparam \plif_exmem.jaddr_l[4] .power_up = "low";
// synopsys translate_on

// Location: FF_X53_Y32_N19
dffeas \plif_exmem.jaddr_l[7] (
	.clk(CPUCLK),
	.d(\plif_exmem.jaddr_l[7]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(exmem_en),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(plif_exmemjaddr_l_7),
	.prn(vcc));
// synopsys translate_off
defparam \plif_exmem.jaddr_l[7] .is_wysiwyg = "true";
defparam \plif_exmem.jaddr_l[7] .power_up = "low";
// synopsys translate_on

// Location: FF_X57_Y29_N13
dffeas \plif_exmem.extimm_l[7] (
	.clk(CPUCLK),
	.d(gnd),
	.asdata(plif_idexextimm_l_7),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(exmem_en),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(plif_exmemextimm_l_7),
	.prn(vcc));
// synopsys translate_off
defparam \plif_exmem.extimm_l[7] .is_wysiwyg = "true";
defparam \plif_exmem.extimm_l[7] .power_up = "low";
// synopsys translate_on

// Location: FF_X53_Y32_N25
dffeas \plif_exmem.extimm_l[6] (
	.clk(CPUCLK),
	.d(gnd),
	.asdata(plif_idexextimm_l_6),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(exmem_en),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(plif_exmemextimm_l_6),
	.prn(vcc));
// synopsys translate_off
defparam \plif_exmem.extimm_l[6] .is_wysiwyg = "true";
defparam \plif_exmem.extimm_l[6] .power_up = "low";
// synopsys translate_on

// Location: FF_X58_Y32_N11
dffeas \plif_exmem.jaddr_l[6] (
	.clk(CPUCLK),
	.d(gnd),
	.asdata(plif_idexjaddr_l_6),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(exmem_en),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(plif_exmemjaddr_l_6),
	.prn(vcc));
// synopsys translate_off
defparam \plif_exmem.jaddr_l[6] .is_wysiwyg = "true";
defparam \plif_exmem.jaddr_l[6] .power_up = "low";
// synopsys translate_on

// Location: FF_X58_Y32_N1
dffeas \plif_exmem.jaddr_l[9] (
	.clk(CPUCLK),
	.d(\plif_exmem.jaddr_l[9]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(exmem_en),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(plif_exmemjaddr_l_9),
	.prn(vcc));
// synopsys translate_off
defparam \plif_exmem.jaddr_l[9] .is_wysiwyg = "true";
defparam \plif_exmem.jaddr_l[9] .power_up = "low";
// synopsys translate_on

// Location: FF_X58_Y32_N31
dffeas \plif_exmem.extimm_l[9] (
	.clk(CPUCLK),
	.d(gnd),
	.asdata(plif_idexextimm_l_9),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(exmem_en),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(plif_exmemextimm_l_9),
	.prn(vcc));
// synopsys translate_off
defparam \plif_exmem.extimm_l[9] .is_wysiwyg = "true";
defparam \plif_exmem.extimm_l[9] .power_up = "low";
// synopsys translate_on

// Location: FF_X58_Y32_N25
dffeas \plif_exmem.extimm_l[8] (
	.clk(CPUCLK),
	.d(gnd),
	.asdata(plif_idexextimm_l_8),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(exmem_en),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(plif_exmemextimm_l_8),
	.prn(vcc));
// synopsys translate_off
defparam \plif_exmem.extimm_l[8] .is_wysiwyg = "true";
defparam \plif_exmem.extimm_l[8] .power_up = "low";
// synopsys translate_on

// Location: FF_X58_Y34_N5
dffeas \plif_exmem.jaddr_l[8] (
	.clk(CPUCLK),
	.d(\plif_exmem.jaddr_l[8]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(exmem_en),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(plif_exmemjaddr_l_8),
	.prn(vcc));
// synopsys translate_off
defparam \plif_exmem.jaddr_l[8] .is_wysiwyg = "true";
defparam \plif_exmem.jaddr_l[8] .power_up = "low";
// synopsys translate_on

// Location: FF_X58_Y32_N19
dffeas \plif_exmem.jaddr_l[11] (
	.clk(CPUCLK),
	.d(\plif_exmem.jaddr_l[11]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(exmem_en),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(plif_exmemjaddr_l_11),
	.prn(vcc));
// synopsys translate_off
defparam \plif_exmem.jaddr_l[11] .is_wysiwyg = "true";
defparam \plif_exmem.jaddr_l[11] .power_up = "low";
// synopsys translate_on

// Location: FF_X58_Y32_N21
dffeas \plif_exmem.extimm_l[11] (
	.clk(CPUCLK),
	.d(gnd),
	.asdata(plif_idexextimm_l_11),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(exmem_en),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(plif_exmemextimm_l_11),
	.prn(vcc));
// synopsys translate_off
defparam \plif_exmem.extimm_l[11] .is_wysiwyg = "true";
defparam \plif_exmem.extimm_l[11] .power_up = "low";
// synopsys translate_on

// Location: FF_X58_Y32_N23
dffeas \plif_exmem.extimm_l[10] (
	.clk(CPUCLK),
	.d(\plif_exmem.extimm_l[10]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(exmem_en),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(plif_exmemextimm_l_10),
	.prn(vcc));
// synopsys translate_off
defparam \plif_exmem.extimm_l[10] .is_wysiwyg = "true";
defparam \plif_exmem.extimm_l[10] .power_up = "low";
// synopsys translate_on

// Location: FF_X50_Y33_N27
dffeas \plif_exmem.jaddr_l[10] (
	.clk(CPUCLK),
	.d(gnd),
	.asdata(plif_idexjaddr_l_10),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(exmem_en),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(plif_exmemjaddr_l_10),
	.prn(vcc));
// synopsys translate_off
defparam \plif_exmem.jaddr_l[10] .is_wysiwyg = "true";
defparam \plif_exmem.jaddr_l[10] .power_up = "low";
// synopsys translate_on

// Location: FF_X58_Y32_N5
dffeas \plif_exmem.jaddr_l[13] (
	.clk(CPUCLK),
	.d(\plif_exmem.jaddr_l[13]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(exmem_en),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(plif_exmemjaddr_l_13),
	.prn(vcc));
// synopsys translate_off
defparam \plif_exmem.jaddr_l[13] .is_wysiwyg = "true";
defparam \plif_exmem.jaddr_l[13] .power_up = "low";
// synopsys translate_on

// Location: FF_X56_Y32_N15
dffeas \plif_exmem.extimm_l[13] (
	.clk(CPUCLK),
	.d(gnd),
	.asdata(plif_idexextimm_l_13),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(exmem_en),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(plif_exmemextimm_l_13),
	.prn(vcc));
// synopsys translate_off
defparam \plif_exmem.extimm_l[13] .is_wysiwyg = "true";
defparam \plif_exmem.extimm_l[13] .power_up = "low";
// synopsys translate_on

// Location: FF_X60_Y31_N1
dffeas \plif_exmem.extimm_l[12] (
	.clk(CPUCLK),
	.d(\plif_exmem.extimm_l[12]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(exmem_en),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(plif_exmemextimm_l_12),
	.prn(vcc));
// synopsys translate_off
defparam \plif_exmem.extimm_l[12] .is_wysiwyg = "true";
defparam \plif_exmem.extimm_l[12] .power_up = "low";
// synopsys translate_on

// Location: FF_X50_Y32_N23
dffeas \plif_exmem.jaddr_l[12] (
	.clk(CPUCLK),
	.d(\plif_exmem.jaddr_l[12]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(exmem_en),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(plif_exmemjaddr_l_12),
	.prn(vcc));
// synopsys translate_off
defparam \plif_exmem.jaddr_l[12] .is_wysiwyg = "true";
defparam \plif_exmem.jaddr_l[12] .power_up = "low";
// synopsys translate_on

// Location: FF_X60_Y31_N3
dffeas \plif_exmem.jaddr_l[15] (
	.clk(CPUCLK),
	.d(\plif_exmem.jaddr_l[15]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(exmem_en),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(plif_exmemjaddr_l_15),
	.prn(vcc));
// synopsys translate_off
defparam \plif_exmem.jaddr_l[15] .is_wysiwyg = "true";
defparam \plif_exmem.jaddr_l[15] .power_up = "low";
// synopsys translate_on

// Location: FF_X60_Y31_N29
dffeas \plif_exmem.extimm_l[15] (
	.clk(CPUCLK),
	.d(\plif_exmem.extimm_l[15]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(exmem_en),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(plif_exmemextimm_l_15),
	.prn(vcc));
// synopsys translate_off
defparam \plif_exmem.extimm_l[15] .is_wysiwyg = "true";
defparam \plif_exmem.extimm_l[15] .power_up = "low";
// synopsys translate_on

// Location: FF_X60_Y31_N11
dffeas \plif_exmem.extimm_l[14] (
	.clk(CPUCLK),
	.d(\plif_exmem.extimm_l[14]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(exmem_en),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(plif_exmemextimm_l_14),
	.prn(vcc));
// synopsys translate_off
defparam \plif_exmem.extimm_l[14] .is_wysiwyg = "true";
defparam \plif_exmem.extimm_l[14] .power_up = "low";
// synopsys translate_on

// Location: FF_X50_Y33_N5
dffeas \plif_exmem.jaddr_l[14] (
	.clk(CPUCLK),
	.d(\plif_exmem.jaddr_l[14]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(exmem_en),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(plif_exmemjaddr_l_14),
	.prn(vcc));
// synopsys translate_off
defparam \plif_exmem.jaddr_l[14] .is_wysiwyg = "true";
defparam \plif_exmem.jaddr_l[14] .power_up = "low";
// synopsys translate_on

// Location: FF_X58_Y31_N11
dffeas \plif_exmem.jaddr_l[17] (
	.clk(CPUCLK),
	.d(\plif_exmem.jaddr_l[17]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(exmem_en),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(plif_exmemjaddr_l_17),
	.prn(vcc));
// synopsys translate_off
defparam \plif_exmem.jaddr_l[17] .is_wysiwyg = "true";
defparam \plif_exmem.jaddr_l[17] .power_up = "low";
// synopsys translate_on

// Location: FF_X55_Y31_N21
dffeas \plif_exmem.extimm_l[17] (
	.clk(CPUCLK),
	.d(gnd),
	.asdata(plif_idexextimm_l_17),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(exmem_en),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(plif_exmemextimm_l_17),
	.prn(vcc));
// synopsys translate_off
defparam \plif_exmem.extimm_l[17] .is_wysiwyg = "true";
defparam \plif_exmem.extimm_l[17] .power_up = "low";
// synopsys translate_on

// Location: FF_X56_Y28_N11
dffeas \plif_exmem.extimm_l[16] (
	.clk(CPUCLK),
	.d(\plif_exmem.extimm_l[16]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(exmem_en),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(plif_exmemextimm_l_16),
	.prn(vcc));
// synopsys translate_off
defparam \plif_exmem.extimm_l[16] .is_wysiwyg = "true";
defparam \plif_exmem.extimm_l[16] .power_up = "low";
// synopsys translate_on

// Location: FF_X50_Y33_N7
dffeas \plif_exmem.jaddr_l[16] (
	.clk(CPUCLK),
	.d(\plif_exmem.jaddr_l[16]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(exmem_en),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(plif_exmemjaddr_l_16),
	.prn(vcc));
// synopsys translate_off
defparam \plif_exmem.jaddr_l[16] .is_wysiwyg = "true";
defparam \plif_exmem.jaddr_l[16] .power_up = "low";
// synopsys translate_on

// Location: FF_X59_Y37_N27
dffeas \plif_exmem.jaddr_l[19] (
	.clk(CPUCLK),
	.d(\plif_exmem.jaddr_l[19]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(exmem_en),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(plif_exmemjaddr_l_19),
	.prn(vcc));
// synopsys translate_off
defparam \plif_exmem.jaddr_l[19] .is_wysiwyg = "true";
defparam \plif_exmem.jaddr_l[19] .power_up = "low";
// synopsys translate_on

// Location: FF_X56_Y31_N17
dffeas \plif_exmem.extimm_l[19] (
	.clk(CPUCLK),
	.d(gnd),
	.asdata(plif_idexextimm_l_19),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(exmem_en),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(plif_exmemextimm_l_19),
	.prn(vcc));
// synopsys translate_off
defparam \plif_exmem.extimm_l[19] .is_wysiwyg = "true";
defparam \plif_exmem.extimm_l[19] .power_up = "low";
// synopsys translate_on

// Location: FF_X55_Y31_N11
dffeas \plif_exmem.extimm_l[18] (
	.clk(CPUCLK),
	.d(\plif_exmem.extimm_l[18]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(exmem_en),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(plif_exmemextimm_l_18),
	.prn(vcc));
// synopsys translate_off
defparam \plif_exmem.extimm_l[18] .is_wysiwyg = "true";
defparam \plif_exmem.extimm_l[18] .power_up = "low";
// synopsys translate_on

// Location: FF_X59_Y37_N17
dffeas \plif_exmem.jaddr_l[18] (
	.clk(CPUCLK),
	.d(gnd),
	.asdata(plif_idexjaddr_l_18),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(exmem_en),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(plif_exmemjaddr_l_18),
	.prn(vcc));
// synopsys translate_off
defparam \plif_exmem.jaddr_l[18] .is_wysiwyg = "true";
defparam \plif_exmem.jaddr_l[18] .power_up = "low";
// synopsys translate_on

// Location: FF_X55_Y31_N17
dffeas \plif_exmem.jaddr_l[21] (
	.clk(CPUCLK),
	.d(\plif_exmem.jaddr_l[21]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(exmem_en),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(plif_exmemjaddr_l_21),
	.prn(vcc));
// synopsys translate_off
defparam \plif_exmem.jaddr_l[21] .is_wysiwyg = "true";
defparam \plif_exmem.jaddr_l[21] .power_up = "low";
// synopsys translate_on

// Location: FF_X57_Y32_N27
dffeas \plif_exmem.extimm_l[21] (
	.clk(CPUCLK),
	.d(\plif_exmem.extimm_l[21]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(exmem_en),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(plif_exmemextimm_l_21),
	.prn(vcc));
// synopsys translate_off
defparam \plif_exmem.extimm_l[21] .is_wysiwyg = "true";
defparam \plif_exmem.extimm_l[21] .power_up = "low";
// synopsys translate_on

// Location: FF_X56_Y31_N11
dffeas \plif_exmem.extimm_l[20] (
	.clk(CPUCLK),
	.d(gnd),
	.asdata(plif_idexextimm_l_20),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(exmem_en),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(plif_exmemextimm_l_20),
	.prn(vcc));
// synopsys translate_off
defparam \plif_exmem.extimm_l[20] .is_wysiwyg = "true";
defparam \plif_exmem.extimm_l[20] .power_up = "low";
// synopsys translate_on

// Location: FF_X59_Y37_N7
dffeas \plif_exmem.jaddr_l[20] (
	.clk(CPUCLK),
	.d(\plif_exmem.jaddr_l[20]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(exmem_en),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(plif_exmemjaddr_l_20),
	.prn(vcc));
// synopsys translate_off
defparam \plif_exmem.jaddr_l[20] .is_wysiwyg = "true";
defparam \plif_exmem.jaddr_l[20] .power_up = "low";
// synopsys translate_on

// Location: FF_X59_Y37_N13
dffeas \plif_exmem.jaddr_l[23] (
	.clk(CPUCLK),
	.d(\plif_exmem.jaddr_l[23]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(exmem_en),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(plif_exmemjaddr_l_23),
	.prn(vcc));
// synopsys translate_off
defparam \plif_exmem.jaddr_l[23] .is_wysiwyg = "true";
defparam \plif_exmem.jaddr_l[23] .power_up = "low";
// synopsys translate_on

// Location: FF_X55_Y31_N3
dffeas \plif_exmem.extimm_l[23] (
	.clk(CPUCLK),
	.d(gnd),
	.asdata(plif_idexextimm_l_23),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(exmem_en),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(plif_exmemextimm_l_23),
	.prn(vcc));
// synopsys translate_off
defparam \plif_exmem.extimm_l[23] .is_wysiwyg = "true";
defparam \plif_exmem.extimm_l[23] .power_up = "low";
// synopsys translate_on

// Location: FF_X55_Y31_N5
dffeas \plif_exmem.extimm_l[22] (
	.clk(CPUCLK),
	.d(\plif_exmem.extimm_l[22]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(exmem_en),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(plif_exmemextimm_l_22),
	.prn(vcc));
// synopsys translate_off
defparam \plif_exmem.extimm_l[22] .is_wysiwyg = "true";
defparam \plif_exmem.extimm_l[22] .power_up = "low";
// synopsys translate_on

// Location: FF_X50_Y33_N29
dffeas \plif_exmem.jaddr_l[22] (
	.clk(CPUCLK),
	.d(\plif_exmem.jaddr_l[22]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(exmem_en),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(plif_exmemjaddr_l_22),
	.prn(vcc));
// synopsys translate_off
defparam \plif_exmem.jaddr_l[22] .is_wysiwyg = "true";
defparam \plif_exmem.jaddr_l[22] .power_up = "low";
// synopsys translate_on

// Location: FF_X55_Y31_N19
dffeas \plif_exmem.jaddr_l[25] (
	.clk(CPUCLK),
	.d(\plif_exmem.jaddr_l[25]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(exmem_en),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(plif_exmemjaddr_l_25),
	.prn(vcc));
// synopsys translate_off
defparam \plif_exmem.jaddr_l[25] .is_wysiwyg = "true";
defparam \plif_exmem.jaddr_l[25] .power_up = "low";
// synopsys translate_on

// Location: FF_X56_Y31_N19
dffeas \plif_exmem.extimm_l[25] (
	.clk(CPUCLK),
	.d(gnd),
	.asdata(plif_idexextimm_l_25),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(exmem_en),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(plif_exmemextimm_l_25),
	.prn(vcc));
// synopsys translate_off
defparam \plif_exmem.extimm_l[25] .is_wysiwyg = "true";
defparam \plif_exmem.extimm_l[25] .power_up = "low";
// synopsys translate_on

// Location: FF_X56_Y28_N1
dffeas \plif_exmem.extimm_l[24] (
	.clk(CPUCLK),
	.d(gnd),
	.asdata(plif_idexextimm_l_24),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(exmem_en),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(plif_exmemextimm_l_24),
	.prn(vcc));
// synopsys translate_off
defparam \plif_exmem.extimm_l[24] .is_wysiwyg = "true";
defparam \plif_exmem.extimm_l[24] .power_up = "low";
// synopsys translate_on

// Location: FF_X59_Y37_N23
dffeas \plif_exmem.jaddr_l[24] (
	.clk(CPUCLK),
	.d(\plif_exmem.jaddr_l[24]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(exmem_en),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(plif_exmemjaddr_l_24),
	.prn(vcc));
// synopsys translate_off
defparam \plif_exmem.jaddr_l[24] .is_wysiwyg = "true";
defparam \plif_exmem.jaddr_l[24] .power_up = "low";
// synopsys translate_on

// Location: FF_X57_Y32_N31
dffeas \plif_exmem.extimm_l[27] (
	.clk(CPUCLK),
	.d(gnd),
	.asdata(plif_idexextimm_l_27),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(exmem_en),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(plif_exmemextimm_l_27),
	.prn(vcc));
// synopsys translate_off
defparam \plif_exmem.extimm_l[27] .is_wysiwyg = "true";
defparam \plif_exmem.extimm_l[27] .power_up = "low";
// synopsys translate_on

// Location: FF_X56_Y28_N27
dffeas \plif_exmem.extimm_l[26] (
	.clk(CPUCLK),
	.d(gnd),
	.asdata(plif_idexextimm_l_26),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(exmem_en),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(plif_exmemextimm_l_26),
	.prn(vcc));
// synopsys translate_off
defparam \plif_exmem.extimm_l[26] .is_wysiwyg = "true";
defparam \plif_exmem.extimm_l[26] .power_up = "low";
// synopsys translate_on

// Location: FF_X57_Y28_N9
dffeas \plif_exmem.extimm_l[29] (
	.clk(CPUCLK),
	.d(gnd),
	.asdata(plif_idexextimm_l_29),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(exmem_en),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(plif_exmemextimm_l_29),
	.prn(vcc));
// synopsys translate_off
defparam \plif_exmem.extimm_l[29] .is_wysiwyg = "true";
defparam \plif_exmem.extimm_l[29] .power_up = "low";
// synopsys translate_on

// Location: FF_X58_Y31_N9
dffeas \plif_exmem.extimm_l[28] (
	.clk(CPUCLK),
	.d(gnd),
	.asdata(plif_idexextimm_l_28),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(exmem_en),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(plif_exmemextimm_l_28),
	.prn(vcc));
// synopsys translate_off
defparam \plif_exmem.extimm_l[28] .is_wysiwyg = "true";
defparam \plif_exmem.extimm_l[28] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X53_Y39_N16
cycloneive_lcell_comb \plif_exmem.porto_l[1]~feeder (
// Equation(s):
// \plif_exmem.porto_l[1]~feeder_combout  = Selector30

	.dataa(gnd),
	.datab(gnd),
	.datac(Selector30),
	.datad(gnd),
	.cin(gnd),
	.combout(\plif_exmem.porto_l[1]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \plif_exmem.porto_l[1]~feeder .lut_mask = 16'hF0F0;
defparam \plif_exmem.porto_l[1]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X50_Y41_N16
cycloneive_lcell_comb \plif_exmem.porto_l[5]~feeder (
// Equation(s):
// \plif_exmem.porto_l[5]~feeder_combout  = Selector26

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(Selector26),
	.cin(gnd),
	.combout(\plif_exmem.porto_l[5]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \plif_exmem.porto_l[5]~feeder .lut_mask = 16'hFF00;
defparam \plif_exmem.porto_l[5]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y42_N0
cycloneive_lcell_comb \plif_exmem.porto_l[7]~feeder (
// Equation(s):
// \plif_exmem.porto_l[7]~feeder_combout  = Selector24

	.dataa(gnd),
	.datab(gnd),
	.datac(Selector24),
	.datad(gnd),
	.cin(gnd),
	.combout(\plif_exmem.porto_l[7]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \plif_exmem.porto_l[7]~feeder .lut_mask = 16'hF0F0;
defparam \plif_exmem.porto_l[7]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y40_N28
cycloneive_lcell_comb \plif_exmem.porto_l[8]~feeder (
// Equation(s):
// \plif_exmem.porto_l[8]~feeder_combout  = Selector23

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(Selector23),
	.cin(gnd),
	.combout(\plif_exmem.porto_l[8]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \plif_exmem.porto_l[8]~feeder .lut_mask = 16'hFF00;
defparam \plif_exmem.porto_l[8]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y37_N16
cycloneive_lcell_comb \plif_exmem.porto_l[11]~feeder (
// Equation(s):
// \plif_exmem.porto_l[11]~feeder_combout  = Selector20

	.dataa(gnd),
	.datab(gnd),
	.datac(Selector20),
	.datad(gnd),
	.cin(gnd),
	.combout(\plif_exmem.porto_l[11]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \plif_exmem.porto_l[11]~feeder .lut_mask = 16'hF0F0;
defparam \plif_exmem.porto_l[11]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y40_N2
cycloneive_lcell_comb \plif_exmem.porto_l[12]~feeder (
// Equation(s):
// \plif_exmem.porto_l[12]~feeder_combout  = Selector19

	.dataa(gnd),
	.datab(gnd),
	.datac(Selector19),
	.datad(gnd),
	.cin(gnd),
	.combout(\plif_exmem.porto_l[12]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \plif_exmem.porto_l[12]~feeder .lut_mask = 16'hF0F0;
defparam \plif_exmem.porto_l[12]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y39_N30
cycloneive_lcell_comb \plif_exmem.porto_l[14]~feeder (
// Equation(s):
// \plif_exmem.porto_l[14]~feeder_combout  = Selector17

	.dataa(gnd),
	.datab(gnd),
	.datac(Selector17),
	.datad(gnd),
	.cin(gnd),
	.combout(\plif_exmem.porto_l[14]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \plif_exmem.porto_l[14]~feeder .lut_mask = 16'hF0F0;
defparam \plif_exmem.porto_l[14]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X52_Y35_N24
cycloneive_lcell_comb \plif_exmem.porto_l[16]~feeder (
// Equation(s):
// \plif_exmem.porto_l[16]~feeder_combout  = Selector15

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(Selector15),
	.cin(gnd),
	.combout(\plif_exmem.porto_l[16]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \plif_exmem.porto_l[16]~feeder .lut_mask = 16'hFF00;
defparam \plif_exmem.porto_l[16]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y42_N20
cycloneive_lcell_comb \plif_exmem.porto_l[21]~feeder (
// Equation(s):
// \plif_exmem.porto_l[21]~feeder_combout  = Selector10

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(Selector10),
	.cin(gnd),
	.combout(\plif_exmem.porto_l[21]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \plif_exmem.porto_l[21]~feeder .lut_mask = 16'hFF00;
defparam \plif_exmem.porto_l[21]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y39_N22
cycloneive_lcell_comb \plif_exmem.porto_l[20]~feeder (
// Equation(s):
// \plif_exmem.porto_l[20]~feeder_combout  = Selector11

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(Selector11),
	.cin(gnd),
	.combout(\plif_exmem.porto_l[20]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \plif_exmem.porto_l[20]~feeder .lut_mask = 16'hFF00;
defparam \plif_exmem.porto_l[20]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y32_N30
cycloneive_lcell_comb \plif_exmem.pcsrc_l[1]~feeder (
// Equation(s):
// \plif_exmem.pcsrc_l[1]~feeder_combout  = plif_idexpcsrc_l_1

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(plif_idexpcsrc_l_1),
	.cin(gnd),
	.combout(\plif_exmem.pcsrc_l[1]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \plif_exmem.pcsrc_l[1]~feeder .lut_mask = 16'hFF00;
defparam \plif_exmem.pcsrc_l[1]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y32_N22
cycloneive_lcell_comb \plif_exmem.pcsrc_l[0]~feeder (
// Equation(s):
// \plif_exmem.pcsrc_l[0]~feeder_combout  = plif_idexpcsrc_l_0

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(plif_idexpcsrc_l_0),
	.cin(gnd),
	.combout(\plif_exmem.pcsrc_l[0]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \plif_exmem.pcsrc_l[0]~feeder .lut_mask = 16'hFF00;
defparam \plif_exmem.pcsrc_l[0]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y32_N16
cycloneive_lcell_comb \plif_exmem.regsrc_l[0]~feeder (
// Equation(s):
// \plif_exmem.regsrc_l[0]~feeder_combout  = plif_idexregsrc_l_0

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(plif_idexregsrc_l_0),
	.cin(gnd),
	.combout(\plif_exmem.regsrc_l[0]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \plif_exmem.regsrc_l[0]~feeder .lut_mask = 16'hFF00;
defparam \plif_exmem.regsrc_l[0]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y31_N26
cycloneive_lcell_comb \plif_exmem.rtnaddr_l[31]~feeder (
// Equation(s):
// \plif_exmem.rtnaddr_l[31]~feeder_combout  = plif_idexrtnaddr_l_31

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(plif_idexrtnaddr_l_31),
	.cin(gnd),
	.combout(\plif_exmem.rtnaddr_l[31]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \plif_exmem.rtnaddr_l[31]~feeder .lut_mask = 16'hFF00;
defparam \plif_exmem.rtnaddr_l[31]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y32_N8
cycloneive_lcell_comb \plif_exmem.rtnaddr_l[27]~feeder (
// Equation(s):
// \plif_exmem.rtnaddr_l[27]~feeder_combout  = plif_idexrtnaddr_l_27

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(plif_idexrtnaddr_l_27),
	.cin(gnd),
	.combout(\plif_exmem.rtnaddr_l[27]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \plif_exmem.rtnaddr_l[27]~feeder .lut_mask = 16'hFF00;
defparam \plif_exmem.rtnaddr_l[27]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y32_N14
cycloneive_lcell_comb \plif_exmem.rtnaddr_l[24]~feeder (
// Equation(s):
// \plif_exmem.rtnaddr_l[24]~feeder_combout  = plif_idexrtnaddr_l_24

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(plif_idexrtnaddr_l_24),
	.cin(gnd),
	.combout(\plif_exmem.rtnaddr_l[24]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \plif_exmem.rtnaddr_l[24]~feeder .lut_mask = 16'hFF00;
defparam \plif_exmem.rtnaddr_l[24]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X52_Y39_N24
cycloneive_lcell_comb \plif_exmem.rtnaddr_l[23]~feeder (
// Equation(s):
// \plif_exmem.rtnaddr_l[23]~feeder_combout  = plif_idexrtnaddr_l_23

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(plif_idexrtnaddr_l_23),
	.cin(gnd),
	.combout(\plif_exmem.rtnaddr_l[23]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \plif_exmem.rtnaddr_l[23]~feeder .lut_mask = 16'hFF00;
defparam \plif_exmem.rtnaddr_l[23]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y31_N12
cycloneive_lcell_comb \plif_exmem.rtnaddr_l[21]~feeder (
// Equation(s):
// \plif_exmem.rtnaddr_l[21]~feeder_combout  = plif_idexrtnaddr_l_21

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(plif_idexrtnaddr_l_21),
	.cin(gnd),
	.combout(\plif_exmem.rtnaddr_l[21]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \plif_exmem.rtnaddr_l[21]~feeder .lut_mask = 16'hFF00;
defparam \plif_exmem.rtnaddr_l[21]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y32_N16
cycloneive_lcell_comb \plif_exmem.rtnaddr_l[20]~feeder (
// Equation(s):
// \plif_exmem.rtnaddr_l[20]~feeder_combout  = plif_idexrtnaddr_l_20

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(plif_idexrtnaddr_l_20),
	.cin(gnd),
	.combout(\plif_exmem.rtnaddr_l[20]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \plif_exmem.rtnaddr_l[20]~feeder .lut_mask = 16'hFF00;
defparam \plif_exmem.rtnaddr_l[20]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y30_N4
cycloneive_lcell_comb \plif_exmem.rtnaddr_l[19]~feeder (
// Equation(s):
// \plif_exmem.rtnaddr_l[19]~feeder_combout  = plif_idexrtnaddr_l_19

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(plif_idexrtnaddr_l_19),
	.cin(gnd),
	.combout(\plif_exmem.rtnaddr_l[19]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \plif_exmem.rtnaddr_l[19]~feeder .lut_mask = 16'hFF00;
defparam \plif_exmem.rtnaddr_l[19]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y30_N8
cycloneive_lcell_comb \plif_exmem.rtnaddr_l[17]~feeder (
// Equation(s):
// \plif_exmem.rtnaddr_l[17]~feeder_combout  = plif_idexrtnaddr_l_17

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(plif_idexrtnaddr_l_17),
	.cin(gnd),
	.combout(\plif_exmem.rtnaddr_l[17]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \plif_exmem.rtnaddr_l[17]~feeder .lut_mask = 16'hFF00;
defparam \plif_exmem.rtnaddr_l[17]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y30_N12
cycloneive_lcell_comb \plif_exmem.rtnaddr_l[15]~feeder (
// Equation(s):
// \plif_exmem.rtnaddr_l[15]~feeder_combout  = plif_idexrtnaddr_l_15

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(plif_idexrtnaddr_l_15),
	.cin(gnd),
	.combout(\plif_exmem.rtnaddr_l[15]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \plif_exmem.rtnaddr_l[15]~feeder .lut_mask = 16'hFF00;
defparam \plif_exmem.rtnaddr_l[15]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y31_N18
cycloneive_lcell_comb \plif_exmem.rtnaddr_l[13]~feeder (
// Equation(s):
// \plif_exmem.rtnaddr_l[13]~feeder_combout  = plif_idexrtnaddr_l_13

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(plif_idexrtnaddr_l_13),
	.cin(gnd),
	.combout(\plif_exmem.rtnaddr_l[13]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \plif_exmem.rtnaddr_l[13]~feeder .lut_mask = 16'hFF00;
defparam \plif_exmem.rtnaddr_l[13]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y34_N30
cycloneive_lcell_comb \plif_exmem.rtnaddr_l[12]~feeder (
// Equation(s):
// \plif_exmem.rtnaddr_l[12]~feeder_combout  = plif_idexrtnaddr_l_12

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(plif_idexrtnaddr_l_12),
	.cin(gnd),
	.combout(\plif_exmem.rtnaddr_l[12]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \plif_exmem.rtnaddr_l[12]~feeder .lut_mask = 16'hFF00;
defparam \plif_exmem.rtnaddr_l[12]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y31_N4
cycloneive_lcell_comb \plif_exmem.rtnaddr_l[11]~feeder (
// Equation(s):
// \plif_exmem.rtnaddr_l[11]~feeder_combout  = plif_idexrtnaddr_l_11

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(plif_idexrtnaddr_l_11),
	.cin(gnd),
	.combout(\plif_exmem.rtnaddr_l[11]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \plif_exmem.rtnaddr_l[11]~feeder .lut_mask = 16'hFF00;
defparam \plif_exmem.rtnaddr_l[11]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y31_N12
cycloneive_lcell_comb \plif_exmem.rtnaddr_l[9]~feeder (
// Equation(s):
// \plif_exmem.rtnaddr_l[9]~feeder_combout  = plif_idexrtnaddr_l_9

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(plif_idexrtnaddr_l_9),
	.cin(gnd),
	.combout(\plif_exmem.rtnaddr_l[9]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \plif_exmem.rtnaddr_l[9]~feeder .lut_mask = 16'hFF00;
defparam \plif_exmem.rtnaddr_l[9]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y31_N26
cycloneive_lcell_comb \plif_exmem.rtnaddr_l[8]~feeder (
// Equation(s):
// \plif_exmem.rtnaddr_l[8]~feeder_combout  = plif_idexrtnaddr_l_8

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(plif_idexrtnaddr_l_8),
	.cin(gnd),
	.combout(\plif_exmem.rtnaddr_l[8]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \plif_exmem.rtnaddr_l[8]~feeder .lut_mask = 16'hFF00;
defparam \plif_exmem.rtnaddr_l[8]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y31_N16
cycloneive_lcell_comb \plif_exmem.rtnaddr_l[7]~feeder (
// Equation(s):
// \plif_exmem.rtnaddr_l[7]~feeder_combout  = plif_idexrtnaddr_l_7

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(plif_idexrtnaddr_l_7),
	.cin(gnd),
	.combout(\plif_exmem.rtnaddr_l[7]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \plif_exmem.rtnaddr_l[7]~feeder .lut_mask = 16'hFF00;
defparam \plif_exmem.rtnaddr_l[7]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X50_Y41_N4
cycloneive_lcell_comb \plif_exmem.rtnaddr_l[2]~feeder (
// Equation(s):
// \plif_exmem.rtnaddr_l[2]~feeder_combout  = plif_idexrtnaddr_l_2

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(plif_idexrtnaddr_l_2),
	.cin(gnd),
	.combout(\plif_exmem.rtnaddr_l[2]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \plif_exmem.rtnaddr_l[2]~feeder .lut_mask = 16'hFF00;
defparam \plif_exmem.rtnaddr_l[2]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X50_Y41_N20
cycloneive_lcell_comb \plif_exmem.rtnaddr_l[4]~feeder (
// Equation(s):
// \plif_exmem.rtnaddr_l[4]~feeder_combout  = plif_idexrtnaddr_l_4

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(plif_idexrtnaddr_l_4),
	.cin(gnd),
	.combout(\plif_exmem.rtnaddr_l[4]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \plif_exmem.rtnaddr_l[4]~feeder .lut_mask = 16'hFF00;
defparam \plif_exmem.rtnaddr_l[4]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X50_Y41_N30
cycloneive_lcell_comb \plif_exmem.rtnaddr_l[3]~feeder (
// Equation(s):
// \plif_exmem.rtnaddr_l[3]~feeder_combout  = plif_idexrtnaddr_l_3

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(plif_idexrtnaddr_l_3),
	.cin(gnd),
	.combout(\plif_exmem.rtnaddr_l[3]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \plif_exmem.rtnaddr_l[3]~feeder .lut_mask = 16'hFF00;
defparam \plif_exmem.rtnaddr_l[3]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y32_N6
cycloneive_lcell_comb \plif_exmem.extimm_l[3]~feeder (
// Equation(s):
// \plif_exmem.extimm_l[3]~feeder_combout  = plif_idexextimm_l_3

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(plif_idexextimm_l_3),
	.cin(gnd),
	.combout(\plif_exmem.extimm_l[3]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \plif_exmem.extimm_l[3]~feeder .lut_mask = 16'hFF00;
defparam \plif_exmem.extimm_l[3]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X50_Y33_N8
cycloneive_lcell_comb \plif_exmem.jaddr_l[2]~feeder (
// Equation(s):
// \plif_exmem.jaddr_l[2]~feeder_combout  = plif_idexjaddr_l_2

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(plif_idexjaddr_l_2),
	.cin(gnd),
	.combout(\plif_exmem.jaddr_l[2]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \plif_exmem.jaddr_l[2]~feeder .lut_mask = 16'hFF00;
defparam \plif_exmem.jaddr_l[2]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y41_N30
cycloneive_lcell_comb \plif_exmem.extimm_l[4]~feeder (
// Equation(s):
// \plif_exmem.extimm_l[4]~feeder_combout  = plif_idexextimm_l_4

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(plif_idexextimm_l_4),
	.cin(gnd),
	.combout(\plif_exmem.extimm_l[4]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \plif_exmem.extimm_l[4]~feeder .lut_mask = 16'hFF00;
defparam \plif_exmem.extimm_l[4]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y32_N18
cycloneive_lcell_comb \plif_exmem.jaddr_l[7]~feeder (
// Equation(s):
// \plif_exmem.jaddr_l[7]~feeder_combout  = plif_idexjaddr_l_7

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(plif_idexjaddr_l_7),
	.cin(gnd),
	.combout(\plif_exmem.jaddr_l[7]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \plif_exmem.jaddr_l[7]~feeder .lut_mask = 16'hFF00;
defparam \plif_exmem.jaddr_l[7]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y32_N0
cycloneive_lcell_comb \plif_exmem.jaddr_l[9]~feeder (
// Equation(s):
// \plif_exmem.jaddr_l[9]~feeder_combout  = plif_idexjaddr_l_9

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(plif_idexjaddr_l_9),
	.cin(gnd),
	.combout(\plif_exmem.jaddr_l[9]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \plif_exmem.jaddr_l[9]~feeder .lut_mask = 16'hFF00;
defparam \plif_exmem.jaddr_l[9]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y34_N4
cycloneive_lcell_comb \plif_exmem.jaddr_l[8]~feeder (
// Equation(s):
// \plif_exmem.jaddr_l[8]~feeder_combout  = plif_idexjaddr_l_8

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(plif_idexjaddr_l_8),
	.cin(gnd),
	.combout(\plif_exmem.jaddr_l[8]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \plif_exmem.jaddr_l[8]~feeder .lut_mask = 16'hFF00;
defparam \plif_exmem.jaddr_l[8]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y32_N18
cycloneive_lcell_comb \plif_exmem.jaddr_l[11]~feeder (
// Equation(s):
// \plif_exmem.jaddr_l[11]~feeder_combout  = plif_idexjaddr_l_11

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(plif_idexjaddr_l_11),
	.cin(gnd),
	.combout(\plif_exmem.jaddr_l[11]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \plif_exmem.jaddr_l[11]~feeder .lut_mask = 16'hFF00;
defparam \plif_exmem.jaddr_l[11]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y32_N22
cycloneive_lcell_comb \plif_exmem.extimm_l[10]~feeder (
// Equation(s):
// \plif_exmem.extimm_l[10]~feeder_combout  = plif_idexextimm_l_10

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(plif_idexextimm_l_10),
	.cin(gnd),
	.combout(\plif_exmem.extimm_l[10]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \plif_exmem.extimm_l[10]~feeder .lut_mask = 16'hFF00;
defparam \plif_exmem.extimm_l[10]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y32_N4
cycloneive_lcell_comb \plif_exmem.jaddr_l[13]~feeder (
// Equation(s):
// \plif_exmem.jaddr_l[13]~feeder_combout  = plif_idexjaddr_l_13

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(plif_idexjaddr_l_13),
	.cin(gnd),
	.combout(\plif_exmem.jaddr_l[13]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \plif_exmem.jaddr_l[13]~feeder .lut_mask = 16'hFF00;
defparam \plif_exmem.jaddr_l[13]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y31_N0
cycloneive_lcell_comb \plif_exmem.extimm_l[12]~feeder (
// Equation(s):
// \plif_exmem.extimm_l[12]~feeder_combout  = plif_idexextimm_l_12

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(plif_idexextimm_l_12),
	.cin(gnd),
	.combout(\plif_exmem.extimm_l[12]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \plif_exmem.extimm_l[12]~feeder .lut_mask = 16'hFF00;
defparam \plif_exmem.extimm_l[12]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X50_Y32_N22
cycloneive_lcell_comb \plif_exmem.jaddr_l[12]~feeder (
// Equation(s):
// \plif_exmem.jaddr_l[12]~feeder_combout  = plif_idexjaddr_l_12

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(plif_idexjaddr_l_12),
	.cin(gnd),
	.combout(\plif_exmem.jaddr_l[12]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \plif_exmem.jaddr_l[12]~feeder .lut_mask = 16'hFF00;
defparam \plif_exmem.jaddr_l[12]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y31_N2
cycloneive_lcell_comb \plif_exmem.jaddr_l[15]~feeder (
// Equation(s):
// \plif_exmem.jaddr_l[15]~feeder_combout  = plif_idexjaddr_l_15

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(plif_idexjaddr_l_15),
	.cin(gnd),
	.combout(\plif_exmem.jaddr_l[15]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \plif_exmem.jaddr_l[15]~feeder .lut_mask = 16'hFF00;
defparam \plif_exmem.jaddr_l[15]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y31_N28
cycloneive_lcell_comb \plif_exmem.extimm_l[15]~feeder (
// Equation(s):
// \plif_exmem.extimm_l[15]~feeder_combout  = plif_idexextimm_l_15

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(plif_idexextimm_l_15),
	.cin(gnd),
	.combout(\plif_exmem.extimm_l[15]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \plif_exmem.extimm_l[15]~feeder .lut_mask = 16'hFF00;
defparam \plif_exmem.extimm_l[15]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y31_N10
cycloneive_lcell_comb \plif_exmem.extimm_l[14]~feeder (
// Equation(s):
// \plif_exmem.extimm_l[14]~feeder_combout  = plif_idexextimm_l_14

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(plif_idexextimm_l_14),
	.cin(gnd),
	.combout(\plif_exmem.extimm_l[14]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \plif_exmem.extimm_l[14]~feeder .lut_mask = 16'hFF00;
defparam \plif_exmem.extimm_l[14]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X50_Y33_N4
cycloneive_lcell_comb \plif_exmem.jaddr_l[14]~feeder (
// Equation(s):
// \plif_exmem.jaddr_l[14]~feeder_combout  = plif_idexjaddr_l_14

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(plif_idexjaddr_l_14),
	.cin(gnd),
	.combout(\plif_exmem.jaddr_l[14]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \plif_exmem.jaddr_l[14]~feeder .lut_mask = 16'hFF00;
defparam \plif_exmem.jaddr_l[14]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y31_N10
cycloneive_lcell_comb \plif_exmem.jaddr_l[17]~feeder (
// Equation(s):
// \plif_exmem.jaddr_l[17]~feeder_combout  = plif_idexjaddr_l_17

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(plif_idexjaddr_l_17),
	.cin(gnd),
	.combout(\plif_exmem.jaddr_l[17]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \plif_exmem.jaddr_l[17]~feeder .lut_mask = 16'hFF00;
defparam \plif_exmem.jaddr_l[17]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y28_N10
cycloneive_lcell_comb \plif_exmem.extimm_l[16]~feeder (
// Equation(s):
// \plif_exmem.extimm_l[16]~feeder_combout  = plif_idexextimm_l_16

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(plif_idexextimm_l_16),
	.cin(gnd),
	.combout(\plif_exmem.extimm_l[16]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \plif_exmem.extimm_l[16]~feeder .lut_mask = 16'hFF00;
defparam \plif_exmem.extimm_l[16]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X50_Y33_N6
cycloneive_lcell_comb \plif_exmem.jaddr_l[16]~feeder (
// Equation(s):
// \plif_exmem.jaddr_l[16]~feeder_combout  = plif_idexjaddr_l_16

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(plif_idexjaddr_l_16),
	.cin(gnd),
	.combout(\plif_exmem.jaddr_l[16]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \plif_exmem.jaddr_l[16]~feeder .lut_mask = 16'hFF00;
defparam \plif_exmem.jaddr_l[16]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y37_N26
cycloneive_lcell_comb \plif_exmem.jaddr_l[19]~feeder (
// Equation(s):
// \plif_exmem.jaddr_l[19]~feeder_combout  = plif_idexjaddr_l_19

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(plif_idexjaddr_l_19),
	.cin(gnd),
	.combout(\plif_exmem.jaddr_l[19]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \plif_exmem.jaddr_l[19]~feeder .lut_mask = 16'hFF00;
defparam \plif_exmem.jaddr_l[19]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y31_N10
cycloneive_lcell_comb \plif_exmem.extimm_l[18]~feeder (
// Equation(s):
// \plif_exmem.extimm_l[18]~feeder_combout  = plif_idexextimm_l_18

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(plif_idexextimm_l_18),
	.cin(gnd),
	.combout(\plif_exmem.extimm_l[18]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \plif_exmem.extimm_l[18]~feeder .lut_mask = 16'hFF00;
defparam \plif_exmem.extimm_l[18]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y31_N16
cycloneive_lcell_comb \plif_exmem.jaddr_l[21]~feeder (
// Equation(s):
// \plif_exmem.jaddr_l[21]~feeder_combout  = plif_idexjaddr_l_21

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(plif_idexjaddr_l_21),
	.cin(gnd),
	.combout(\plif_exmem.jaddr_l[21]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \plif_exmem.jaddr_l[21]~feeder .lut_mask = 16'hFF00;
defparam \plif_exmem.jaddr_l[21]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y32_N26
cycloneive_lcell_comb \plif_exmem.extimm_l[21]~feeder (
// Equation(s):
// \plif_exmem.extimm_l[21]~feeder_combout  = plif_idexextimm_l_21

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(plif_idexextimm_l_21),
	.cin(gnd),
	.combout(\plif_exmem.extimm_l[21]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \plif_exmem.extimm_l[21]~feeder .lut_mask = 16'hFF00;
defparam \plif_exmem.extimm_l[21]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y37_N6
cycloneive_lcell_comb \plif_exmem.jaddr_l[20]~feeder (
// Equation(s):
// \plif_exmem.jaddr_l[20]~feeder_combout  = plif_idexjaddr_l_20

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(plif_idexjaddr_l_20),
	.cin(gnd),
	.combout(\plif_exmem.jaddr_l[20]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \plif_exmem.jaddr_l[20]~feeder .lut_mask = 16'hFF00;
defparam \plif_exmem.jaddr_l[20]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y37_N12
cycloneive_lcell_comb \plif_exmem.jaddr_l[23]~feeder (
// Equation(s):
// \plif_exmem.jaddr_l[23]~feeder_combout  = plif_idexjaddr_l_23

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(plif_idexjaddr_l_23),
	.cin(gnd),
	.combout(\plif_exmem.jaddr_l[23]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \plif_exmem.jaddr_l[23]~feeder .lut_mask = 16'hFF00;
defparam \plif_exmem.jaddr_l[23]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y31_N4
cycloneive_lcell_comb \plif_exmem.extimm_l[22]~feeder (
// Equation(s):
// \plif_exmem.extimm_l[22]~feeder_combout  = plif_idexextimm_l_22

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(plif_idexextimm_l_22),
	.cin(gnd),
	.combout(\plif_exmem.extimm_l[22]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \plif_exmem.extimm_l[22]~feeder .lut_mask = 16'hFF00;
defparam \plif_exmem.extimm_l[22]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X50_Y33_N28
cycloneive_lcell_comb \plif_exmem.jaddr_l[22]~feeder (
// Equation(s):
// \plif_exmem.jaddr_l[22]~feeder_combout  = plif_idexjaddr_l_22

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(plif_idexjaddr_l_22),
	.cin(gnd),
	.combout(\plif_exmem.jaddr_l[22]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \plif_exmem.jaddr_l[22]~feeder .lut_mask = 16'hFF00;
defparam \plif_exmem.jaddr_l[22]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y31_N18
cycloneive_lcell_comb \plif_exmem.jaddr_l[25]~feeder (
// Equation(s):
// \plif_exmem.jaddr_l[25]~feeder_combout  = plif_idexjaddr_l_25

	.dataa(gnd),
	.datab(gnd),
	.datac(plif_idexjaddr_l_25),
	.datad(gnd),
	.cin(gnd),
	.combout(\plif_exmem.jaddr_l[25]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \plif_exmem.jaddr_l[25]~feeder .lut_mask = 16'hF0F0;
defparam \plif_exmem.jaddr_l[25]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y37_N22
cycloneive_lcell_comb \plif_exmem.jaddr_l[24]~feeder (
// Equation(s):
// \plif_exmem.jaddr_l[24]~feeder_combout  = plif_idexjaddr_l_24

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(plif_idexjaddr_l_24),
	.cin(gnd),
	.combout(\plif_exmem.jaddr_l[24]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \plif_exmem.jaddr_l[24]~feeder .lut_mask = 16'hFF00;
defparam \plif_exmem.jaddr_l[24]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

endmodule

module pipeline_idex (
	plif_exmemdmemWEN_l,
	plif_exmemdmemREN_l,
	always1,
	plif_idexhlt_l,
	plif_memwbpcsrc_l_1,
	plif_memwbpcsrc_l_0,
	plif_idexpcsrc_l_1,
	plif_idexpcsrc_l_0,
	ifid_sRST,
	plif_idexaluop_l_3,
	plif_idexaluop_l_2,
	plif_idexaluop_l_1,
	plif_idexaluop_l_0,
	plif_idexextimm_l_31,
	plif_idexalusrc_l,
	plif_idexrsel2_l_1,
	plif_idexrsel2_l_0,
	plif_idexrsel2_l_2,
	plif_idexrsel2_l_3,
	plif_idexrsel2_l_4,
	plif_idexrdat2_l_31,
	plif_idexextimm_l_30,
	plif_idexrdat2_l_30,
	plif_idexextimm_l_29,
	plif_idexrdat2_l_29,
	plif_idexextimm_l_28,
	plif_idexrdat2_l_28,
	plif_idexextimm_l_27,
	plif_idexrdat2_l_27,
	plif_idexextimm_l_26,
	plif_idexrdat2_l_26,
	plif_idexextimm_l_25,
	plif_idexrdat2_l_25,
	plif_idexextimm_l_24,
	plif_idexrdat2_l_24,
	plif_idexextimm_l_23,
	plif_idexrdat2_l_23,
	plif_idexextimm_l_22,
	plif_idexrdat2_l_22,
	plif_idexextimm_l_21,
	plif_idexrdat2_l_21,
	plif_idexextimm_l_20,
	plif_idexrdat2_l_20,
	plif_idexextimm_l_19,
	plif_idexrdat2_l_19,
	plif_idexextimm_l_18,
	plif_idexrdat2_l_18,
	plif_idexextimm_l_17,
	plif_idexrdat2_l_17,
	plif_idexextimm_l_16,
	plif_idexrdat2_l_16,
	plif_idexextimm_l_15,
	plif_idexrdat2_l_15,
	plif_idexrdat2_l_14,
	plif_idexextimm_l_14,
	plif_idexextimm_l_13,
	plif_idexrdat2_l_13,
	plif_idexrdat2_l_12,
	plif_idexextimm_l_12,
	plif_idexextimm_l_11,
	plif_idexrdat2_l_11,
	plif_idexrdat2_l_10,
	plif_idexextimm_l_10,
	plif_idexextimm_l_9,
	plif_idexrdat2_l_9,
	plif_idexrdat2_l_8,
	plif_idexextimm_l_8,
	plif_idexextimm_l_7,
	plif_idexrdat2_l_7,
	plif_idexrdat2_l_6,
	plif_idexextimm_l_6,
	plif_idexextimm_l_5,
	plif_idexrdat2_l_5,
	plif_idexrsel1_l_4,
	plif_idexrsel1_l_1,
	plif_idexrsel1_l_0,
	plif_idexrsel1_l_2,
	plif_idexrsel1_l_3,
	plif_idexrdat1_l_2,
	plif_idexrdat1_l_1,
	plif_idexrdat2_l_0,
	plif_idexextimm_l_0,
	plif_idexextimm_l_1,
	plif_idexrdat2_l_1,
	plif_idexrdat1_l_4,
	plif_idexrdat1_l_3,
	plif_idexrdat2_l_2,
	plif_idexextimm_l_2,
	plif_idexrdat1_l_8,
	plif_idexrdat1_l_7,
	plif_idexrdat1_l_6,
	plif_idexrdat1_l_5,
	plif_idexextimm_l_3,
	plif_idexrdat2_l_3,
	plif_idexrdat1_l_16,
	plif_idexrdat1_l_15,
	plif_idexrdat1_l_14,
	plif_idexrdat1_l_13,
	plif_idexrdat1_l_12,
	plif_idexrdat1_l_11,
	plif_idexrdat1_l_10,
	plif_idexrdat1_l_9,
	plif_idexrdat2_l_4,
	plif_idexextimm_l_4,
	plif_idexrdat1_l_31,
	plif_idexrdat1_l_29,
	plif_idexrdat1_l_30,
	plif_idexrdat1_l_28,
	plif_idexrdat1_l_27,
	plif_idexrdat1_l_26,
	plif_idexrdat1_l_25,
	plif_idexrdat1_l_24,
	plif_idexrdat1_l_23,
	plif_idexrdat1_l_22,
	plif_idexrdat1_l_21,
	plif_idexrdat1_l_20,
	plif_idexrdat1_l_19,
	plif_idexrdat1_l_18,
	plif_idexrdat1_l_17,
	plif_idexrdat1_l_0,
	plif_idexdmemREN_l,
	plif_idexwsel_l_0,
	plif_idexwsel_l_1,
	plif_ifidinstr_l_31,
	plif_ifidinstr_l_29,
	plif_ifidinstr_l_27,
	plif_ifidinstr_l_26,
	plif_ifidinstr_l_28,
	Equal16,
	plif_ifidinstr_l_30,
	Equal22,
	plif_ifidinstr_l_5,
	plif_ifidinstr_l_1,
	plif_ifidinstr_l_0,
	plif_ifidinstr_l_2,
	plif_ifidinstr_l_3,
	WideNor0,
	Equal11,
	Equal26,
	plif_ifidinstr_l_4,
	Equal21,
	WideOr14,
	Equal13,
	aluop_l,
	WideNor1,
	Selector22,
	Selector4,
	plif_ifidinstr_l_22,
	plif_ifidinstr_l_21,
	plif_idexwsel_l_2,
	plif_idexwsel_l_3,
	plif_ifidinstr_l_24,
	plif_ifidinstr_l_23,
	plif_idexwsel_l_4,
	plif_ifidinstr_l_25,
	Selector1,
	Equal6,
	Selector11,
	Selector21,
	Selector9,
	plif_ifidinstr_l_17,
	plif_ifidinstr_l_16,
	plif_ifidinstr_l_19,
	plif_ifidinstr_l_18,
	plif_ifidinstr_l_20,
	Selector6,
	plif_idexdmemWEN_l,
	Equal23,
	idex_sRST,
	idex_sRST1,
	pcsrc,
	Equal1,
	Equal20,
	WideNor11,
	Equal19,
	Equal12,
	Equal18,
	Selector221,
	plif_ifidinstr_l_15,
	WideOr141,
	WideOr15,
	WideOr16,
	plif_idexregen_l,
	Mux32,
	Mux321,
	extimm_30,
	plif_ifidinstr_l_14,
	Equal0,
	Mux33,
	Mux331,
	plif_ifidinstr_l_13,
	Mux34,
	Mux341,
	plif_ifidinstr_l_12,
	Mux35,
	Mux351,
	plif_ifidinstr_l_11,
	Mux36,
	Mux361,
	plif_ifidinstr_l_10,
	Mux37,
	Mux371,
	plif_ifidinstr_l_9,
	Mux38,
	Mux381,
	plif_ifidinstr_l_8,
	Mux39,
	Mux391,
	plif_ifidinstr_l_7,
	Mux40,
	Mux401,
	plif_ifidinstr_l_6,
	Mux41,
	Mux411,
	Mux42,
	Mux421,
	Selector14,
	Mux43,
	Mux431,
	Selector15,
	Mux44,
	Mux441,
	Selector16,
	Mux45,
	Mux451,
	Selector17,
	Mux46,
	Mux461,
	Selector18,
	Mux47,
	Mux471,
	Mux48,
	Mux481,
	Mux49,
	Mux491,
	Mux50,
	Mux501,
	Mux51,
	Mux511,
	Mux52,
	Mux521,
	Mux53,
	Mux531,
	Mux54,
	Mux541,
	Mux55,
	Mux551,
	Mux56,
	Mux561,
	Mux57,
	Mux571,
	Mux58,
	Mux581,
	Mux29,
	Mux291,
	Mux30,
	Mux301,
	Mux63,
	Mux631,
	Mux62,
	Mux621,
	Mux27,
	Mux271,
	Mux28,
	Mux281,
	Mux61,
	Mux611,
	Mux23,
	Mux231,
	Mux24,
	Mux241,
	Mux25,
	Mux251,
	Mux26,
	Mux261,
	Mux60,
	Mux601,
	Mux15,
	Mux151,
	Mux16,
	Mux161,
	Mux17,
	Mux171,
	Mux18,
	Mux181,
	Mux19,
	Mux191,
	Mux20,
	Mux201,
	Mux21,
	Mux211,
	Mux22,
	Mux221,
	Mux59,
	Mux591,
	Mux0,
	Mux01,
	Mux2,
	Mux210,
	Mux1,
	Mux11,
	Mux3,
	Mux31,
	Mux4,
	Mux410,
	Mux5,
	Mux510,
	Mux6,
	Mux64,
	Mux7,
	Mux71,
	Mux8,
	Mux81,
	Mux9,
	Mux91,
	Mux10,
	Mux101,
	Mux111,
	Mux112,
	Mux12,
	Mux121,
	Mux13,
	Mux131,
	Mux14,
	Mux141,
	Mux311,
	Mux312,
	Selector24,
	plif_idexregsrc_l_0,
	plif_idexregsrc_l_1,
	plif_idexrtnaddr_l_31,
	plif_idexrtnaddr_l_30,
	plif_idexrtnaddr_l_29,
	plif_idexrtnaddr_l_28,
	plif_idexrtnaddr_l_27,
	plif_idexrtnaddr_l_26,
	plif_idexrtnaddr_l_25,
	plif_idexrtnaddr_l_24,
	plif_idexrtnaddr_l_23,
	plif_idexrtnaddr_l_22,
	plif_idexrtnaddr_l_21,
	plif_idexrtnaddr_l_20,
	plif_idexrtnaddr_l_19,
	plif_idexrtnaddr_l_18,
	plif_idexrtnaddr_l_17,
	plif_idexrtnaddr_l_16,
	plif_idexrtnaddr_l_15,
	plif_idexrtnaddr_l_14,
	plif_idexrtnaddr_l_13,
	plif_idexrtnaddr_l_12,
	plif_idexrtnaddr_l_11,
	plif_idexrtnaddr_l_10,
	plif_idexrtnaddr_l_9,
	plif_idexrtnaddr_l_8,
	plif_idexrtnaddr_l_7,
	plif_idexrtnaddr_l_6,
	plif_idexrtnaddr_l_5,
	plif_idexrtnaddr_l_2,
	plif_idexrtnaddr_l_1,
	plif_idexrtnaddr_l_0,
	plif_idexrtnaddr_l_4,
	plif_idexrtnaddr_l_3,
	plif_idexbtype_l,
	plif_idexjaddr_l_1,
	plif_idexjaddr_l_0,
	plif_idexjaddr_l_3,
	plif_idexjaddr_l_2,
	plif_idexjaddr_l_5,
	plif_idexjaddr_l_4,
	plif_idexjaddr_l_7,
	plif_idexjaddr_l_6,
	plif_idexjaddr_l_9,
	plif_idexjaddr_l_8,
	plif_idexjaddr_l_11,
	plif_idexjaddr_l_10,
	plif_idexjaddr_l_13,
	plif_idexjaddr_l_12,
	plif_idexjaddr_l_15,
	plif_idexjaddr_l_14,
	plif_idexjaddr_l_17,
	plif_idexjaddr_l_16,
	plif_idexjaddr_l_19,
	plif_idexjaddr_l_18,
	plif_idexjaddr_l_21,
	plif_idexjaddr_l_20,
	plif_idexjaddr_l_23,
	plif_idexjaddr_l_22,
	plif_idexjaddr_l_25,
	plif_idexjaddr_l_24,
	plif_ifidrtnaddr_l_31,
	plif_ifidrtnaddr_l_30,
	plif_ifidrtnaddr_l_29,
	plif_ifidrtnaddr_l_28,
	plif_ifidrtnaddr_l_27,
	plif_ifidrtnaddr_l_26,
	plif_ifidrtnaddr_l_25,
	plif_ifidrtnaddr_l_24,
	plif_ifidrtnaddr_l_23,
	plif_ifidrtnaddr_l_22,
	plif_ifidrtnaddr_l_21,
	plif_ifidrtnaddr_l_20,
	plif_ifidrtnaddr_l_19,
	plif_ifidrtnaddr_l_18,
	plif_ifidrtnaddr_l_17,
	plif_ifidrtnaddr_l_16,
	plif_ifidrtnaddr_l_15,
	plif_ifidrtnaddr_l_14,
	plif_ifidrtnaddr_l_13,
	plif_ifidrtnaddr_l_12,
	plif_ifidrtnaddr_l_11,
	plif_ifidrtnaddr_l_10,
	plif_ifidrtnaddr_l_9,
	plif_ifidrtnaddr_l_8,
	plif_ifidrtnaddr_l_7,
	plif_ifidrtnaddr_l_6,
	plif_ifidrtnaddr_l_5,
	plif_ifidrtnaddr_l_2,
	plif_ifidrtnaddr_l_1,
	plif_ifidrtnaddr_l_0,
	plif_ifidrtnaddr_l_4,
	plif_ifidrtnaddr_l_3,
	Equal121,
	idex_sRST2,
	Selector0,
	Equal25,
	CPUCLK,
	nRST,
	devpor,
	devclrn,
	devoe);
input 	plif_exmemdmemWEN_l;
input 	plif_exmemdmemREN_l;
input 	always1;
output 	plif_idexhlt_l;
input 	plif_memwbpcsrc_l_1;
input 	plif_memwbpcsrc_l_0;
output 	plif_idexpcsrc_l_1;
output 	plif_idexpcsrc_l_0;
input 	ifid_sRST;
output 	plif_idexaluop_l_3;
output 	plif_idexaluop_l_2;
output 	plif_idexaluop_l_1;
output 	plif_idexaluop_l_0;
output 	plif_idexextimm_l_31;
output 	plif_idexalusrc_l;
output 	plif_idexrsel2_l_1;
output 	plif_idexrsel2_l_0;
output 	plif_idexrsel2_l_2;
output 	plif_idexrsel2_l_3;
output 	plif_idexrsel2_l_4;
output 	plif_idexrdat2_l_31;
output 	plif_idexextimm_l_30;
output 	plif_idexrdat2_l_30;
output 	plif_idexextimm_l_29;
output 	plif_idexrdat2_l_29;
output 	plif_idexextimm_l_28;
output 	plif_idexrdat2_l_28;
output 	plif_idexextimm_l_27;
output 	plif_idexrdat2_l_27;
output 	plif_idexextimm_l_26;
output 	plif_idexrdat2_l_26;
output 	plif_idexextimm_l_25;
output 	plif_idexrdat2_l_25;
output 	plif_idexextimm_l_24;
output 	plif_idexrdat2_l_24;
output 	plif_idexextimm_l_23;
output 	plif_idexrdat2_l_23;
output 	plif_idexextimm_l_22;
output 	plif_idexrdat2_l_22;
output 	plif_idexextimm_l_21;
output 	plif_idexrdat2_l_21;
output 	plif_idexextimm_l_20;
output 	plif_idexrdat2_l_20;
output 	plif_idexextimm_l_19;
output 	plif_idexrdat2_l_19;
output 	plif_idexextimm_l_18;
output 	plif_idexrdat2_l_18;
output 	plif_idexextimm_l_17;
output 	plif_idexrdat2_l_17;
output 	plif_idexextimm_l_16;
output 	plif_idexrdat2_l_16;
output 	plif_idexextimm_l_15;
output 	plif_idexrdat2_l_15;
output 	plif_idexrdat2_l_14;
output 	plif_idexextimm_l_14;
output 	plif_idexextimm_l_13;
output 	plif_idexrdat2_l_13;
output 	plif_idexrdat2_l_12;
output 	plif_idexextimm_l_12;
output 	plif_idexextimm_l_11;
output 	plif_idexrdat2_l_11;
output 	plif_idexrdat2_l_10;
output 	plif_idexextimm_l_10;
output 	plif_idexextimm_l_9;
output 	plif_idexrdat2_l_9;
output 	plif_idexrdat2_l_8;
output 	plif_idexextimm_l_8;
output 	plif_idexextimm_l_7;
output 	plif_idexrdat2_l_7;
output 	plif_idexrdat2_l_6;
output 	plif_idexextimm_l_6;
output 	plif_idexextimm_l_5;
output 	plif_idexrdat2_l_5;
output 	plif_idexrsel1_l_4;
output 	plif_idexrsel1_l_1;
output 	plif_idexrsel1_l_0;
output 	plif_idexrsel1_l_2;
output 	plif_idexrsel1_l_3;
output 	plif_idexrdat1_l_2;
output 	plif_idexrdat1_l_1;
output 	plif_idexrdat2_l_0;
output 	plif_idexextimm_l_0;
output 	plif_idexextimm_l_1;
output 	plif_idexrdat2_l_1;
output 	plif_idexrdat1_l_4;
output 	plif_idexrdat1_l_3;
output 	plif_idexrdat2_l_2;
output 	plif_idexextimm_l_2;
output 	plif_idexrdat1_l_8;
output 	plif_idexrdat1_l_7;
output 	plif_idexrdat1_l_6;
output 	plif_idexrdat1_l_5;
output 	plif_idexextimm_l_3;
output 	plif_idexrdat2_l_3;
output 	plif_idexrdat1_l_16;
output 	plif_idexrdat1_l_15;
output 	plif_idexrdat1_l_14;
output 	plif_idexrdat1_l_13;
output 	plif_idexrdat1_l_12;
output 	plif_idexrdat1_l_11;
output 	plif_idexrdat1_l_10;
output 	plif_idexrdat1_l_9;
output 	plif_idexrdat2_l_4;
output 	plif_idexextimm_l_4;
output 	plif_idexrdat1_l_31;
output 	plif_idexrdat1_l_29;
output 	plif_idexrdat1_l_30;
output 	plif_idexrdat1_l_28;
output 	plif_idexrdat1_l_27;
output 	plif_idexrdat1_l_26;
output 	plif_idexrdat1_l_25;
output 	plif_idexrdat1_l_24;
output 	plif_idexrdat1_l_23;
output 	plif_idexrdat1_l_22;
output 	plif_idexrdat1_l_21;
output 	plif_idexrdat1_l_20;
output 	plif_idexrdat1_l_19;
output 	plif_idexrdat1_l_18;
output 	plif_idexrdat1_l_17;
output 	plif_idexrdat1_l_0;
output 	plif_idexdmemREN_l;
output 	plif_idexwsel_l_0;
output 	plif_idexwsel_l_1;
input 	plif_ifidinstr_l_31;
input 	plif_ifidinstr_l_29;
input 	plif_ifidinstr_l_27;
input 	plif_ifidinstr_l_26;
input 	plif_ifidinstr_l_28;
input 	Equal16;
input 	plif_ifidinstr_l_30;
input 	Equal22;
input 	plif_ifidinstr_l_5;
input 	plif_ifidinstr_l_1;
input 	plif_ifidinstr_l_0;
input 	plif_ifidinstr_l_2;
input 	plif_ifidinstr_l_3;
input 	WideNor0;
input 	Equal11;
input 	Equal26;
input 	plif_ifidinstr_l_4;
input 	Equal21;
input 	WideOr14;
input 	Equal13;
output 	aluop_l;
input 	WideNor1;
input 	Selector22;
input 	Selector4;
input 	plif_ifidinstr_l_22;
input 	plif_ifidinstr_l_21;
output 	plif_idexwsel_l_2;
output 	plif_idexwsel_l_3;
input 	plif_ifidinstr_l_24;
input 	plif_ifidinstr_l_23;
output 	plif_idexwsel_l_4;
input 	plif_ifidinstr_l_25;
input 	Selector1;
input 	Equal6;
input 	Selector11;
input 	Selector21;
input 	Selector9;
input 	plif_ifidinstr_l_17;
input 	plif_ifidinstr_l_16;
input 	plif_ifidinstr_l_19;
input 	plif_ifidinstr_l_18;
input 	plif_ifidinstr_l_20;
input 	Selector6;
output 	plif_idexdmemWEN_l;
input 	Equal23;
input 	idex_sRST;
input 	idex_sRST1;
input 	pcsrc;
input 	Equal1;
input 	Equal20;
input 	WideNor11;
input 	Equal19;
input 	Equal12;
input 	Equal18;
input 	Selector221;
input 	plif_ifidinstr_l_15;
input 	WideOr141;
input 	WideOr15;
input 	WideOr16;
output 	plif_idexregen_l;
input 	Mux32;
input 	Mux321;
input 	extimm_30;
input 	plif_ifidinstr_l_14;
input 	Equal0;
input 	Mux33;
input 	Mux331;
input 	plif_ifidinstr_l_13;
input 	Mux34;
input 	Mux341;
input 	plif_ifidinstr_l_12;
input 	Mux35;
input 	Mux351;
input 	plif_ifidinstr_l_11;
input 	Mux36;
input 	Mux361;
input 	plif_ifidinstr_l_10;
input 	Mux37;
input 	Mux371;
input 	plif_ifidinstr_l_9;
input 	Mux38;
input 	Mux381;
input 	plif_ifidinstr_l_8;
input 	Mux39;
input 	Mux391;
input 	plif_ifidinstr_l_7;
input 	Mux40;
input 	Mux401;
input 	plif_ifidinstr_l_6;
input 	Mux41;
input 	Mux411;
input 	Mux42;
input 	Mux421;
input 	Selector14;
input 	Mux43;
input 	Mux431;
input 	Selector15;
input 	Mux44;
input 	Mux441;
input 	Selector16;
input 	Mux45;
input 	Mux451;
input 	Selector17;
input 	Mux46;
input 	Mux461;
input 	Selector18;
input 	Mux47;
input 	Mux471;
input 	Mux48;
input 	Mux481;
input 	Mux49;
input 	Mux491;
input 	Mux50;
input 	Mux501;
input 	Mux51;
input 	Mux511;
input 	Mux52;
input 	Mux521;
input 	Mux53;
input 	Mux531;
input 	Mux54;
input 	Mux541;
input 	Mux55;
input 	Mux551;
input 	Mux56;
input 	Mux561;
input 	Mux57;
input 	Mux571;
input 	Mux58;
input 	Mux581;
input 	Mux29;
input 	Mux291;
input 	Mux30;
input 	Mux301;
input 	Mux63;
input 	Mux631;
input 	Mux62;
input 	Mux621;
input 	Mux27;
input 	Mux271;
input 	Mux28;
input 	Mux281;
input 	Mux61;
input 	Mux611;
input 	Mux23;
input 	Mux231;
input 	Mux24;
input 	Mux241;
input 	Mux25;
input 	Mux251;
input 	Mux26;
input 	Mux261;
input 	Mux60;
input 	Mux601;
input 	Mux15;
input 	Mux151;
input 	Mux16;
input 	Mux161;
input 	Mux17;
input 	Mux171;
input 	Mux18;
input 	Mux181;
input 	Mux19;
input 	Mux191;
input 	Mux20;
input 	Mux201;
input 	Mux21;
input 	Mux211;
input 	Mux22;
input 	Mux221;
input 	Mux59;
input 	Mux591;
input 	Mux0;
input 	Mux01;
input 	Mux2;
input 	Mux210;
input 	Mux1;
input 	Mux11;
input 	Mux3;
input 	Mux31;
input 	Mux4;
input 	Mux410;
input 	Mux5;
input 	Mux510;
input 	Mux6;
input 	Mux64;
input 	Mux7;
input 	Mux71;
input 	Mux8;
input 	Mux81;
input 	Mux9;
input 	Mux91;
input 	Mux10;
input 	Mux101;
input 	Mux111;
input 	Mux112;
input 	Mux12;
input 	Mux121;
input 	Mux13;
input 	Mux131;
input 	Mux14;
input 	Mux141;
input 	Mux311;
input 	Mux312;
input 	Selector24;
output 	plif_idexregsrc_l_0;
output 	plif_idexregsrc_l_1;
output 	plif_idexrtnaddr_l_31;
output 	plif_idexrtnaddr_l_30;
output 	plif_idexrtnaddr_l_29;
output 	plif_idexrtnaddr_l_28;
output 	plif_idexrtnaddr_l_27;
output 	plif_idexrtnaddr_l_26;
output 	plif_idexrtnaddr_l_25;
output 	plif_idexrtnaddr_l_24;
output 	plif_idexrtnaddr_l_23;
output 	plif_idexrtnaddr_l_22;
output 	plif_idexrtnaddr_l_21;
output 	plif_idexrtnaddr_l_20;
output 	plif_idexrtnaddr_l_19;
output 	plif_idexrtnaddr_l_18;
output 	plif_idexrtnaddr_l_17;
output 	plif_idexrtnaddr_l_16;
output 	plif_idexrtnaddr_l_15;
output 	plif_idexrtnaddr_l_14;
output 	plif_idexrtnaddr_l_13;
output 	plif_idexrtnaddr_l_12;
output 	plif_idexrtnaddr_l_11;
output 	plif_idexrtnaddr_l_10;
output 	plif_idexrtnaddr_l_9;
output 	plif_idexrtnaddr_l_8;
output 	plif_idexrtnaddr_l_7;
output 	plif_idexrtnaddr_l_6;
output 	plif_idexrtnaddr_l_5;
output 	plif_idexrtnaddr_l_2;
output 	plif_idexrtnaddr_l_1;
output 	plif_idexrtnaddr_l_0;
output 	plif_idexrtnaddr_l_4;
output 	plif_idexrtnaddr_l_3;
output 	plif_idexbtype_l;
output 	plif_idexjaddr_l_1;
output 	plif_idexjaddr_l_0;
output 	plif_idexjaddr_l_3;
output 	plif_idexjaddr_l_2;
output 	plif_idexjaddr_l_5;
output 	plif_idexjaddr_l_4;
output 	plif_idexjaddr_l_7;
output 	plif_idexjaddr_l_6;
output 	plif_idexjaddr_l_9;
output 	plif_idexjaddr_l_8;
output 	plif_idexjaddr_l_11;
output 	plif_idexjaddr_l_10;
output 	plif_idexjaddr_l_13;
output 	plif_idexjaddr_l_12;
output 	plif_idexjaddr_l_15;
output 	plif_idexjaddr_l_14;
output 	plif_idexjaddr_l_17;
output 	plif_idexjaddr_l_16;
output 	plif_idexjaddr_l_19;
output 	plif_idexjaddr_l_18;
output 	plif_idexjaddr_l_21;
output 	plif_idexjaddr_l_20;
output 	plif_idexjaddr_l_23;
output 	plif_idexjaddr_l_22;
output 	plif_idexjaddr_l_25;
output 	plif_idexjaddr_l_24;
input 	plif_ifidrtnaddr_l_31;
input 	plif_ifidrtnaddr_l_30;
input 	plif_ifidrtnaddr_l_29;
input 	plif_ifidrtnaddr_l_28;
input 	plif_ifidrtnaddr_l_27;
input 	plif_ifidrtnaddr_l_26;
input 	plif_ifidrtnaddr_l_25;
input 	plif_ifidrtnaddr_l_24;
input 	plif_ifidrtnaddr_l_23;
input 	plif_ifidrtnaddr_l_22;
input 	plif_ifidrtnaddr_l_21;
input 	plif_ifidrtnaddr_l_20;
input 	plif_ifidrtnaddr_l_19;
input 	plif_ifidrtnaddr_l_18;
input 	plif_ifidrtnaddr_l_17;
input 	plif_ifidrtnaddr_l_16;
input 	plif_ifidrtnaddr_l_15;
input 	plif_ifidrtnaddr_l_14;
input 	plif_ifidrtnaddr_l_13;
input 	plif_ifidrtnaddr_l_12;
input 	plif_ifidrtnaddr_l_11;
input 	plif_ifidrtnaddr_l_10;
input 	plif_ifidrtnaddr_l_9;
input 	plif_ifidrtnaddr_l_8;
input 	plif_ifidrtnaddr_l_7;
input 	plif_ifidrtnaddr_l_6;
input 	plif_ifidrtnaddr_l_5;
input 	plif_ifidrtnaddr_l_2;
input 	plif_ifidrtnaddr_l_1;
input 	plif_ifidrtnaddr_l_0;
input 	plif_ifidrtnaddr_l_4;
input 	plif_ifidrtnaddr_l_3;
input 	Equal121;
input 	idex_sRST2;
input 	Selector0;
input 	Equal25;
input 	CPUCLK;
input 	nRST;

// Design Ports Information

input 	devpor;
input 	devclrn;
input 	devoe;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
assign unknown = 1'bx;

wire \hlt_l~0_combout ;
wire \plif_idex.aluop_l[1]~9_combout ;
wire \plif_idex.aluop_l[1]~8_combout ;
wire \pcsrc_l~0_combout ;
wire \pcsrc_l~1_combout ;
wire \pcsrc_l~2_combout ;
wire \aluop_l~2_combout ;
wire \aluop_l~1_combout ;
wire \aluop_l~3_combout ;
wire \aluop_l~4_combout ;
wire \aluop_l~6_combout ;
wire \aluop_l~5_combout ;
wire \aluop_l~7_combout ;
wire \aluop_l~8_combout ;
wire \extimm_l~0_combout ;
wire \extimm_l~1_combout ;
wire \alusrc_l~0_combout ;
wire \rsel2_l~10_combout ;
wire \rsel2_l~11_combout ;
wire \rsel2_l~12_combout ;
wire \rsel2_l~13_combout ;
wire \rsel2_l~14_combout ;
wire \rdat2_l~0_combout ;
wire \extimm_l~2_combout ;
wire \extimm_l~3_combout ;
wire \rdat2_l~1_combout ;
wire \extimm_l~4_combout ;
wire \rdat2_l~2_combout ;
wire \extimm_l~5_combout ;
wire \rdat2_l~3_combout ;
wire \extimm_l~6_combout ;
wire \rdat2_l~4_combout ;
wire \extimm_l~7_combout ;
wire \rdat2_l~5_combout ;
wire \extimm_l~8_combout ;
wire \rdat2_l~6_combout ;
wire \extimm_l~9_combout ;
wire \rdat2_l~7_combout ;
wire \extimm_l~10_combout ;
wire \rdat2_l~8_combout ;
wire \extimm_l~11_combout ;
wire \rdat2_l~9_combout ;
wire \extimm_l~12_combout ;
wire \rdat2_l~10_combout ;
wire \extimm_l~13_combout ;
wire \rdat2_l~11_combout ;
wire \extimm_l~14_combout ;
wire \rdat2_l~12_combout ;
wire \extimm_l~15_combout ;
wire \rdat2_l~13_combout ;
wire \extimm_l~16_combout ;
wire \rdat2_l~14_combout ;
wire \extimm_l~17_combout ;
wire \rdat2_l~15_combout ;
wire \extimm_l~18_combout ;
wire \extimm_l~19_combout ;
wire \rdat2_l~16_combout ;
wire \rdat2_l~17_combout ;
wire \extimm_l~20_combout ;
wire \extimm_l~21_combout ;
wire \rdat2_l~18_combout ;
wire \rdat2_l~19_combout ;
wire \extimm_l~22_combout ;
wire \extimm_l~23_combout ;
wire \rdat2_l~20_combout ;
wire \rdat2_l~21_combout ;
wire \extimm_l~24_combout ;
wire \extimm_l~25_combout ;
wire \rdat2_l~22_combout ;
wire \rdat2_l~23_combout ;
wire \extimm_l~26_combout ;
wire \extimm_l~27_combout ;
wire \rdat2_l~24_combout ;
wire \rdat2_l~25_combout ;
wire \extimm_l~28_combout ;
wire \extimm_l~29_combout ;
wire \rdat2_l~26_combout ;
wire \rsel1_l~10_combout ;
wire \rsel1_l~11_combout ;
wire \rsel1_l~12_combout ;
wire \rsel1_l~13_combout ;
wire \rsel1_l~14_combout ;
wire \rdat1_l~0_combout ;
wire \rdat1_l~1_combout ;
wire \rdat2_l~27_combout ;
wire \extimm_l~30_combout ;
wire \extimm_l~31_combout ;
wire \rdat2_l~28_combout ;
wire \rdat1_l~2_combout ;
wire \rdat1_l~3_combout ;
wire \rdat2_l~29_combout ;
wire \extimm_l~32_combout ;
wire \rdat1_l~4_combout ;
wire \rdat1_l~5_combout ;
wire \rdat1_l~6_combout ;
wire \rdat1_l~7_combout ;
wire \extimm_l~33_combout ;
wire \rdat2_l~30_combout ;
wire \rdat1_l~8_combout ;
wire \rdat1_l~9_combout ;
wire \rdat1_l~10_combout ;
wire \rdat1_l~11_combout ;
wire \rdat1_l~12_combout ;
wire \rdat1_l~13_combout ;
wire \rdat1_l~14_combout ;
wire \rdat1_l~15_combout ;
wire \rdat2_l~31_combout ;
wire \extimm_l~34_combout ;
wire \plif_idex.extimm_l[4]~feeder_combout ;
wire \rdat1_l~16_combout ;
wire \rdat1_l~17_combout ;
wire \rdat1_l~18_combout ;
wire \rdat1_l~19_combout ;
wire \rdat1_l~20_combout ;
wire \rdat1_l~21_combout ;
wire \rdat1_l~22_combout ;
wire \rdat1_l~23_combout ;
wire \rdat1_l~24_combout ;
wire \rdat1_l~25_combout ;
wire \rdat1_l~26_combout ;
wire \rdat1_l~27_combout ;
wire \rdat1_l~28_combout ;
wire \rdat1_l~29_combout ;
wire \rdat1_l~30_combout ;
wire \rdat1_l~31_combout ;
wire \dmemREN_l~0_combout ;
wire \wsel_l~1_combout ;
wire \wsel_l~2_combout ;
wire \wsel_l~0_combout ;
wire \wsel_l~3_combout ;
wire \wsel_l~4_combout ;
wire \wsel_l~5_combout ;
wire \wsel_l~6_combout ;
wire \wsel_l~7_combout ;
wire \wsel_l~8_combout ;
wire \wsel_l~9_combout ;
wire \wsel_l~10_combout ;
wire \dmemWEN_l~0_combout ;
wire \regen_l~0_combout ;
wire \regsrc_l~0_combout ;
wire \regsrc_l~1_combout ;
wire \rtnaddr_l~0_combout ;
wire \rtnaddr_l~1_combout ;
wire \rtnaddr_l~2_combout ;
wire \rtnaddr_l~3_combout ;
wire \rtnaddr_l~4_combout ;
wire \rtnaddr_l~5_combout ;
wire \rtnaddr_l~6_combout ;
wire \rtnaddr_l~7_combout ;
wire \rtnaddr_l~8_combout ;
wire \rtnaddr_l~9_combout ;
wire \rtnaddr_l~10_combout ;
wire \rtnaddr_l~11_combout ;
wire \rtnaddr_l~12_combout ;
wire \rtnaddr_l~13_combout ;
wire \rtnaddr_l~14_combout ;
wire \rtnaddr_l~15_combout ;
wire \rtnaddr_l~16_combout ;
wire \rtnaddr_l~17_combout ;
wire \rtnaddr_l~18_combout ;
wire \rtnaddr_l~19_combout ;
wire \rtnaddr_l~20_combout ;
wire \rtnaddr_l~21_combout ;
wire \rtnaddr_l~22_combout ;
wire \rtnaddr_l~23_combout ;
wire \rtnaddr_l~24_combout ;
wire \rtnaddr_l~25_combout ;
wire \rtnaddr_l~26_combout ;
wire \rtnaddr_l~27_combout ;
wire \rtnaddr_l~28_combout ;
wire \rtnaddr_l~29_combout ;
wire \rtnaddr_l~30_combout ;
wire \rtnaddr_l~31_combout ;
wire \btype_l~0_combout ;
wire \jaddr_l~0_combout ;
wire \jaddr_l~1_combout ;
wire \jaddr_l~2_combout ;
wire \jaddr_l~3_combout ;
wire \jaddr_l~4_combout ;
wire \jaddr_l~5_combout ;
wire \jaddr_l~6_combout ;
wire \jaddr_l~7_combout ;
wire \jaddr_l~8_combout ;
wire \jaddr_l~9_combout ;
wire \jaddr_l~10_combout ;
wire \jaddr_l~11_combout ;
wire \jaddr_l~12_combout ;
wire \jaddr_l~13_combout ;
wire \jaddr_l~14_combout ;
wire \jaddr_l~15_combout ;
wire \jaddr_l~16_combout ;
wire \jaddr_l~17_combout ;
wire \jaddr_l~18_combout ;
wire \jaddr_l~19_combout ;
wire \jaddr_l~20_combout ;
wire \jaddr_l~21_combout ;
wire \jaddr_l~22_combout ;
wire \jaddr_l~23_combout ;
wire \jaddr_l~24_combout ;
wire \jaddr_l~25_combout ;


// Location: FF_X59_Y30_N25
dffeas \plif_idex.hlt_l (
	.clk(CPUCLK),
	.d(\hlt_l~0_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\plif_idex.aluop_l[1]~8_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(plif_idexhlt_l),
	.prn(vcc));
// synopsys translate_off
defparam \plif_idex.hlt_l .is_wysiwyg = "true";
defparam \plif_idex.hlt_l .power_up = "low";
// synopsys translate_on

// Location: FF_X56_Y30_N5
dffeas \plif_idex.pcsrc_l[1] (
	.clk(CPUCLK),
	.d(\pcsrc_l~1_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\plif_idex.aluop_l[1]~8_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(plif_idexpcsrc_l_1),
	.prn(vcc));
// synopsys translate_off
defparam \plif_idex.pcsrc_l[1] .is_wysiwyg = "true";
defparam \plif_idex.pcsrc_l[1] .power_up = "low";
// synopsys translate_on

// Location: FF_X56_Y30_N19
dffeas \plif_idex.pcsrc_l[0] (
	.clk(CPUCLK),
	.d(\pcsrc_l~2_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\plif_idex.aluop_l[1]~8_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(plif_idexpcsrc_l_0),
	.prn(vcc));
// synopsys translate_off
defparam \plif_idex.pcsrc_l[0] .is_wysiwyg = "true";
defparam \plif_idex.pcsrc_l[0] .power_up = "low";
// synopsys translate_on

// Location: FF_X56_Y30_N29
dffeas \plif_idex.aluop_l[3] (
	.clk(CPUCLK),
	.d(\aluop_l~3_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\plif_idex.aluop_l[1]~8_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(plif_idexaluop_l_3),
	.prn(vcc));
// synopsys translate_off
defparam \plif_idex.aluop_l[3] .is_wysiwyg = "true";
defparam \plif_idex.aluop_l[3] .power_up = "low";
// synopsys translate_on

// Location: FF_X56_Y30_N11
dffeas \plif_idex.aluop_l[2] (
	.clk(CPUCLK),
	.d(\aluop_l~4_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\plif_idex.aluop_l[1]~8_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(plif_idexaluop_l_2),
	.prn(vcc));
// synopsys translate_off
defparam \plif_idex.aluop_l[2] .is_wysiwyg = "true";
defparam \plif_idex.aluop_l[2] .power_up = "low";
// synopsys translate_on

// Location: FF_X57_Y33_N17
dffeas \plif_idex.aluop_l[1] (
	.clk(CPUCLK),
	.d(\aluop_l~7_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\plif_idex.aluop_l[1]~8_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(plif_idexaluop_l_1),
	.prn(vcc));
// synopsys translate_off
defparam \plif_idex.aluop_l[1] .is_wysiwyg = "true";
defparam \plif_idex.aluop_l[1] .power_up = "low";
// synopsys translate_on

// Location: FF_X56_Y30_N1
dffeas \plif_idex.aluop_l[0] (
	.clk(CPUCLK),
	.d(\aluop_l~8_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\plif_idex.aluop_l[1]~8_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(plif_idexaluop_l_0),
	.prn(vcc));
// synopsys translate_off
defparam \plif_idex.aluop_l[0] .is_wysiwyg = "true";
defparam \plif_idex.aluop_l[0] .power_up = "low";
// synopsys translate_on

// Location: FF_X58_Y33_N29
dffeas \plif_idex.extimm_l[31] (
	.clk(CPUCLK),
	.d(\extimm_l~1_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\plif_idex.aluop_l[1]~8_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(plif_idexextimm_l_31),
	.prn(vcc));
// synopsys translate_off
defparam \plif_idex.extimm_l[31] .is_wysiwyg = "true";
defparam \plif_idex.extimm_l[31] .power_up = "low";
// synopsys translate_on

// Location: FF_X57_Y33_N11
dffeas \plif_idex.alusrc_l (
	.clk(CPUCLK),
	.d(\alusrc_l~0_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\plif_idex.aluop_l[1]~8_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(plif_idexalusrc_l),
	.prn(vcc));
// synopsys translate_off
defparam \plif_idex.alusrc_l .is_wysiwyg = "true";
defparam \plif_idex.alusrc_l .power_up = "low";
// synopsys translate_on

// Location: FF_X58_Y37_N17
dffeas \plif_idex.rsel2_l[1] (
	.clk(CPUCLK),
	.d(\rsel2_l~10_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\plif_idex.aluop_l[1]~8_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(plif_idexrsel2_l_1),
	.prn(vcc));
// synopsys translate_off
defparam \plif_idex.rsel2_l[1] .is_wysiwyg = "true";
defparam \plif_idex.rsel2_l[1] .power_up = "low";
// synopsys translate_on

// Location: FF_X58_Y37_N7
dffeas \plif_idex.rsel2_l[0] (
	.clk(CPUCLK),
	.d(\rsel2_l~11_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\plif_idex.aluop_l[1]~8_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(plif_idexrsel2_l_0),
	.prn(vcc));
// synopsys translate_off
defparam \plif_idex.rsel2_l[0] .is_wysiwyg = "true";
defparam \plif_idex.rsel2_l[0] .power_up = "low";
// synopsys translate_on

// Location: FF_X58_Y37_N29
dffeas \plif_idex.rsel2_l[2] (
	.clk(CPUCLK),
	.d(\rsel2_l~12_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\plif_idex.aluop_l[1]~8_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(plif_idexrsel2_l_2),
	.prn(vcc));
// synopsys translate_off
defparam \plif_idex.rsel2_l[2] .is_wysiwyg = "true";
defparam \plif_idex.rsel2_l[2] .power_up = "low";
// synopsys translate_on

// Location: FF_X58_Y37_N23
dffeas \plif_idex.rsel2_l[3] (
	.clk(CPUCLK),
	.d(\rsel2_l~13_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\plif_idex.aluop_l[1]~8_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(plif_idexrsel2_l_3),
	.prn(vcc));
// synopsys translate_off
defparam \plif_idex.rsel2_l[3] .is_wysiwyg = "true";
defparam \plif_idex.rsel2_l[3] .power_up = "low";
// synopsys translate_on

// Location: FF_X58_Y37_N25
dffeas \plif_idex.rsel2_l[4] (
	.clk(CPUCLK),
	.d(\rsel2_l~14_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\plif_idex.aluop_l[1]~8_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(plif_idexrsel2_l_4),
	.prn(vcc));
// synopsys translate_off
defparam \plif_idex.rsel2_l[4] .is_wysiwyg = "true";
defparam \plif_idex.rsel2_l[4] .power_up = "low";
// synopsys translate_on

// Location: FF_X67_Y35_N25
dffeas \plif_idex.rdat2_l[31] (
	.clk(CPUCLK),
	.d(\rdat2_l~0_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\plif_idex.aluop_l[1]~8_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(plif_idexrdat2_l_31),
	.prn(vcc));
// synopsys translate_off
defparam \plif_idex.rdat2_l[31] .is_wysiwyg = "true";
defparam \plif_idex.rdat2_l[31] .power_up = "low";
// synopsys translate_on

// Location: FF_X58_Y31_N13
dffeas \plif_idex.extimm_l[30] (
	.clk(CPUCLK),
	.d(\extimm_l~3_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\plif_idex.aluop_l[1]~8_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(plif_idexextimm_l_30),
	.prn(vcc));
// synopsys translate_off
defparam \plif_idex.extimm_l[30] .is_wysiwyg = "true";
defparam \plif_idex.extimm_l[30] .power_up = "low";
// synopsys translate_on

// Location: FF_X61_Y39_N17
dffeas \plif_idex.rdat2_l[30] (
	.clk(CPUCLK),
	.d(\rdat2_l~1_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\plif_idex.aluop_l[1]~8_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(plif_idexrdat2_l_30),
	.prn(vcc));
// synopsys translate_off
defparam \plif_idex.rdat2_l[30] .is_wysiwyg = "true";
defparam \plif_idex.rdat2_l[30] .power_up = "low";
// synopsys translate_on

// Location: FF_X57_Y32_N5
dffeas \plif_idex.extimm_l[29] (
	.clk(CPUCLK),
	.d(\extimm_l~4_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\plif_idex.aluop_l[1]~8_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(plif_idexextimm_l_29),
	.prn(vcc));
// synopsys translate_off
defparam \plif_idex.extimm_l[29] .is_wysiwyg = "true";
defparam \plif_idex.extimm_l[29] .power_up = "low";
// synopsys translate_on

// Location: FF_X61_Y32_N9
dffeas \plif_idex.rdat2_l[29] (
	.clk(CPUCLK),
	.d(\rdat2_l~2_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\plif_idex.aluop_l[1]~8_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(plif_idexrdat2_l_29),
	.prn(vcc));
// synopsys translate_off
defparam \plif_idex.rdat2_l[29] .is_wysiwyg = "true";
defparam \plif_idex.rdat2_l[29] .power_up = "low";
// synopsys translate_on

// Location: FF_X58_Y31_N31
dffeas \plif_idex.extimm_l[28] (
	.clk(CPUCLK),
	.d(\extimm_l~5_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\plif_idex.aluop_l[1]~8_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(plif_idexextimm_l_28),
	.prn(vcc));
// synopsys translate_off
defparam \plif_idex.extimm_l[28] .is_wysiwyg = "true";
defparam \plif_idex.extimm_l[28] .power_up = "low";
// synopsys translate_on

// Location: FF_X67_Y35_N15
dffeas \plif_idex.rdat2_l[28] (
	.clk(CPUCLK),
	.d(\rdat2_l~3_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\plif_idex.aluop_l[1]~8_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(plif_idexrdat2_l_28),
	.prn(vcc));
// synopsys translate_off
defparam \plif_idex.rdat2_l[28] .is_wysiwyg = "true";
defparam \plif_idex.rdat2_l[28] .power_up = "low";
// synopsys translate_on

// Location: FF_X57_Y32_N23
dffeas \plif_idex.extimm_l[27] (
	.clk(CPUCLK),
	.d(\extimm_l~6_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\plif_idex.aluop_l[1]~8_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(plif_idexextimm_l_27),
	.prn(vcc));
// synopsys translate_off
defparam \plif_idex.extimm_l[27] .is_wysiwyg = "true";
defparam \plif_idex.extimm_l[27] .power_up = "low";
// synopsys translate_on

// Location: FF_X61_Y39_N31
dffeas \plif_idex.rdat2_l[27] (
	.clk(CPUCLK),
	.d(\rdat2_l~4_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\plif_idex.aluop_l[1]~8_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(plif_idexrdat2_l_27),
	.prn(vcc));
// synopsys translate_off
defparam \plif_idex.rdat2_l[27] .is_wysiwyg = "true";
defparam \plif_idex.rdat2_l[27] .power_up = "low";
// synopsys translate_on

// Location: FF_X57_Y32_N25
dffeas \plif_idex.extimm_l[26] (
	.clk(CPUCLK),
	.d(\extimm_l~7_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\plif_idex.aluop_l[1]~8_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(plif_idexextimm_l_26),
	.prn(vcc));
// synopsys translate_off
defparam \plif_idex.extimm_l[26] .is_wysiwyg = "true";
defparam \plif_idex.extimm_l[26] .power_up = "low";
// synopsys translate_on

// Location: FF_X61_Y32_N23
dffeas \plif_idex.rdat2_l[26] (
	.clk(CPUCLK),
	.d(\rdat2_l~5_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\plif_idex.aluop_l[1]~8_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(plif_idexrdat2_l_26),
	.prn(vcc));
// synopsys translate_off
defparam \plif_idex.rdat2_l[26] .is_wysiwyg = "true";
defparam \plif_idex.rdat2_l[26] .power_up = "low";
// synopsys translate_on

// Location: FF_X57_Y32_N11
dffeas \plif_idex.extimm_l[25] (
	.clk(CPUCLK),
	.d(\extimm_l~8_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\plif_idex.aluop_l[1]~8_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(plif_idexextimm_l_25),
	.prn(vcc));
// synopsys translate_off
defparam \plif_idex.extimm_l[25] .is_wysiwyg = "true";
defparam \plif_idex.extimm_l[25] .power_up = "low";
// synopsys translate_on

// Location: FF_X65_Y32_N21
dffeas \plif_idex.rdat2_l[25] (
	.clk(CPUCLK),
	.d(\rdat2_l~6_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\plif_idex.aluop_l[1]~8_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(plif_idexrdat2_l_25),
	.prn(vcc));
// synopsys translate_off
defparam \plif_idex.rdat2_l[25] .is_wysiwyg = "true";
defparam \plif_idex.rdat2_l[25] .power_up = "low";
// synopsys translate_on

// Location: FF_X57_Y32_N9
dffeas \plif_idex.extimm_l[24] (
	.clk(CPUCLK),
	.d(\extimm_l~9_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\plif_idex.aluop_l[1]~8_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(plif_idexextimm_l_24),
	.prn(vcc));
// synopsys translate_off
defparam \plif_idex.extimm_l[24] .is_wysiwyg = "true";
defparam \plif_idex.extimm_l[24] .power_up = "low";
// synopsys translate_on

// Location: FF_X65_Y32_N31
dffeas \plif_idex.rdat2_l[24] (
	.clk(CPUCLK),
	.d(\rdat2_l~7_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\plif_idex.aluop_l[1]~8_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(plif_idexrdat2_l_24),
	.prn(vcc));
// synopsys translate_off
defparam \plif_idex.rdat2_l[24] .is_wysiwyg = "true";
defparam \plif_idex.rdat2_l[24] .power_up = "low";
// synopsys translate_on

// Location: FF_X57_Y32_N7
dffeas \plif_idex.extimm_l[23] (
	.clk(CPUCLK),
	.d(\extimm_l~10_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\plif_idex.aluop_l[1]~8_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(plif_idexextimm_l_23),
	.prn(vcc));
// synopsys translate_off
defparam \plif_idex.extimm_l[23] .is_wysiwyg = "true";
defparam \plif_idex.extimm_l[23] .power_up = "low";
// synopsys translate_on

// Location: FF_X67_Y30_N25
dffeas \plif_idex.rdat2_l[23] (
	.clk(CPUCLK),
	.d(\rdat2_l~8_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\plif_idex.aluop_l[1]~8_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(plif_idexrdat2_l_23),
	.prn(vcc));
// synopsys translate_off
defparam \plif_idex.rdat2_l[23] .is_wysiwyg = "true";
defparam \plif_idex.rdat2_l[23] .power_up = "low";
// synopsys translate_on

// Location: FF_X57_Y32_N13
dffeas \plif_idex.extimm_l[22] (
	.clk(CPUCLK),
	.d(\extimm_l~11_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\plif_idex.aluop_l[1]~8_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(plif_idexextimm_l_22),
	.prn(vcc));
// synopsys translate_off
defparam \plif_idex.extimm_l[22] .is_wysiwyg = "true";
defparam \plif_idex.extimm_l[22] .power_up = "low";
// synopsys translate_on

// Location: FF_X67_Y30_N15
dffeas \plif_idex.rdat2_l[22] (
	.clk(CPUCLK),
	.d(\rdat2_l~9_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\plif_idex.aluop_l[1]~8_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(plif_idexrdat2_l_22),
	.prn(vcc));
// synopsys translate_off
defparam \plif_idex.rdat2_l[22] .is_wysiwyg = "true";
defparam \plif_idex.rdat2_l[22] .power_up = "low";
// synopsys translate_on

// Location: FF_X57_Y32_N3
dffeas \plif_idex.extimm_l[21] (
	.clk(CPUCLK),
	.d(\extimm_l~12_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\plif_idex.aluop_l[1]~8_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(plif_idexextimm_l_21),
	.prn(vcc));
// synopsys translate_off
defparam \plif_idex.extimm_l[21] .is_wysiwyg = "true";
defparam \plif_idex.extimm_l[21] .power_up = "low";
// synopsys translate_on

// Location: FF_X67_Y30_N1
dffeas \plif_idex.rdat2_l[21] (
	.clk(CPUCLK),
	.d(\rdat2_l~10_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\plif_idex.aluop_l[1]~8_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(plif_idexrdat2_l_21),
	.prn(vcc));
// synopsys translate_off
defparam \plif_idex.rdat2_l[21] .is_wysiwyg = "true";
defparam \plif_idex.rdat2_l[21] .power_up = "low";
// synopsys translate_on

// Location: FF_X57_Y33_N29
dffeas \plif_idex.extimm_l[20] (
	.clk(CPUCLK),
	.d(\extimm_l~13_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\plif_idex.aluop_l[1]~8_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(plif_idexextimm_l_20),
	.prn(vcc));
// synopsys translate_off
defparam \plif_idex.extimm_l[20] .is_wysiwyg = "true";
defparam \plif_idex.extimm_l[20] .power_up = "low";
// synopsys translate_on

// Location: FF_X60_Y39_N1
dffeas \plif_idex.rdat2_l[20] (
	.clk(CPUCLK),
	.d(\rdat2_l~11_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\plif_idex.aluop_l[1]~8_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(plif_idexrdat2_l_20),
	.prn(vcc));
// synopsys translate_off
defparam \plif_idex.rdat2_l[20] .is_wysiwyg = "true";
defparam \plif_idex.rdat2_l[20] .power_up = "low";
// synopsys translate_on

// Location: FF_X57_Y33_N27
dffeas \plif_idex.extimm_l[19] (
	.clk(CPUCLK),
	.d(\extimm_l~14_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\plif_idex.aluop_l[1]~8_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(plif_idexextimm_l_19),
	.prn(vcc));
// synopsys translate_off
defparam \plif_idex.extimm_l[19] .is_wysiwyg = "true";
defparam \plif_idex.extimm_l[19] .power_up = "low";
// synopsys translate_on

// Location: FF_X60_Y39_N15
dffeas \plif_idex.rdat2_l[19] (
	.clk(CPUCLK),
	.d(\rdat2_l~12_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\plif_idex.aluop_l[1]~8_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(plif_idexrdat2_l_19),
	.prn(vcc));
// synopsys translate_off
defparam \plif_idex.rdat2_l[19] .is_wysiwyg = "true";
defparam \plif_idex.rdat2_l[19] .power_up = "low";
// synopsys translate_on

// Location: FF_X58_Y33_N19
dffeas \plif_idex.extimm_l[18] (
	.clk(CPUCLK),
	.d(\extimm_l~15_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\plif_idex.aluop_l[1]~8_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(plif_idexextimm_l_18),
	.prn(vcc));
// synopsys translate_off
defparam \plif_idex.extimm_l[18] .is_wysiwyg = "true";
defparam \plif_idex.extimm_l[18] .power_up = "low";
// synopsys translate_on

// Location: FF_X63_Y39_N21
dffeas \plif_idex.rdat2_l[18] (
	.clk(CPUCLK),
	.d(\rdat2_l~13_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\plif_idex.aluop_l[1]~8_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(plif_idexrdat2_l_18),
	.prn(vcc));
// synopsys translate_off
defparam \plif_idex.rdat2_l[18] .is_wysiwyg = "true";
defparam \plif_idex.rdat2_l[18] .power_up = "low";
// synopsys translate_on

// Location: FF_X58_Y31_N29
dffeas \plif_idex.extimm_l[17] (
	.clk(CPUCLK),
	.d(\extimm_l~16_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\plif_idex.aluop_l[1]~8_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(plif_idexextimm_l_17),
	.prn(vcc));
// synopsys translate_off
defparam \plif_idex.extimm_l[17] .is_wysiwyg = "true";
defparam \plif_idex.extimm_l[17] .power_up = "low";
// synopsys translate_on

// Location: FF_X67_Y40_N25
dffeas \plif_idex.rdat2_l[17] (
	.clk(CPUCLK),
	.d(\rdat2_l~14_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\plif_idex.aluop_l[1]~8_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(plif_idexrdat2_l_17),
	.prn(vcc));
// synopsys translate_off
defparam \plif_idex.rdat2_l[17] .is_wysiwyg = "true";
defparam \plif_idex.rdat2_l[17] .power_up = "low";
// synopsys translate_on

// Location: FF_X58_Y31_N23
dffeas \plif_idex.extimm_l[16] (
	.clk(CPUCLK),
	.d(\extimm_l~17_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\plif_idex.aluop_l[1]~8_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(plif_idexextimm_l_16),
	.prn(vcc));
// synopsys translate_off
defparam \plif_idex.extimm_l[16] .is_wysiwyg = "true";
defparam \plif_idex.extimm_l[16] .power_up = "low";
// synopsys translate_on

// Location: FF_X67_Y40_N3
dffeas \plif_idex.rdat2_l[16] (
	.clk(CPUCLK),
	.d(\rdat2_l~15_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\plif_idex.aluop_l[1]~8_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(plif_idexrdat2_l_16),
	.prn(vcc));
// synopsys translate_off
defparam \plif_idex.rdat2_l[16] .is_wysiwyg = "true";
defparam \plif_idex.rdat2_l[16] .power_up = "low";
// synopsys translate_on

// Location: FF_X57_Y30_N17
dffeas \plif_idex.extimm_l[15] (
	.clk(CPUCLK),
	.d(\extimm_l~19_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\plif_idex.aluop_l[1]~8_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(plif_idexextimm_l_15),
	.prn(vcc));
// synopsys translate_off
defparam \plif_idex.extimm_l[15] .is_wysiwyg = "true";
defparam \plif_idex.extimm_l[15] .power_up = "low";
// synopsys translate_on

// Location: FF_X70_Y35_N25
dffeas \plif_idex.rdat2_l[15] (
	.clk(CPUCLK),
	.d(\rdat2_l~16_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\plif_idex.aluop_l[1]~8_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(plif_idexrdat2_l_15),
	.prn(vcc));
// synopsys translate_off
defparam \plif_idex.rdat2_l[15] .is_wysiwyg = "true";
defparam \plif_idex.rdat2_l[15] .power_up = "low";
// synopsys translate_on

// Location: FF_X66_Y30_N21
dffeas \plif_idex.rdat2_l[14] (
	.clk(CPUCLK),
	.d(\rdat2_l~17_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\plif_idex.aluop_l[1]~8_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(plif_idexrdat2_l_14),
	.prn(vcc));
// synopsys translate_off
defparam \plif_idex.rdat2_l[14] .is_wysiwyg = "true";
defparam \plif_idex.rdat2_l[14] .power_up = "low";
// synopsys translate_on

// Location: FF_X57_Y30_N15
dffeas \plif_idex.extimm_l[14] (
	.clk(CPUCLK),
	.d(\extimm_l~20_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\plif_idex.aluop_l[1]~8_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(plif_idexextimm_l_14),
	.prn(vcc));
// synopsys translate_off
defparam \plif_idex.extimm_l[14] .is_wysiwyg = "true";
defparam \plif_idex.extimm_l[14] .power_up = "low";
// synopsys translate_on

// Location: FF_X57_Y30_N9
dffeas \plif_idex.extimm_l[13] (
	.clk(CPUCLK),
	.d(\extimm_l~21_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\plif_idex.aluop_l[1]~8_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(plif_idexextimm_l_13),
	.prn(vcc));
// synopsys translate_off
defparam \plif_idex.extimm_l[13] .is_wysiwyg = "true";
defparam \plif_idex.extimm_l[13] .power_up = "low";
// synopsys translate_on

// Location: FF_X57_Y38_N11
dffeas \plif_idex.rdat2_l[13] (
	.clk(CPUCLK),
	.d(\rdat2_l~18_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\plif_idex.aluop_l[1]~8_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(plif_idexrdat2_l_13),
	.prn(vcc));
// synopsys translate_off
defparam \plif_idex.rdat2_l[13] .is_wysiwyg = "true";
defparam \plif_idex.rdat2_l[13] .power_up = "low";
// synopsys translate_on

// Location: FF_X61_Y30_N25
dffeas \plif_idex.rdat2_l[12] (
	.clk(CPUCLK),
	.d(\rdat2_l~19_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\plif_idex.aluop_l[1]~8_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(plif_idexrdat2_l_12),
	.prn(vcc));
// synopsys translate_off
defparam \plif_idex.rdat2_l[12] .is_wysiwyg = "true";
defparam \plif_idex.rdat2_l[12] .power_up = "low";
// synopsys translate_on

// Location: FF_X57_Y30_N19
dffeas \plif_idex.extimm_l[12] (
	.clk(CPUCLK),
	.d(\extimm_l~22_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\plif_idex.aluop_l[1]~8_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(plif_idexextimm_l_12),
	.prn(vcc));
// synopsys translate_off
defparam \plif_idex.extimm_l[12] .is_wysiwyg = "true";
defparam \plif_idex.extimm_l[12] .power_up = "low";
// synopsys translate_on

// Location: FF_X57_Y30_N25
dffeas \plif_idex.extimm_l[11] (
	.clk(CPUCLK),
	.d(\extimm_l~23_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\plif_idex.aluop_l[1]~8_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(plif_idexextimm_l_11),
	.prn(vcc));
// synopsys translate_off
defparam \plif_idex.extimm_l[11] .is_wysiwyg = "true";
defparam \plif_idex.extimm_l[11] .power_up = "low";
// synopsys translate_on

// Location: FF_X58_Y38_N3
dffeas \plif_idex.rdat2_l[11] (
	.clk(CPUCLK),
	.d(\rdat2_l~20_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\plif_idex.aluop_l[1]~8_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(plif_idexrdat2_l_11),
	.prn(vcc));
// synopsys translate_off
defparam \plif_idex.rdat2_l[11] .is_wysiwyg = "true";
defparam \plif_idex.rdat2_l[11] .power_up = "low";
// synopsys translate_on

// Location: FF_X68_Y40_N21
dffeas \plif_idex.rdat2_l[10] (
	.clk(CPUCLK),
	.d(\rdat2_l~21_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\plif_idex.aluop_l[1]~8_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(plif_idexrdat2_l_10),
	.prn(vcc));
// synopsys translate_off
defparam \plif_idex.rdat2_l[10] .is_wysiwyg = "true";
defparam \plif_idex.rdat2_l[10] .power_up = "low";
// synopsys translate_on

// Location: FF_X57_Y30_N7
dffeas \plif_idex.extimm_l[10] (
	.clk(CPUCLK),
	.d(\extimm_l~24_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\plif_idex.aluop_l[1]~8_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(plif_idexextimm_l_10),
	.prn(vcc));
// synopsys translate_off
defparam \plif_idex.extimm_l[10] .is_wysiwyg = "true";
defparam \plif_idex.extimm_l[10] .power_up = "low";
// synopsys translate_on

// Location: FF_X57_Y30_N21
dffeas \plif_idex.extimm_l[9] (
	.clk(CPUCLK),
	.d(\extimm_l~25_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\plif_idex.aluop_l[1]~8_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(plif_idexextimm_l_9),
	.prn(vcc));
// synopsys translate_off
defparam \plif_idex.extimm_l[9] .is_wysiwyg = "true";
defparam \plif_idex.extimm_l[9] .power_up = "low";
// synopsys translate_on

// Location: FF_X68_Y40_N31
dffeas \plif_idex.rdat2_l[9] (
	.clk(CPUCLK),
	.d(\rdat2_l~22_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\plif_idex.aluop_l[1]~8_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(plif_idexrdat2_l_9),
	.prn(vcc));
// synopsys translate_off
defparam \plif_idex.rdat2_l[9] .is_wysiwyg = "true";
defparam \plif_idex.rdat2_l[9] .power_up = "low";
// synopsys translate_on

// Location: FF_X58_Y36_N25
dffeas \plif_idex.rdat2_l[8] (
	.clk(CPUCLK),
	.d(\rdat2_l~23_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\plif_idex.aluop_l[1]~8_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(plif_idexrdat2_l_8),
	.prn(vcc));
// synopsys translate_off
defparam \plif_idex.rdat2_l[8] .is_wysiwyg = "true";
defparam \plif_idex.rdat2_l[8] .power_up = "low";
// synopsys translate_on

// Location: FF_X57_Y30_N23
dffeas \plif_idex.extimm_l[8] (
	.clk(CPUCLK),
	.d(\extimm_l~26_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\plif_idex.aluop_l[1]~8_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(plif_idexextimm_l_8),
	.prn(vcc));
// synopsys translate_off
defparam \plif_idex.extimm_l[8] .is_wysiwyg = "true";
defparam \plif_idex.extimm_l[8] .power_up = "low";
// synopsys translate_on

// Location: FF_X57_Y30_N1
dffeas \plif_idex.extimm_l[7] (
	.clk(CPUCLK),
	.d(\extimm_l~27_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\plif_idex.aluop_l[1]~8_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(plif_idexextimm_l_7),
	.prn(vcc));
// synopsys translate_off
defparam \plif_idex.extimm_l[7] .is_wysiwyg = "true";
defparam \plif_idex.extimm_l[7] .power_up = "low";
// synopsys translate_on

// Location: FF_X56_Y38_N23
dffeas \plif_idex.rdat2_l[7] (
	.clk(CPUCLK),
	.d(\rdat2_l~24_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\plif_idex.aluop_l[1]~8_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(plif_idexrdat2_l_7),
	.prn(vcc));
// synopsys translate_off
defparam \plif_idex.rdat2_l[7] .is_wysiwyg = "true";
defparam \plif_idex.rdat2_l[7] .power_up = "low";
// synopsys translate_on

// Location: FF_X65_Y30_N21
dffeas \plif_idex.rdat2_l[6] (
	.clk(CPUCLK),
	.d(\rdat2_l~25_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\plif_idex.aluop_l[1]~8_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(plif_idexrdat2_l_6),
	.prn(vcc));
// synopsys translate_off
defparam \plif_idex.rdat2_l[6] .is_wysiwyg = "true";
defparam \plif_idex.rdat2_l[6] .power_up = "low";
// synopsys translate_on

// Location: FF_X57_Y30_N3
dffeas \plif_idex.extimm_l[6] (
	.clk(CPUCLK),
	.d(\extimm_l~28_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\plif_idex.aluop_l[1]~8_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(plif_idexextimm_l_6),
	.prn(vcc));
// synopsys translate_off
defparam \plif_idex.extimm_l[6] .is_wysiwyg = "true";
defparam \plif_idex.extimm_l[6] .power_up = "low";
// synopsys translate_on

// Location: FF_X57_Y30_N29
dffeas \plif_idex.extimm_l[5] (
	.clk(CPUCLK),
	.d(\extimm_l~29_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\plif_idex.aluop_l[1]~8_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(plif_idexextimm_l_5),
	.prn(vcc));
// synopsys translate_off
defparam \plif_idex.extimm_l[5] .is_wysiwyg = "true";
defparam \plif_idex.extimm_l[5] .power_up = "low";
// synopsys translate_on

// Location: FF_X65_Y30_N23
dffeas \plif_idex.rdat2_l[5] (
	.clk(CPUCLK),
	.d(\rdat2_l~26_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\plif_idex.aluop_l[1]~8_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(plif_idexrdat2_l_5),
	.prn(vcc));
// synopsys translate_off
defparam \plif_idex.rdat2_l[5] .is_wysiwyg = "true";
defparam \plif_idex.rdat2_l[5] .power_up = "low";
// synopsys translate_on

// Location: FF_X56_Y37_N13
dffeas \plif_idex.rsel1_l[4] (
	.clk(CPUCLK),
	.d(\rsel1_l~10_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\plif_idex.aluop_l[1]~8_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(plif_idexrsel1_l_4),
	.prn(vcc));
// synopsys translate_off
defparam \plif_idex.rsel1_l[4] .is_wysiwyg = "true";
defparam \plif_idex.rsel1_l[4] .power_up = "low";
// synopsys translate_on

// Location: FF_X56_Y37_N9
dffeas \plif_idex.rsel1_l[1] (
	.clk(CPUCLK),
	.d(\rsel1_l~11_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\plif_idex.aluop_l[1]~8_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(plif_idexrsel1_l_1),
	.prn(vcc));
// synopsys translate_off
defparam \plif_idex.rsel1_l[1] .is_wysiwyg = "true";
defparam \plif_idex.rsel1_l[1] .power_up = "low";
// synopsys translate_on

// Location: FF_X56_Y37_N7
dffeas \plif_idex.rsel1_l[0] (
	.clk(CPUCLK),
	.d(\rsel1_l~12_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\plif_idex.aluop_l[1]~8_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(plif_idexrsel1_l_0),
	.prn(vcc));
// synopsys translate_off
defparam \plif_idex.rsel1_l[0] .is_wysiwyg = "true";
defparam \plif_idex.rsel1_l[0] .power_up = "low";
// synopsys translate_on

// Location: FF_X56_Y37_N19
dffeas \plif_idex.rsel1_l[2] (
	.clk(CPUCLK),
	.d(\rsel1_l~13_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\plif_idex.aluop_l[1]~8_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(plif_idexrsel1_l_2),
	.prn(vcc));
// synopsys translate_off
defparam \plif_idex.rsel1_l[2] .is_wysiwyg = "true";
defparam \plif_idex.rsel1_l[2] .power_up = "low";
// synopsys translate_on

// Location: FF_X56_Y37_N25
dffeas \plif_idex.rsel1_l[3] (
	.clk(CPUCLK),
	.d(\rsel1_l~14_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\plif_idex.aluop_l[1]~8_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(plif_idexrsel1_l_3),
	.prn(vcc));
// synopsys translate_off
defparam \plif_idex.rsel1_l[3] .is_wysiwyg = "true";
defparam \plif_idex.rsel1_l[3] .power_up = "low";
// synopsys translate_on

// Location: FF_X63_Y32_N5
dffeas \plif_idex.rdat1_l[2] (
	.clk(CPUCLK),
	.d(\rdat1_l~0_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\plif_idex.aluop_l[1]~8_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(plif_idexrdat1_l_2),
	.prn(vcc));
// synopsys translate_off
defparam \plif_idex.rdat1_l[2] .is_wysiwyg = "true";
defparam \plif_idex.rdat1_l[2] .power_up = "low";
// synopsys translate_on

// Location: FF_X65_Y31_N25
dffeas \plif_idex.rdat1_l[1] (
	.clk(CPUCLK),
	.d(\rdat1_l~1_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\plif_idex.aluop_l[1]~8_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(plif_idexrdat1_l_1),
	.prn(vcc));
// synopsys translate_off
defparam \plif_idex.rdat1_l[1] .is_wysiwyg = "true";
defparam \plif_idex.rdat1_l[1] .power_up = "low";
// synopsys translate_on

// Location: FF_X59_Y35_N25
dffeas \plif_idex.rdat2_l[0] (
	.clk(CPUCLK),
	.d(\rdat2_l~27_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\plif_idex.aluop_l[1]~8_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(plif_idexrdat2_l_0),
	.prn(vcc));
// synopsys translate_off
defparam \plif_idex.rdat2_l[0] .is_wysiwyg = "true";
defparam \plif_idex.rdat2_l[0] .power_up = "low";
// synopsys translate_on

// Location: FF_X58_Y33_N9
dffeas \plif_idex.extimm_l[0] (
	.clk(CPUCLK),
	.d(\extimm_l~30_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\plif_idex.aluop_l[1]~8_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(plif_idexextimm_l_0),
	.prn(vcc));
// synopsys translate_off
defparam \plif_idex.extimm_l[0] .is_wysiwyg = "true";
defparam \plif_idex.extimm_l[0] .power_up = "low";
// synopsys translate_on

// Location: FF_X59_Y37_N21
dffeas \plif_idex.extimm_l[1] (
	.clk(CPUCLK),
	.d(\extimm_l~31_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\plif_idex.aluop_l[1]~8_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(plif_idexextimm_l_1),
	.prn(vcc));
// synopsys translate_off
defparam \plif_idex.extimm_l[1] .is_wysiwyg = "true";
defparam \plif_idex.extimm_l[1] .power_up = "low";
// synopsys translate_on

// Location: FF_X59_Y35_N11
dffeas \plif_idex.rdat2_l[1] (
	.clk(CPUCLK),
	.d(\rdat2_l~28_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\plif_idex.aluop_l[1]~8_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(plif_idexrdat2_l_1),
	.prn(vcc));
// synopsys translate_off
defparam \plif_idex.rdat2_l[1] .is_wysiwyg = "true";
defparam \plif_idex.rdat2_l[1] .power_up = "low";
// synopsys translate_on

// Location: FF_X59_Y34_N1
dffeas \plif_idex.rdat1_l[4] (
	.clk(CPUCLK),
	.d(\rdat1_l~2_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\plif_idex.aluop_l[1]~8_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(plif_idexrdat1_l_4),
	.prn(vcc));
// synopsys translate_off
defparam \plif_idex.rdat1_l[4] .is_wysiwyg = "true";
defparam \plif_idex.rdat1_l[4] .power_up = "low";
// synopsys translate_on

// Location: FF_X70_Y37_N25
dffeas \plif_idex.rdat1_l[3] (
	.clk(CPUCLK),
	.d(\rdat1_l~3_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\plif_idex.aluop_l[1]~8_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(plif_idexrdat1_l_3),
	.prn(vcc));
// synopsys translate_off
defparam \plif_idex.rdat1_l[3] .is_wysiwyg = "true";
defparam \plif_idex.rdat1_l[3] .power_up = "low";
// synopsys translate_on

// Location: FF_X59_Y35_N29
dffeas \plif_idex.rdat2_l[2] (
	.clk(CPUCLK),
	.d(\rdat2_l~29_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\plif_idex.aluop_l[1]~8_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(plif_idexrdat2_l_2),
	.prn(vcc));
// synopsys translate_off
defparam \plif_idex.rdat2_l[2] .is_wysiwyg = "true";
defparam \plif_idex.rdat2_l[2] .power_up = "low";
// synopsys translate_on

// Location: FF_X58_Y36_N11
dffeas \plif_idex.extimm_l[2] (
	.clk(CPUCLK),
	.d(\extimm_l~32_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\plif_idex.aluop_l[1]~8_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(plif_idexextimm_l_2),
	.prn(vcc));
// synopsys translate_off
defparam \plif_idex.extimm_l[2] .is_wysiwyg = "true";
defparam \plif_idex.extimm_l[2] .power_up = "low";
// synopsys translate_on

// Location: FF_X68_Y36_N21
dffeas \plif_idex.rdat1_l[8] (
	.clk(CPUCLK),
	.d(\rdat1_l~4_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\plif_idex.aluop_l[1]~8_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(plif_idexrdat1_l_8),
	.prn(vcc));
// synopsys translate_off
defparam \plif_idex.rdat1_l[8] .is_wysiwyg = "true";
defparam \plif_idex.rdat1_l[8] .power_up = "low";
// synopsys translate_on

// Location: FF_X60_Y40_N29
dffeas \plif_idex.rdat1_l[7] (
	.clk(CPUCLK),
	.d(\rdat1_l~5_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\plif_idex.aluop_l[1]~8_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(plif_idexrdat1_l_7),
	.prn(vcc));
// synopsys translate_off
defparam \plif_idex.rdat1_l[7] .is_wysiwyg = "true";
defparam \plif_idex.rdat1_l[7] .power_up = "low";
// synopsys translate_on

// Location: FF_X67_Y36_N17
dffeas \plif_idex.rdat1_l[6] (
	.clk(CPUCLK),
	.d(\rdat1_l~6_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\plif_idex.aluop_l[1]~8_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(plif_idexrdat1_l_6),
	.prn(vcc));
// synopsys translate_off
defparam \plif_idex.rdat1_l[6] .is_wysiwyg = "true";
defparam \plif_idex.rdat1_l[6] .power_up = "low";
// synopsys translate_on

// Location: FF_X67_Y36_N27
dffeas \plif_idex.rdat1_l[5] (
	.clk(CPUCLK),
	.d(\rdat1_l~7_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\plif_idex.aluop_l[1]~8_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(plif_idexrdat1_l_5),
	.prn(vcc));
// synopsys translate_off
defparam \plif_idex.rdat1_l[5] .is_wysiwyg = "true";
defparam \plif_idex.rdat1_l[5] .power_up = "low";
// synopsys translate_on

// Location: FF_X58_Y36_N29
dffeas \plif_idex.extimm_l[3] (
	.clk(CPUCLK),
	.d(\extimm_l~33_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\plif_idex.aluop_l[1]~8_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(plif_idexextimm_l_3),
	.prn(vcc));
// synopsys translate_off
defparam \plif_idex.extimm_l[3] .is_wysiwyg = "true";
defparam \plif_idex.extimm_l[3] .power_up = "low";
// synopsys translate_on

// Location: FF_X58_Y36_N3
dffeas \plif_idex.rdat2_l[3] (
	.clk(CPUCLK),
	.d(\rdat2_l~30_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\plif_idex.aluop_l[1]~8_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(plif_idexrdat2_l_3),
	.prn(vcc));
// synopsys translate_off
defparam \plif_idex.rdat2_l[3] .is_wysiwyg = "true";
defparam \plif_idex.rdat2_l[3] .power_up = "low";
// synopsys translate_on

// Location: FF_X63_Y36_N1
dffeas \plif_idex.rdat1_l[16] (
	.clk(CPUCLK),
	.d(\rdat1_l~8_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\plif_idex.aluop_l[1]~8_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(plif_idexrdat1_l_16),
	.prn(vcc));
// synopsys translate_off
defparam \plif_idex.rdat1_l[16] .is_wysiwyg = "true";
defparam \plif_idex.rdat1_l[16] .power_up = "low";
// synopsys translate_on

// Location: FF_X58_Y40_N23
dffeas \plif_idex.rdat1_l[15] (
	.clk(CPUCLK),
	.d(\rdat1_l~9_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\plif_idex.aluop_l[1]~8_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(plif_idexrdat1_l_15),
	.prn(vcc));
// synopsys translate_off
defparam \plif_idex.rdat1_l[15] .is_wysiwyg = "true";
defparam \plif_idex.rdat1_l[15] .power_up = "low";
// synopsys translate_on

// Location: FF_X66_Y30_N15
dffeas \plif_idex.rdat1_l[14] (
	.clk(CPUCLK),
	.d(\rdat1_l~10_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\plif_idex.aluop_l[1]~8_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(plif_idexrdat1_l_14),
	.prn(vcc));
// synopsys translate_off
defparam \plif_idex.rdat1_l[14] .is_wysiwyg = "true";
defparam \plif_idex.rdat1_l[14] .power_up = "low";
// synopsys translate_on

// Location: FF_X63_Y38_N5
dffeas \plif_idex.rdat1_l[13] (
	.clk(CPUCLK),
	.d(\rdat1_l~11_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\plif_idex.aluop_l[1]~8_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(plif_idexrdat1_l_13),
	.prn(vcc));
// synopsys translate_off
defparam \plif_idex.rdat1_l[13] .is_wysiwyg = "true";
defparam \plif_idex.rdat1_l[13] .power_up = "low";
// synopsys translate_on

// Location: FF_X61_Y30_N3
dffeas \plif_idex.rdat1_l[12] (
	.clk(CPUCLK),
	.d(\rdat1_l~12_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\plif_idex.aluop_l[1]~8_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(plif_idexrdat1_l_12),
	.prn(vcc));
// synopsys translate_off
defparam \plif_idex.rdat1_l[12] .is_wysiwyg = "true";
defparam \plif_idex.rdat1_l[12] .power_up = "low";
// synopsys translate_on

// Location: FF_X63_Y38_N19
dffeas \plif_idex.rdat1_l[11] (
	.clk(CPUCLK),
	.d(\rdat1_l~13_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\plif_idex.aluop_l[1]~8_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(plif_idexrdat1_l_11),
	.prn(vcc));
// synopsys translate_off
defparam \plif_idex.rdat1_l[11] .is_wysiwyg = "true";
defparam \plif_idex.rdat1_l[11] .power_up = "low";
// synopsys translate_on

// Location: FF_X70_Y36_N5
dffeas \plif_idex.rdat1_l[10] (
	.clk(CPUCLK),
	.d(\rdat1_l~14_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\plif_idex.aluop_l[1]~8_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(plif_idexrdat1_l_10),
	.prn(vcc));
// synopsys translate_off
defparam \plif_idex.rdat1_l[10] .is_wysiwyg = "true";
defparam \plif_idex.rdat1_l[10] .power_up = "low";
// synopsys translate_on

// Location: FF_X57_Y41_N13
dffeas \plif_idex.rdat1_l[9] (
	.clk(CPUCLK),
	.d(\rdat1_l~15_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\plif_idex.aluop_l[1]~8_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(plif_idexrdat1_l_9),
	.prn(vcc));
// synopsys translate_off
defparam \plif_idex.rdat1_l[9] .is_wysiwyg = "true";
defparam \plif_idex.rdat1_l[9] .power_up = "low";
// synopsys translate_on

// Location: FF_X58_Y41_N15
dffeas \plif_idex.rdat2_l[4] (
	.clk(CPUCLK),
	.d(\rdat2_l~31_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\plif_idex.aluop_l[1]~8_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(plif_idexrdat2_l_4),
	.prn(vcc));
// synopsys translate_off
defparam \plif_idex.rdat2_l[4] .is_wysiwyg = "true";
defparam \plif_idex.rdat2_l[4] .power_up = "low";
// synopsys translate_on

// Location: FF_X58_Y41_N21
dffeas \plif_idex.extimm_l[4] (
	.clk(CPUCLK),
	.d(\plif_idex.extimm_l[4]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\plif_idex.aluop_l[1]~8_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(plif_idexextimm_l_4),
	.prn(vcc));
// synopsys translate_off
defparam \plif_idex.extimm_l[4] .is_wysiwyg = "true";
defparam \plif_idex.extimm_l[4] .power_up = "low";
// synopsys translate_on

// Location: FF_X61_Y33_N25
dffeas \plif_idex.rdat1_l[31] (
	.clk(CPUCLK),
	.d(\rdat1_l~16_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\plif_idex.aluop_l[1]~8_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(plif_idexrdat1_l_31),
	.prn(vcc));
// synopsys translate_off
defparam \plif_idex.rdat1_l[31] .is_wysiwyg = "true";
defparam \plif_idex.rdat1_l[31] .power_up = "low";
// synopsys translate_on

// Location: FF_X61_Y33_N3
dffeas \plif_idex.rdat1_l[29] (
	.clk(CPUCLK),
	.d(\rdat1_l~17_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\plif_idex.aluop_l[1]~8_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(plif_idexrdat1_l_29),
	.prn(vcc));
// synopsys translate_off
defparam \plif_idex.rdat1_l[29] .is_wysiwyg = "true";
defparam \plif_idex.rdat1_l[29] .power_up = "low";
// synopsys translate_on

// Location: FF_X61_Y33_N9
dffeas \plif_idex.rdat1_l[30] (
	.clk(CPUCLK),
	.d(\rdat1_l~18_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\plif_idex.aluop_l[1]~8_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(plif_idexrdat1_l_30),
	.prn(vcc));
// synopsys translate_off
defparam \plif_idex.rdat1_l[30] .is_wysiwyg = "true";
defparam \plif_idex.rdat1_l[30] .power_up = "low";
// synopsys translate_on

// Location: FF_X63_Y39_N27
dffeas \plif_idex.rdat1_l[28] (
	.clk(CPUCLK),
	.d(\rdat1_l~19_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\plif_idex.aluop_l[1]~8_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(plif_idexrdat1_l_28),
	.prn(vcc));
// synopsys translate_off
defparam \plif_idex.rdat1_l[28] .is_wysiwyg = "true";
defparam \plif_idex.rdat1_l[28] .power_up = "low";
// synopsys translate_on

// Location: FF_X63_Y39_N5
dffeas \plif_idex.rdat1_l[27] (
	.clk(CPUCLK),
	.d(\rdat1_l~20_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\plif_idex.aluop_l[1]~8_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(plif_idexrdat1_l_27),
	.prn(vcc));
// synopsys translate_off
defparam \plif_idex.rdat1_l[27] .is_wysiwyg = "true";
defparam \plif_idex.rdat1_l[27] .power_up = "low";
// synopsys translate_on

// Location: FF_X63_Y32_N7
dffeas \plif_idex.rdat1_l[26] (
	.clk(CPUCLK),
	.d(\rdat1_l~21_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\plif_idex.aluop_l[1]~8_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(plif_idexrdat1_l_26),
	.prn(vcc));
// synopsys translate_off
defparam \plif_idex.rdat1_l[26] .is_wysiwyg = "true";
defparam \plif_idex.rdat1_l[26] .power_up = "low";
// synopsys translate_on

// Location: FF_X65_Y31_N15
dffeas \plif_idex.rdat1_l[25] (
	.clk(CPUCLK),
	.d(\rdat1_l~22_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\plif_idex.aluop_l[1]~8_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(plif_idexrdat1_l_25),
	.prn(vcc));
// synopsys translate_off
defparam \plif_idex.rdat1_l[25] .is_wysiwyg = "true";
defparam \plif_idex.rdat1_l[25] .power_up = "low";
// synopsys translate_on

// Location: FF_X59_Y34_N23
dffeas \plif_idex.rdat1_l[24] (
	.clk(CPUCLK),
	.d(\rdat1_l~23_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\plif_idex.aluop_l[1]~8_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(plif_idexrdat1_l_24),
	.prn(vcc));
// synopsys translate_off
defparam \plif_idex.rdat1_l[24] .is_wysiwyg = "true";
defparam \plif_idex.rdat1_l[24] .power_up = "low";
// synopsys translate_on

// Location: FF_X70_Y37_N11
dffeas \plif_idex.rdat1_l[23] (
	.clk(CPUCLK),
	.d(\rdat1_l~24_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\plif_idex.aluop_l[1]~8_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(plif_idexrdat1_l_23),
	.prn(vcc));
// synopsys translate_off
defparam \plif_idex.rdat1_l[23] .is_wysiwyg = "true";
defparam \plif_idex.rdat1_l[23] .power_up = "low";
// synopsys translate_on

// Location: FF_X68_Y36_N15
dffeas \plif_idex.rdat1_l[22] (
	.clk(CPUCLK),
	.d(\rdat1_l~25_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\plif_idex.aluop_l[1]~8_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(plif_idexrdat1_l_22),
	.prn(vcc));
// synopsys translate_off
defparam \plif_idex.rdat1_l[22] .is_wysiwyg = "true";
defparam \plif_idex.rdat1_l[22] .power_up = "low";
// synopsys translate_on

// Location: FF_X59_Y38_N19
dffeas \plif_idex.rdat1_l[21] (
	.clk(CPUCLK),
	.d(\rdat1_l~26_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\plif_idex.aluop_l[1]~8_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(plif_idexrdat1_l_21),
	.prn(vcc));
// synopsys translate_off
defparam \plif_idex.rdat1_l[21] .is_wysiwyg = "true";
defparam \plif_idex.rdat1_l[21] .power_up = "low";
// synopsys translate_on

// Location: FF_X60_Y40_N31
dffeas \plif_idex.rdat1_l[20] (
	.clk(CPUCLK),
	.d(\rdat1_l~27_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\plif_idex.aluop_l[1]~8_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(plif_idexrdat1_l_20),
	.prn(vcc));
// synopsys translate_off
defparam \plif_idex.rdat1_l[20] .is_wysiwyg = "true";
defparam \plif_idex.rdat1_l[20] .power_up = "low";
// synopsys translate_on

// Location: FF_X67_Y36_N13
dffeas \plif_idex.rdat1_l[19] (
	.clk(CPUCLK),
	.d(\rdat1_l~28_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\plif_idex.aluop_l[1]~8_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(plif_idexrdat1_l_19),
	.prn(vcc));
// synopsys translate_off
defparam \plif_idex.rdat1_l[19] .is_wysiwyg = "true";
defparam \plif_idex.rdat1_l[19] .power_up = "low";
// synopsys translate_on

// Location: FF_X63_Y36_N11
dffeas \plif_idex.rdat1_l[18] (
	.clk(CPUCLK),
	.d(\rdat1_l~29_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\plif_idex.aluop_l[1]~8_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(plif_idexrdat1_l_18),
	.prn(vcc));
// synopsys translate_off
defparam \plif_idex.rdat1_l[18] .is_wysiwyg = "true";
defparam \plif_idex.rdat1_l[18] .power_up = "low";
// synopsys translate_on

// Location: FF_X56_Y40_N17
dffeas \plif_idex.rdat1_l[17] (
	.clk(CPUCLK),
	.d(\rdat1_l~30_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\plif_idex.aluop_l[1]~8_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(plif_idexrdat1_l_17),
	.prn(vcc));
// synopsys translate_off
defparam \plif_idex.rdat1_l[17] .is_wysiwyg = "true";
defparam \plif_idex.rdat1_l[17] .power_up = "low";
// synopsys translate_on

// Location: FF_X55_Y40_N17
dffeas \plif_idex.rdat1_l[0] (
	.clk(CPUCLK),
	.d(\rdat1_l~31_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\plif_idex.aluop_l[1]~8_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(plif_idexrdat1_l_0),
	.prn(vcc));
// synopsys translate_off
defparam \plif_idex.rdat1_l[0] .is_wysiwyg = "true";
defparam \plif_idex.rdat1_l[0] .power_up = "low";
// synopsys translate_on

// Location: FF_X58_Y33_N23
dffeas \plif_idex.dmemREN_l (
	.clk(CPUCLK),
	.d(\dmemREN_l~0_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\plif_idex.aluop_l[1]~8_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(plif_idexdmemREN_l),
	.prn(vcc));
// synopsys translate_off
defparam \plif_idex.dmemREN_l .is_wysiwyg = "true";
defparam \plif_idex.dmemREN_l .power_up = "low";
// synopsys translate_on

// Location: FF_X60_Y32_N9
dffeas \plif_idex.wsel_l[0] (
	.clk(CPUCLK),
	.d(\wsel_l~2_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\plif_idex.aluop_l[1]~8_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(plif_idexwsel_l_0),
	.prn(vcc));
// synopsys translate_off
defparam \plif_idex.wsel_l[0] .is_wysiwyg = "true";
defparam \plif_idex.wsel_l[0] .power_up = "low";
// synopsys translate_on

// Location: FF_X60_Y32_N23
dffeas \plif_idex.wsel_l[1] (
	.clk(CPUCLK),
	.d(\wsel_l~4_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\plif_idex.aluop_l[1]~8_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(plif_idexwsel_l_1),
	.prn(vcc));
// synopsys translate_off
defparam \plif_idex.wsel_l[1] .is_wysiwyg = "true";
defparam \plif_idex.wsel_l[1] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X59_Y30_N4
cycloneive_lcell_comb \aluop_l~0 (
// Equation(s):
// aluop_l = (((plif_ifidinstr_l_26 & plif_ifidinstr_l_27)) # (!plif_ifidinstr_l_28)) # (!Equal13)

	.dataa(plif_ifidinstr_l_26),
	.datab(Equal13),
	.datac(plif_ifidinstr_l_28),
	.datad(plif_ifidinstr_l_27),
	.cin(gnd),
	.combout(aluop_l),
	.cout());
// synopsys translate_off
defparam \aluop_l~0 .lut_mask = 16'hBF3F;
defparam \aluop_l~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X60_Y32_N27
dffeas \plif_idex.wsel_l[2] (
	.clk(CPUCLK),
	.d(\wsel_l~6_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\plif_idex.aluop_l[1]~8_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(plif_idexwsel_l_2),
	.prn(vcc));
// synopsys translate_off
defparam \plif_idex.wsel_l[2] .is_wysiwyg = "true";
defparam \plif_idex.wsel_l[2] .power_up = "low";
// synopsys translate_on

// Location: FF_X60_Y32_N25
dffeas \plif_idex.wsel_l[3] (
	.clk(CPUCLK),
	.d(\wsel_l~8_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\plif_idex.aluop_l[1]~8_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(plif_idexwsel_l_3),
	.prn(vcc));
// synopsys translate_off
defparam \plif_idex.wsel_l[3] .is_wysiwyg = "true";
defparam \plif_idex.wsel_l[3] .power_up = "low";
// synopsys translate_on

// Location: FF_X60_Y32_N5
dffeas \plif_idex.wsel_l[4] (
	.clk(CPUCLK),
	.d(\wsel_l~10_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\plif_idex.aluop_l[1]~8_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(plif_idexwsel_l_4),
	.prn(vcc));
// synopsys translate_off
defparam \plif_idex.wsel_l[4] .is_wysiwyg = "true";
defparam \plif_idex.wsel_l[4] .power_up = "low";
// synopsys translate_on

// Location: FF_X56_Y30_N27
dffeas \plif_idex.dmemWEN_l (
	.clk(CPUCLK),
	.d(\dmemWEN_l~0_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\plif_idex.aluop_l[1]~8_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(plif_idexdmemWEN_l),
	.prn(vcc));
// synopsys translate_off
defparam \plif_idex.dmemWEN_l .is_wysiwyg = "true";
defparam \plif_idex.dmemWEN_l .power_up = "low";
// synopsys translate_on

// Location: FF_X60_Y32_N1
dffeas \plif_idex.regen_l (
	.clk(CPUCLK),
	.d(\regen_l~0_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\plif_idex.aluop_l[1]~8_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(plif_idexregen_l),
	.prn(vcc));
// synopsys translate_off
defparam \plif_idex.regen_l .is_wysiwyg = "true";
defparam \plif_idex.regen_l .power_up = "low";
// synopsys translate_on

// Location: FF_X57_Y32_N21
dffeas \plif_idex.regsrc_l[0] (
	.clk(CPUCLK),
	.d(\regsrc_l~0_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\plif_idex.aluop_l[1]~8_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(plif_idexregsrc_l_0),
	.prn(vcc));
// synopsys translate_off
defparam \plif_idex.regsrc_l[0] .is_wysiwyg = "true";
defparam \plif_idex.regsrc_l[0] .power_up = "low";
// synopsys translate_on

// Location: FF_X58_Y33_N21
dffeas \plif_idex.regsrc_l[1] (
	.clk(CPUCLK),
	.d(\regsrc_l~1_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\plif_idex.aluop_l[1]~8_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(plif_idexregsrc_l_1),
	.prn(vcc));
// synopsys translate_off
defparam \plif_idex.regsrc_l[1] .is_wysiwyg = "true";
defparam \plif_idex.regsrc_l[1] .power_up = "low";
// synopsys translate_on

// Location: FF_X58_Y31_N27
dffeas \plif_idex.rtnaddr_l[31] (
	.clk(CPUCLK),
	.d(\rtnaddr_l~0_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\plif_idex.aluop_l[1]~8_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(plif_idexrtnaddr_l_31),
	.prn(vcc));
// synopsys translate_off
defparam \plif_idex.rtnaddr_l[31] .is_wysiwyg = "true";
defparam \plif_idex.rtnaddr_l[31] .power_up = "low";
// synopsys translate_on

// Location: FF_X58_Y31_N17
dffeas \plif_idex.rtnaddr_l[30] (
	.clk(CPUCLK),
	.d(\rtnaddr_l~1_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\plif_idex.aluop_l[1]~8_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(plif_idexrtnaddr_l_30),
	.prn(vcc));
// synopsys translate_off
defparam \plif_idex.rtnaddr_l[30] .is_wysiwyg = "true";
defparam \plif_idex.rtnaddr_l[30] .power_up = "low";
// synopsys translate_on

// Location: FF_X58_Y31_N15
dffeas \plif_idex.rtnaddr_l[29] (
	.clk(CPUCLK),
	.d(\rtnaddr_l~2_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\plif_idex.aluop_l[1]~8_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(plif_idexrtnaddr_l_29),
	.prn(vcc));
// synopsys translate_off
defparam \plif_idex.rtnaddr_l[29] .is_wysiwyg = "true";
defparam \plif_idex.rtnaddr_l[29] .power_up = "low";
// synopsys translate_on

// Location: FF_X54_Y31_N11
dffeas \plif_idex.rtnaddr_l[28] (
	.clk(CPUCLK),
	.d(\rtnaddr_l~3_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\plif_idex.aluop_l[1]~8_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(plif_idexrtnaddr_l_28),
	.prn(vcc));
// synopsys translate_off
defparam \plif_idex.rtnaddr_l[28] .is_wysiwyg = "true";
defparam \plif_idex.rtnaddr_l[28] .power_up = "low";
// synopsys translate_on

// Location: FF_X52_Y31_N13
dffeas \plif_idex.rtnaddr_l[27] (
	.clk(CPUCLK),
	.d(\rtnaddr_l~4_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\plif_idex.aluop_l[1]~8_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(plif_idexrtnaddr_l_27),
	.prn(vcc));
// synopsys translate_off
defparam \plif_idex.rtnaddr_l[27] .is_wysiwyg = "true";
defparam \plif_idex.rtnaddr_l[27] .power_up = "low";
// synopsys translate_on

// Location: FF_X52_Y31_N11
dffeas \plif_idex.rtnaddr_l[26] (
	.clk(CPUCLK),
	.d(\rtnaddr_l~5_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\plif_idex.aluop_l[1]~8_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(plif_idexrtnaddr_l_26),
	.prn(vcc));
// synopsys translate_off
defparam \plif_idex.rtnaddr_l[26] .is_wysiwyg = "true";
defparam \plif_idex.rtnaddr_l[26] .power_up = "low";
// synopsys translate_on

// Location: FF_X52_Y31_N21
dffeas \plif_idex.rtnaddr_l[25] (
	.clk(CPUCLK),
	.d(\rtnaddr_l~6_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\plif_idex.aluop_l[1]~8_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(plif_idexrtnaddr_l_25),
	.prn(vcc));
// synopsys translate_off
defparam \plif_idex.rtnaddr_l[25] .is_wysiwyg = "true";
defparam \plif_idex.rtnaddr_l[25] .power_up = "low";
// synopsys translate_on

// Location: FF_X52_Y31_N3
dffeas \plif_idex.rtnaddr_l[24] (
	.clk(CPUCLK),
	.d(\rtnaddr_l~7_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\plif_idex.aluop_l[1]~8_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(plif_idexrtnaddr_l_24),
	.prn(vcc));
// synopsys translate_off
defparam \plif_idex.rtnaddr_l[24] .is_wysiwyg = "true";
defparam \plif_idex.rtnaddr_l[24] .power_up = "low";
// synopsys translate_on

// Location: FF_X52_Y31_N25
dffeas \plif_idex.rtnaddr_l[23] (
	.clk(CPUCLK),
	.d(\rtnaddr_l~8_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\plif_idex.aluop_l[1]~8_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(plif_idexrtnaddr_l_23),
	.prn(vcc));
// synopsys translate_off
defparam \plif_idex.rtnaddr_l[23] .is_wysiwyg = "true";
defparam \plif_idex.rtnaddr_l[23] .power_up = "low";
// synopsys translate_on

// Location: FF_X52_Y31_N7
dffeas \plif_idex.rtnaddr_l[22] (
	.clk(CPUCLK),
	.d(\rtnaddr_l~9_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\plif_idex.aluop_l[1]~8_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(plif_idexrtnaddr_l_22),
	.prn(vcc));
// synopsys translate_off
defparam \plif_idex.rtnaddr_l[22] .is_wysiwyg = "true";
defparam \plif_idex.rtnaddr_l[22] .power_up = "low";
// synopsys translate_on

// Location: FF_X53_Y30_N1
dffeas \plif_idex.rtnaddr_l[21] (
	.clk(CPUCLK),
	.d(\rtnaddr_l~10_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\plif_idex.aluop_l[1]~8_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(plif_idexrtnaddr_l_21),
	.prn(vcc));
// synopsys translate_off
defparam \plif_idex.rtnaddr_l[21] .is_wysiwyg = "true";
defparam \plif_idex.rtnaddr_l[21] .power_up = "low";
// synopsys translate_on

// Location: FF_X53_Y30_N3
dffeas \plif_idex.rtnaddr_l[20] (
	.clk(CPUCLK),
	.d(\rtnaddr_l~11_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\plif_idex.aluop_l[1]~8_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(plif_idexrtnaddr_l_20),
	.prn(vcc));
// synopsys translate_off
defparam \plif_idex.rtnaddr_l[20] .is_wysiwyg = "true";
defparam \plif_idex.rtnaddr_l[20] .power_up = "low";
// synopsys translate_on

// Location: FF_X53_Y30_N25
dffeas \plif_idex.rtnaddr_l[19] (
	.clk(CPUCLK),
	.d(\rtnaddr_l~12_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\plif_idex.aluop_l[1]~8_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(plif_idexrtnaddr_l_19),
	.prn(vcc));
// synopsys translate_off
defparam \plif_idex.rtnaddr_l[19] .is_wysiwyg = "true";
defparam \plif_idex.rtnaddr_l[19] .power_up = "low";
// synopsys translate_on

// Location: FF_X53_Y30_N27
dffeas \plif_idex.rtnaddr_l[18] (
	.clk(CPUCLK),
	.d(\rtnaddr_l~13_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\plif_idex.aluop_l[1]~8_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(plif_idexrtnaddr_l_18),
	.prn(vcc));
// synopsys translate_off
defparam \plif_idex.rtnaddr_l[18] .is_wysiwyg = "true";
defparam \plif_idex.rtnaddr_l[18] .power_up = "low";
// synopsys translate_on

// Location: FF_X53_Y30_N17
dffeas \plif_idex.rtnaddr_l[17] (
	.clk(CPUCLK),
	.d(\rtnaddr_l~14_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\plif_idex.aluop_l[1]~8_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(plif_idexrtnaddr_l_17),
	.prn(vcc));
// synopsys translate_off
defparam \plif_idex.rtnaddr_l[17] .is_wysiwyg = "true";
defparam \plif_idex.rtnaddr_l[17] .power_up = "low";
// synopsys translate_on

// Location: FF_X53_Y30_N23
dffeas \plif_idex.rtnaddr_l[16] (
	.clk(CPUCLK),
	.d(\rtnaddr_l~15_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\plif_idex.aluop_l[1]~8_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(plif_idexrtnaddr_l_16),
	.prn(vcc));
// synopsys translate_off
defparam \plif_idex.rtnaddr_l[16] .is_wysiwyg = "true";
defparam \plif_idex.rtnaddr_l[16] .power_up = "low";
// synopsys translate_on

// Location: FF_X53_Y30_N21
dffeas \plif_idex.rtnaddr_l[15] (
	.clk(CPUCLK),
	.d(\rtnaddr_l~16_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\plif_idex.aluop_l[1]~8_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(plif_idexrtnaddr_l_15),
	.prn(vcc));
// synopsys translate_off
defparam \plif_idex.rtnaddr_l[15] .is_wysiwyg = "true";
defparam \plif_idex.rtnaddr_l[15] .power_up = "low";
// synopsys translate_on

// Location: FF_X53_Y30_N31
dffeas \plif_idex.rtnaddr_l[14] (
	.clk(CPUCLK),
	.d(\rtnaddr_l~17_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\plif_idex.aluop_l[1]~8_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(plif_idexrtnaddr_l_14),
	.prn(vcc));
// synopsys translate_off
defparam \plif_idex.rtnaddr_l[14] .is_wysiwyg = "true";
defparam \plif_idex.rtnaddr_l[14] .power_up = "low";
// synopsys translate_on

// Location: FF_X54_Y31_N21
dffeas \plif_idex.rtnaddr_l[13] (
	.clk(CPUCLK),
	.d(\rtnaddr_l~18_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\plif_idex.aluop_l[1]~8_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(plif_idexrtnaddr_l_13),
	.prn(vcc));
// synopsys translate_off
defparam \plif_idex.rtnaddr_l[13] .is_wysiwyg = "true";
defparam \plif_idex.rtnaddr_l[13] .power_up = "low";
// synopsys translate_on

// Location: FF_X54_Y31_N15
dffeas \plif_idex.rtnaddr_l[12] (
	.clk(CPUCLK),
	.d(\rtnaddr_l~19_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\plif_idex.aluop_l[1]~8_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(plif_idexrtnaddr_l_12),
	.prn(vcc));
// synopsys translate_off
defparam \plif_idex.rtnaddr_l[12] .is_wysiwyg = "true";
defparam \plif_idex.rtnaddr_l[12] .power_up = "low";
// synopsys translate_on

// Location: FF_X54_Y31_N29
dffeas \plif_idex.rtnaddr_l[11] (
	.clk(CPUCLK),
	.d(\rtnaddr_l~20_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\plif_idex.aluop_l[1]~8_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(plif_idexrtnaddr_l_11),
	.prn(vcc));
// synopsys translate_off
defparam \plif_idex.rtnaddr_l[11] .is_wysiwyg = "true";
defparam \plif_idex.rtnaddr_l[11] .power_up = "low";
// synopsys translate_on

// Location: FF_X54_Y31_N31
dffeas \plif_idex.rtnaddr_l[10] (
	.clk(CPUCLK),
	.d(\rtnaddr_l~21_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\plif_idex.aluop_l[1]~8_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(plif_idexrtnaddr_l_10),
	.prn(vcc));
// synopsys translate_off
defparam \plif_idex.rtnaddr_l[10] .is_wysiwyg = "true";
defparam \plif_idex.rtnaddr_l[10] .power_up = "low";
// synopsys translate_on

// Location: FF_X54_Y31_N25
dffeas \plif_idex.rtnaddr_l[9] (
	.clk(CPUCLK),
	.d(\rtnaddr_l~22_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\plif_idex.aluop_l[1]~8_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(plif_idexrtnaddr_l_9),
	.prn(vcc));
// synopsys translate_off
defparam \plif_idex.rtnaddr_l[9] .is_wysiwyg = "true";
defparam \plif_idex.rtnaddr_l[9] .power_up = "low";
// synopsys translate_on

// Location: FF_X54_Y31_N3
dffeas \plif_idex.rtnaddr_l[8] (
	.clk(CPUCLK),
	.d(\rtnaddr_l~23_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\plif_idex.aluop_l[1]~8_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(plif_idexrtnaddr_l_8),
	.prn(vcc));
// synopsys translate_off
defparam \plif_idex.rtnaddr_l[8] .is_wysiwyg = "true";
defparam \plif_idex.rtnaddr_l[8] .power_up = "low";
// synopsys translate_on

// Location: FF_X54_Y31_N1
dffeas \plif_idex.rtnaddr_l[7] (
	.clk(CPUCLK),
	.d(\rtnaddr_l~24_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\plif_idex.aluop_l[1]~8_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(plif_idexrtnaddr_l_7),
	.prn(vcc));
// synopsys translate_off
defparam \plif_idex.rtnaddr_l[7] .is_wysiwyg = "true";
defparam \plif_idex.rtnaddr_l[7] .power_up = "low";
// synopsys translate_on

// Location: FF_X58_Y31_N21
dffeas \plif_idex.rtnaddr_l[6] (
	.clk(CPUCLK),
	.d(\rtnaddr_l~25_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\plif_idex.aluop_l[1]~8_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(plif_idexrtnaddr_l_6),
	.prn(vcc));
// synopsys translate_off
defparam \plif_idex.rtnaddr_l[6] .is_wysiwyg = "true";
defparam \plif_idex.rtnaddr_l[6] .power_up = "low";
// synopsys translate_on

// Location: FF_X54_Y31_N7
dffeas \plif_idex.rtnaddr_l[5] (
	.clk(CPUCLK),
	.d(\rtnaddr_l~26_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\plif_idex.aluop_l[1]~8_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(plif_idexrtnaddr_l_5),
	.prn(vcc));
// synopsys translate_off
defparam \plif_idex.rtnaddr_l[5] .is_wysiwyg = "true";
defparam \plif_idex.rtnaddr_l[5] .power_up = "low";
// synopsys translate_on

// Location: FF_X50_Y41_N1
dffeas \plif_idex.rtnaddr_l[2] (
	.clk(CPUCLK),
	.d(\rtnaddr_l~27_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\plif_idex.aluop_l[1]~8_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(plif_idexrtnaddr_l_2),
	.prn(vcc));
// synopsys translate_off
defparam \plif_idex.rtnaddr_l[2] .is_wysiwyg = "true";
defparam \plif_idex.rtnaddr_l[2] .power_up = "low";
// synopsys translate_on

// Location: FF_X52_Y31_N17
dffeas \plif_idex.rtnaddr_l[1] (
	.clk(CPUCLK),
	.d(\rtnaddr_l~28_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\plif_idex.aluop_l[1]~8_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(plif_idexrtnaddr_l_1),
	.prn(vcc));
// synopsys translate_off
defparam \plif_idex.rtnaddr_l[1] .is_wysiwyg = "true";
defparam \plif_idex.rtnaddr_l[1] .power_up = "low";
// synopsys translate_on

// Location: FF_X50_Y41_N23
dffeas \plif_idex.rtnaddr_l[0] (
	.clk(CPUCLK),
	.d(\rtnaddr_l~29_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\plif_idex.aluop_l[1]~8_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(plif_idexrtnaddr_l_0),
	.prn(vcc));
// synopsys translate_off
defparam \plif_idex.rtnaddr_l[0] .is_wysiwyg = "true";
defparam \plif_idex.rtnaddr_l[0] .power_up = "low";
// synopsys translate_on

// Location: FF_X50_Y41_N29
dffeas \plif_idex.rtnaddr_l[4] (
	.clk(CPUCLK),
	.d(\rtnaddr_l~30_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\plif_idex.aluop_l[1]~8_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(plif_idexrtnaddr_l_4),
	.prn(vcc));
// synopsys translate_off
defparam \plif_idex.rtnaddr_l[4] .is_wysiwyg = "true";
defparam \plif_idex.rtnaddr_l[4] .power_up = "low";
// synopsys translate_on

// Location: FF_X50_Y41_N11
dffeas \plif_idex.rtnaddr_l[3] (
	.clk(CPUCLK),
	.d(\rtnaddr_l~31_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\plif_idex.aluop_l[1]~8_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(plif_idexrtnaddr_l_3),
	.prn(vcc));
// synopsys translate_off
defparam \plif_idex.rtnaddr_l[3] .is_wysiwyg = "true";
defparam \plif_idex.rtnaddr_l[3] .power_up = "low";
// synopsys translate_on

// Location: FF_X56_Y30_N13
dffeas \plif_idex.btype_l (
	.clk(CPUCLK),
	.d(\btype_l~0_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\plif_idex.aluop_l[1]~8_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(plif_idexbtype_l),
	.prn(vcc));
// synopsys translate_off
defparam \plif_idex.btype_l .is_wysiwyg = "true";
defparam \plif_idex.btype_l .power_up = "low";
// synopsys translate_on

// Location: FF_X57_Y30_N31
dffeas \plif_idex.jaddr_l[1] (
	.clk(CPUCLK),
	.d(\jaddr_l~0_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\plif_idex.aluop_l[1]~8_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(plif_idexjaddr_l_1),
	.prn(vcc));
// synopsys translate_off
defparam \plif_idex.jaddr_l[1] .is_wysiwyg = "true";
defparam \plif_idex.jaddr_l[1] .power_up = "low";
// synopsys translate_on

// Location: FF_X58_Y33_N27
dffeas \plif_idex.jaddr_l[0] (
	.clk(CPUCLK),
	.d(\jaddr_l~1_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\plif_idex.aluop_l[1]~8_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(plif_idexjaddr_l_0),
	.prn(vcc));
// synopsys translate_off
defparam \plif_idex.jaddr_l[0] .is_wysiwyg = "true";
defparam \plif_idex.jaddr_l[0] .power_up = "low";
// synopsys translate_on

// Location: FF_X58_Y33_N1
dffeas \plif_idex.jaddr_l[3] (
	.clk(CPUCLK),
	.d(\jaddr_l~2_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\plif_idex.aluop_l[1]~8_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(plif_idexjaddr_l_3),
	.prn(vcc));
// synopsys translate_off
defparam \plif_idex.jaddr_l[3] .is_wysiwyg = "true";
defparam \plif_idex.jaddr_l[3] .power_up = "low";
// synopsys translate_on

// Location: FF_X58_Y33_N15
dffeas \plif_idex.jaddr_l[2] (
	.clk(CPUCLK),
	.d(\jaddr_l~3_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\plif_idex.aluop_l[1]~8_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(plif_idexjaddr_l_2),
	.prn(vcc));
// synopsys translate_off
defparam \plif_idex.jaddr_l[2] .is_wysiwyg = "true";
defparam \plif_idex.jaddr_l[2] .power_up = "low";
// synopsys translate_on

// Location: FF_X57_Y30_N13
dffeas \plif_idex.jaddr_l[5] (
	.clk(CPUCLK),
	.d(\jaddr_l~4_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\plif_idex.aluop_l[1]~8_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(plif_idexjaddr_l_5),
	.prn(vcc));
// synopsys translate_off
defparam \plif_idex.jaddr_l[5] .is_wysiwyg = "true";
defparam \plif_idex.jaddr_l[5] .power_up = "low";
// synopsys translate_on

// Location: FF_X58_Y33_N13
dffeas \plif_idex.jaddr_l[4] (
	.clk(CPUCLK),
	.d(\jaddr_l~5_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\plif_idex.aluop_l[1]~8_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(plif_idexjaddr_l_4),
	.prn(vcc));
// synopsys translate_off
defparam \plif_idex.jaddr_l[4] .is_wysiwyg = "true";
defparam \plif_idex.jaddr_l[4] .power_up = "low";
// synopsys translate_on

// Location: FF_X57_Y32_N15
dffeas \plif_idex.jaddr_l[7] (
	.clk(CPUCLK),
	.d(\jaddr_l~6_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\plif_idex.aluop_l[1]~8_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(plif_idexjaddr_l_7),
	.prn(vcc));
// synopsys translate_off
defparam \plif_idex.jaddr_l[7] .is_wysiwyg = "true";
defparam \plif_idex.jaddr_l[7] .power_up = "low";
// synopsys translate_on

// Location: FF_X58_Y33_N31
dffeas \plif_idex.jaddr_l[6] (
	.clk(CPUCLK),
	.d(\jaddr_l~7_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\plif_idex.aluop_l[1]~8_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(plif_idexjaddr_l_6),
	.prn(vcc));
// synopsys translate_off
defparam \plif_idex.jaddr_l[6] .is_wysiwyg = "true";
defparam \plif_idex.jaddr_l[6] .power_up = "low";
// synopsys translate_on

// Location: FF_X58_Y33_N25
dffeas \plif_idex.jaddr_l[9] (
	.clk(CPUCLK),
	.d(\jaddr_l~8_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\plif_idex.aluop_l[1]~8_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(plif_idexjaddr_l_9),
	.prn(vcc));
// synopsys translate_off
defparam \plif_idex.jaddr_l[9] .is_wysiwyg = "true";
defparam \plif_idex.jaddr_l[9] .power_up = "low";
// synopsys translate_on

// Location: FF_X58_Y33_N7
dffeas \plif_idex.jaddr_l[8] (
	.clk(CPUCLK),
	.d(\jaddr_l~9_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\plif_idex.aluop_l[1]~8_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(plif_idexjaddr_l_8),
	.prn(vcc));
// synopsys translate_off
defparam \plif_idex.jaddr_l[8] .is_wysiwyg = "true";
defparam \plif_idex.jaddr_l[8] .power_up = "low";
// synopsys translate_on

// Location: FF_X58_Y33_N5
dffeas \plif_idex.jaddr_l[11] (
	.clk(CPUCLK),
	.d(\jaddr_l~10_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\plif_idex.aluop_l[1]~8_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(plif_idexjaddr_l_11),
	.prn(vcc));
// synopsys translate_off
defparam \plif_idex.jaddr_l[11] .is_wysiwyg = "true";
defparam \plif_idex.jaddr_l[11] .power_up = "low";
// synopsys translate_on

// Location: FF_X58_Y33_N3
dffeas \plif_idex.jaddr_l[10] (
	.clk(CPUCLK),
	.d(\jaddr_l~11_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\plif_idex.aluop_l[1]~8_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(plif_idexjaddr_l_10),
	.prn(vcc));
// synopsys translate_off
defparam \plif_idex.jaddr_l[10] .is_wysiwyg = "true";
defparam \plif_idex.jaddr_l[10] .power_up = "low";
// synopsys translate_on

// Location: FF_X57_Y32_N29
dffeas \plif_idex.jaddr_l[13] (
	.clk(CPUCLK),
	.d(\jaddr_l~12_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\plif_idex.aluop_l[1]~8_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(plif_idexjaddr_l_13),
	.prn(vcc));
// synopsys translate_off
defparam \plif_idex.jaddr_l[13] .is_wysiwyg = "true";
defparam \plif_idex.jaddr_l[13] .power_up = "low";
// synopsys translate_on

// Location: FF_X58_Y31_N3
dffeas \plif_idex.jaddr_l[12] (
	.clk(CPUCLK),
	.d(\jaddr_l~13_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\plif_idex.aluop_l[1]~8_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(plif_idexjaddr_l_12),
	.prn(vcc));
// synopsys translate_off
defparam \plif_idex.jaddr_l[12] .is_wysiwyg = "true";
defparam \plif_idex.jaddr_l[12] .power_up = "low";
// synopsys translate_on

// Location: FF_X58_Y31_N25
dffeas \plif_idex.jaddr_l[15] (
	.clk(CPUCLK),
	.d(\jaddr_l~14_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\plif_idex.aluop_l[1]~8_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(plif_idexjaddr_l_15),
	.prn(vcc));
// synopsys translate_off
defparam \plif_idex.jaddr_l[15] .is_wysiwyg = "true";
defparam \plif_idex.jaddr_l[15] .power_up = "low";
// synopsys translate_on

// Location: FF_X57_Y30_N27
dffeas \plif_idex.jaddr_l[14] (
	.clk(CPUCLK),
	.d(\jaddr_l~15_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\plif_idex.aluop_l[1]~8_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(plif_idexjaddr_l_14),
	.prn(vcc));
// synopsys translate_off
defparam \plif_idex.jaddr_l[14] .is_wysiwyg = "true";
defparam \plif_idex.jaddr_l[14] .power_up = "low";
// synopsys translate_on

// Location: FF_X58_Y31_N19
dffeas \plif_idex.jaddr_l[17] (
	.clk(CPUCLK),
	.d(\jaddr_l~16_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\plif_idex.aluop_l[1]~8_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(plif_idexjaddr_l_17),
	.prn(vcc));
// synopsys translate_off
defparam \plif_idex.jaddr_l[17] .is_wysiwyg = "true";
defparam \plif_idex.jaddr_l[17] .power_up = "low";
// synopsys translate_on

// Location: FF_X58_Y33_N17
dffeas \plif_idex.jaddr_l[16] (
	.clk(CPUCLK),
	.d(\jaddr_l~17_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\plif_idex.aluop_l[1]~8_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(plif_idexjaddr_l_16),
	.prn(vcc));
// synopsys translate_off
defparam \plif_idex.jaddr_l[16] .is_wysiwyg = "true";
defparam \plif_idex.jaddr_l[16] .power_up = "low";
// synopsys translate_on

// Location: FF_X59_Y37_N11
dffeas \plif_idex.jaddr_l[19] (
	.clk(CPUCLK),
	.d(\jaddr_l~18_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\plif_idex.aluop_l[1]~8_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(plif_idexjaddr_l_19),
	.prn(vcc));
// synopsys translate_off
defparam \plif_idex.jaddr_l[19] .is_wysiwyg = "true";
defparam \plif_idex.jaddr_l[19] .power_up = "low";
// synopsys translate_on

// Location: FF_X59_Y37_N9
dffeas \plif_idex.jaddr_l[18] (
	.clk(CPUCLK),
	.d(\jaddr_l~19_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\plif_idex.aluop_l[1]~8_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(plif_idexjaddr_l_18),
	.prn(vcc));
// synopsys translate_off
defparam \plif_idex.jaddr_l[18] .is_wysiwyg = "true";
defparam \plif_idex.jaddr_l[18] .power_up = "low";
// synopsys translate_on

// Location: FF_X58_Y37_N15
dffeas \plif_idex.jaddr_l[21] (
	.clk(CPUCLK),
	.d(\jaddr_l~20_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\plif_idex.aluop_l[1]~8_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(plif_idexjaddr_l_21),
	.prn(vcc));
// synopsys translate_off
defparam \plif_idex.jaddr_l[21] .is_wysiwyg = "true";
defparam \plif_idex.jaddr_l[21] .power_up = "low";
// synopsys translate_on

// Location: FF_X59_Y37_N19
dffeas \plif_idex.jaddr_l[20] (
	.clk(CPUCLK),
	.d(\jaddr_l~21_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\plif_idex.aluop_l[1]~8_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(plif_idexjaddr_l_20),
	.prn(vcc));
// synopsys translate_off
defparam \plif_idex.jaddr_l[20] .is_wysiwyg = "true";
defparam \plif_idex.jaddr_l[20] .power_up = "low";
// synopsys translate_on

// Location: FF_X59_Y37_N25
dffeas \plif_idex.jaddr_l[23] (
	.clk(CPUCLK),
	.d(\jaddr_l~22_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\plif_idex.aluop_l[1]~8_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(plif_idexjaddr_l_23),
	.prn(vcc));
// synopsys translate_off
defparam \plif_idex.jaddr_l[23] .is_wysiwyg = "true";
defparam \plif_idex.jaddr_l[23] .power_up = "low";
// synopsys translate_on

// Location: FF_X58_Y33_N11
dffeas \plif_idex.jaddr_l[22] (
	.clk(CPUCLK),
	.d(\jaddr_l~23_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\plif_idex.aluop_l[1]~8_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(plif_idexjaddr_l_22),
	.prn(vcc));
// synopsys translate_off
defparam \plif_idex.jaddr_l[22] .is_wysiwyg = "true";
defparam \plif_idex.jaddr_l[22] .power_up = "low";
// synopsys translate_on

// Location: FF_X59_Y37_N15
dffeas \plif_idex.jaddr_l[25] (
	.clk(CPUCLK),
	.d(\jaddr_l~24_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\plif_idex.aluop_l[1]~8_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(plif_idexjaddr_l_25),
	.prn(vcc));
// synopsys translate_off
defparam \plif_idex.jaddr_l[25] .is_wysiwyg = "true";
defparam \plif_idex.jaddr_l[25] .power_up = "low";
// synopsys translate_on

// Location: FF_X59_Y37_N29
dffeas \plif_idex.jaddr_l[24] (
	.clk(CPUCLK),
	.d(\jaddr_l~25_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\plif_idex.aluop_l[1]~8_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(plif_idexjaddr_l_24),
	.prn(vcc));
// synopsys translate_off
defparam \plif_idex.jaddr_l[24] .is_wysiwyg = "true";
defparam \plif_idex.jaddr_l[24] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X59_Y30_N24
cycloneive_lcell_comb \hlt_l~0 (
// Equation(s):
// \hlt_l~0_combout  = (Equal23 & (!idex_sRST1 & (plif_ifidinstr_l_30 & plif_ifidinstr_l_29)))

	.dataa(Equal23),
	.datab(idex_sRST1),
	.datac(plif_ifidinstr_l_30),
	.datad(plif_ifidinstr_l_29),
	.cin(gnd),
	.combout(\hlt_l~0_combout ),
	.cout());
// synopsys translate_off
defparam \hlt_l~0 .lut_mask = 16'h2000;
defparam \hlt_l~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y32_N10
cycloneive_lcell_comb \plif_idex.aluop_l[1]~9 (
// Equation(s):
// \plif_idex.aluop_l[1]~9_combout  = (plif_memwbpcsrc_l_0) # ((plif_memwbpcsrc_l_1) # ((!plif_exmemdmemREN_l & !plif_exmemdmemWEN_l)))

	.dataa(plif_memwbpcsrc_l_0),
	.datab(plif_memwbpcsrc_l_1),
	.datac(plif_exmemdmemREN_l),
	.datad(plif_exmemdmemWEN_l),
	.cin(gnd),
	.combout(\plif_idex.aluop_l[1]~9_combout ),
	.cout());
// synopsys translate_off
defparam \plif_idex.aluop_l[1]~9 .lut_mask = 16'hEEEF;
defparam \plif_idex.aluop_l[1]~9 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y32_N4
cycloneive_lcell_comb \plif_idex.aluop_l[1]~8 (
// Equation(s):
// \plif_idex.aluop_l[1]~8_combout  = (\plif_idex.aluop_l[1]~9_combout ) # ((idex_sRST2) # ((always1) # (!ifid_sRST)))

	.dataa(\plif_idex.aluop_l[1]~9_combout ),
	.datab(idex_sRST2),
	.datac(always1),
	.datad(ifid_sRST),
	.cin(gnd),
	.combout(\plif_idex.aluop_l[1]~8_combout ),
	.cout());
// synopsys translate_off
defparam \plif_idex.aluop_l[1]~8 .lut_mask = 16'hFEFF;
defparam \plif_idex.aluop_l[1]~8 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y30_N24
cycloneive_lcell_comb \pcsrc_l~0 (
// Equation(s):
// \pcsrc_l~0_combout  = (Equal26 & (Equal6 & (plif_ifidinstr_l_3 & !plif_ifidinstr_l_1)))

	.dataa(Equal26),
	.datab(Equal6),
	.datac(plif_ifidinstr_l_3),
	.datad(plif_ifidinstr_l_1),
	.cin(gnd),
	.combout(\pcsrc_l~0_combout ),
	.cout());
// synopsys translate_off
defparam \pcsrc_l~0 .lut_mask = 16'h0080;
defparam \pcsrc_l~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y30_N4
cycloneive_lcell_comb \pcsrc_l~1 (
// Equation(s):
// \pcsrc_l~1_combout  = (!idex_sRST & (!idex_sRST2 & ((\pcsrc_l~0_combout ) # (!pcsrc))))

	.dataa(idex_sRST),
	.datab(pcsrc),
	.datac(\pcsrc_l~0_combout ),
	.datad(idex_sRST2),
	.cin(gnd),
	.combout(\pcsrc_l~1_combout ),
	.cout());
// synopsys translate_off
defparam \pcsrc_l~1 .lut_mask = 16'h0051;
defparam \pcsrc_l~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y30_N18
cycloneive_lcell_comb \pcsrc_l~2 (
// Equation(s):
// \pcsrc_l~2_combout  = (!idex_sRST & (!idex_sRST2 & ((\pcsrc_l~0_combout ) # (!Selector22))))

	.dataa(idex_sRST),
	.datab(Selector22),
	.datac(\pcsrc_l~0_combout ),
	.datad(idex_sRST2),
	.cin(gnd),
	.combout(\pcsrc_l~2_combout ),
	.cout());
// synopsys translate_off
defparam \pcsrc_l~2 .lut_mask = 16'h0051;
defparam \pcsrc_l~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y30_N14
cycloneive_lcell_comb \aluop_l~2 (
// Equation(s):
// \aluop_l~2_combout  = (!plif_ifidinstr_l_4 & (!plif_ifidinstr_l_2 & (plif_ifidinstr_l_5 & WideNor0)))

	.dataa(plif_ifidinstr_l_4),
	.datab(plif_ifidinstr_l_2),
	.datac(plif_ifidinstr_l_5),
	.datad(WideNor0),
	.cin(gnd),
	.combout(\aluop_l~2_combout ),
	.cout());
// synopsys translate_off
defparam \aluop_l~2 .lut_mask = 16'h1000;
defparam \aluop_l~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y30_N8
cycloneive_lcell_comb \aluop_l~1 (
// Equation(s):
// \aluop_l~1_combout  = (!plif_ifidinstr_l_28 & (Equal13 & plif_ifidinstr_l_27))

	.dataa(plif_ifidinstr_l_28),
	.datab(Equal13),
	.datac(gnd),
	.datad(plif_ifidinstr_l_27),
	.cin(gnd),
	.combout(\aluop_l~1_combout ),
	.cout());
// synopsys translate_off
defparam \aluop_l~1 .lut_mask = 16'h4400;
defparam \aluop_l~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y30_N28
cycloneive_lcell_comb \aluop_l~3 (
// Equation(s):
// \aluop_l~3_combout  = (!idex_sRST1 & ((\aluop_l~1_combout ) # ((\aluop_l~2_combout  & Equal26))))

	.dataa(\aluop_l~2_combout ),
	.datab(Equal26),
	.datac(\aluop_l~1_combout ),
	.datad(idex_sRST1),
	.cin(gnd),
	.combout(\aluop_l~3_combout ),
	.cout());
// synopsys translate_off
defparam \aluop_l~3 .lut_mask = 16'h00F8;
defparam \aluop_l~3 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y30_N10
cycloneive_lcell_comb \aluop_l~4 (
// Equation(s):
// \aluop_l~4_combout  = (!idex_sRST1 & (((Equal1 & Equal26)) # (!aluop_l)))

	.dataa(Equal1),
	.datab(Equal26),
	.datac(aluop_l),
	.datad(idex_sRST1),
	.cin(gnd),
	.combout(\aluop_l~4_combout ),
	.cout());
// synopsys translate_off
defparam \aluop_l~4 .lut_mask = 16'h008F;
defparam \aluop_l~4 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y30_N12
cycloneive_lcell_comb \aluop_l~6 (
// Equation(s):
// \aluop_l~6_combout  = (Equal26 & (!Equal12 & ((Selector21)))) # (!Equal26 & (((WideNor1))))

	.dataa(Equal12),
	.datab(WideNor1),
	.datac(Equal26),
	.datad(Selector21),
	.cin(gnd),
	.combout(\aluop_l~6_combout ),
	.cout());
// synopsys translate_off
defparam \aluop_l~6 .lut_mask = 16'h5C0C;
defparam \aluop_l~6 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y30_N10
cycloneive_lcell_comb \aluop_l~5 (
// Equation(s):
// \aluop_l~5_combout  = (WideOr141 & (!Equal19 & ((!Equal13) # (!Equal16))))

	.dataa(Equal16),
	.datab(Equal13),
	.datac(WideOr14),
	.datad(Equal19),
	.cin(gnd),
	.combout(\aluop_l~5_combout ),
	.cout());
// synopsys translate_off
defparam \aluop_l~5 .lut_mask = 16'h0070;
defparam \aluop_l~5 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y33_N16
cycloneive_lcell_comb \aluop_l~7 (
// Equation(s):
// \aluop_l~7_combout  = (!idex_sRST1 & ((\aluop_l~6_combout ) # ((!WideNor11) # (!\aluop_l~5_combout ))))

	.dataa(\aluop_l~6_combout ),
	.datab(\aluop_l~5_combout ),
	.datac(WideNor11),
	.datad(idex_sRST1),
	.cin(gnd),
	.combout(\aluop_l~7_combout ),
	.cout());
// synopsys translate_off
defparam \aluop_l~7 .lut_mask = 16'h00BF;
defparam \aluop_l~7 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y30_N0
cycloneive_lcell_comb \aluop_l~8 (
// Equation(s):
// \aluop_l~8_combout  = (!idex_sRST1 & ((Equal18) # ((Selector221) # (!Selector22))))

	.dataa(Equal18),
	.datab(Selector221),
	.datac(Selector22),
	.datad(idex_sRST1),
	.cin(gnd),
	.combout(\aluop_l~8_combout ),
	.cout());
// synopsys translate_off
defparam \aluop_l~8 .lut_mask = 16'h00EF;
defparam \aluop_l~8 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y33_N22
cycloneive_lcell_comb \extimm_l~0 (
// Equation(s):
// \extimm_l~0_combout  = (!WideOr151 & (plif_ifidinstr_l_15 & ((Equal20) # (WideOr142))))

	.dataa(Equal20),
	.datab(WideOr15),
	.datac(plif_ifidinstr_l_15),
	.datad(WideOr141),
	.cin(gnd),
	.combout(\extimm_l~0_combout ),
	.cout());
// synopsys translate_off
defparam \extimm_l~0 .lut_mask = 16'h3020;
defparam \extimm_l~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y33_N28
cycloneive_lcell_comb \extimm_l~1 (
// Equation(s):
// \extimm_l~1_combout  = (!idex_sRST & (\extimm_l~0_combout  & !idex_sRST2))

	.dataa(idex_sRST),
	.datab(gnd),
	.datac(\extimm_l~0_combout ),
	.datad(idex_sRST2),
	.cin(gnd),
	.combout(\extimm_l~1_combout ),
	.cout());
// synopsys translate_off
defparam \extimm_l~1 .lut_mask = 16'h0050;
defparam \extimm_l~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y33_N10
cycloneive_lcell_comb \alusrc_l~0 (
// Equation(s):
// \alusrc_l~0_combout  = (!idex_sRST1 & ((Selector0) # ((Equal22) # (!WideOr161))))

	.dataa(Selector0),
	.datab(Equal22),
	.datac(idex_sRST1),
	.datad(WideOr16),
	.cin(gnd),
	.combout(\alusrc_l~0_combout ),
	.cout());
// synopsys translate_off
defparam \alusrc_l~0 .lut_mask = 16'h0E0F;
defparam \alusrc_l~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y37_N16
cycloneive_lcell_comb \rsel2_l~10 (
// Equation(s):
// \rsel2_l~10_combout  = (!idex_sRST & (Selector9 & (!idex_sRST2 & plif_ifidinstr_l_17)))

	.dataa(idex_sRST),
	.datab(Selector9),
	.datac(idex_sRST2),
	.datad(plif_ifidinstr_l_17),
	.cin(gnd),
	.combout(\rsel2_l~10_combout ),
	.cout());
// synopsys translate_off
defparam \rsel2_l~10 .lut_mask = 16'h0400;
defparam \rsel2_l~10 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y37_N6
cycloneive_lcell_comb \rsel2_l~11 (
// Equation(s):
// \rsel2_l~11_combout  = (!idex_sRST & (Selector9 & (!idex_sRST2 & plif_ifidinstr_l_16)))

	.dataa(idex_sRST),
	.datab(Selector9),
	.datac(idex_sRST2),
	.datad(plif_ifidinstr_l_16),
	.cin(gnd),
	.combout(\rsel2_l~11_combout ),
	.cout());
// synopsys translate_off
defparam \rsel2_l~11 .lut_mask = 16'h0400;
defparam \rsel2_l~11 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y37_N28
cycloneive_lcell_comb \rsel2_l~12 (
// Equation(s):
// \rsel2_l~12_combout  = (!idex_sRST2 & (plif_ifidinstr_l_18 & (!idex_sRST & Selector9)))

	.dataa(idex_sRST2),
	.datab(plif_ifidinstr_l_18),
	.datac(idex_sRST),
	.datad(Selector9),
	.cin(gnd),
	.combout(\rsel2_l~12_combout ),
	.cout());
// synopsys translate_off
defparam \rsel2_l~12 .lut_mask = 16'h0400;
defparam \rsel2_l~12 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y37_N22
cycloneive_lcell_comb \rsel2_l~13 (
// Equation(s):
// \rsel2_l~13_combout  = (!idex_sRST2 & (Selector9 & (!idex_sRST & plif_ifidinstr_l_19)))

	.dataa(idex_sRST2),
	.datab(Selector9),
	.datac(idex_sRST),
	.datad(plif_ifidinstr_l_19),
	.cin(gnd),
	.combout(\rsel2_l~13_combout ),
	.cout());
// synopsys translate_off
defparam \rsel2_l~13 .lut_mask = 16'h0400;
defparam \rsel2_l~13 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y37_N24
cycloneive_lcell_comb \rsel2_l~14 (
// Equation(s):
// \rsel2_l~14_combout  = (!idex_sRST2 & (plif_ifidinstr_l_20 & (!idex_sRST & Selector9)))

	.dataa(idex_sRST2),
	.datab(plif_ifidinstr_l_20),
	.datac(idex_sRST),
	.datad(Selector9),
	.cin(gnd),
	.combout(\rsel2_l~14_combout ),
	.cout());
// synopsys translate_off
defparam \rsel2_l~14 .lut_mask = 16'h0400;
defparam \rsel2_l~14 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X67_Y35_N24
cycloneive_lcell_comb \rdat2_l~0 (
// Equation(s):
// \rdat2_l~0_combout  = (!idex_sRST1 & ((Selector6 & ((Mux32))) # (!Selector6 & (Mux321))))

	.dataa(Mux321),
	.datab(Selector6),
	.datac(idex_sRST1),
	.datad(Mux32),
	.cin(gnd),
	.combout(\rdat2_l~0_combout ),
	.cout());
// synopsys translate_off
defparam \rdat2_l~0 .lut_mask = 16'h0E02;
defparam \rdat2_l~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y32_N30
cycloneive_lcell_comb \extimm_l~2 (
// Equation(s):
// \extimm_l~2_combout  = (\Equal0~0_combout  & !WideOr151)

	.dataa(gnd),
	.datab(Equal0),
	.datac(gnd),
	.datad(WideOr15),
	.cin(gnd),
	.combout(\extimm_l~2_combout ),
	.cout());
// synopsys translate_off
defparam \extimm_l~2 .lut_mask = 16'h00CC;
defparam \extimm_l~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y31_N12
cycloneive_lcell_comb \extimm_l~3 (
// Equation(s):
// \extimm_l~3_combout  = (!idex_sRST1 & ((\extimm[30]~0_combout ) # ((plif_ifidinstr_l_14 & \extimm_l~2_combout ))))

	.dataa(extimm_30),
	.datab(plif_ifidinstr_l_14),
	.datac(\extimm_l~2_combout ),
	.datad(idex_sRST1),
	.cin(gnd),
	.combout(\extimm_l~3_combout ),
	.cout());
// synopsys translate_off
defparam \extimm_l~3 .lut_mask = 16'h00EA;
defparam \extimm_l~3 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y39_N16
cycloneive_lcell_comb \rdat2_l~1 (
// Equation(s):
// \rdat2_l~1_combout  = (!idex_sRST1 & ((Selector6 & (Mux33)) # (!Selector6 & ((Mux331)))))

	.dataa(Selector6),
	.datab(Mux33),
	.datac(idex_sRST1),
	.datad(Mux331),
	.cin(gnd),
	.combout(\rdat2_l~1_combout ),
	.cout());
// synopsys translate_off
defparam \rdat2_l~1 .lut_mask = 16'h0D08;
defparam \rdat2_l~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y32_N4
cycloneive_lcell_comb \extimm_l~4 (
// Equation(s):
// \extimm_l~4_combout  = (!idex_sRST1 & ((\extimm[30]~0_combout ) # ((plif_ifidinstr_l_13 & \extimm_l~2_combout ))))

	.dataa(plif_ifidinstr_l_13),
	.datab(idex_sRST1),
	.datac(\extimm_l~2_combout ),
	.datad(extimm_30),
	.cin(gnd),
	.combout(\extimm_l~4_combout ),
	.cout());
// synopsys translate_off
defparam \extimm_l~4 .lut_mask = 16'h3320;
defparam \extimm_l~4 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y32_N8
cycloneive_lcell_comb \rdat2_l~2 (
// Equation(s):
// \rdat2_l~2_combout  = (!idex_sRST1 & ((Selector6 & (Mux34)) # (!Selector6 & ((Mux341)))))

	.dataa(Selector6),
	.datab(idex_sRST1),
	.datac(Mux34),
	.datad(Mux341),
	.cin(gnd),
	.combout(\rdat2_l~2_combout ),
	.cout());
// synopsys translate_off
defparam \rdat2_l~2 .lut_mask = 16'h3120;
defparam \rdat2_l~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y31_N30
cycloneive_lcell_comb \extimm_l~5 (
// Equation(s):
// \extimm_l~5_combout  = (!idex_sRST1 & ((\extimm[30]~0_combout ) # ((plif_ifidinstr_l_12 & \extimm_l~2_combout ))))

	.dataa(extimm_30),
	.datab(plif_ifidinstr_l_12),
	.datac(\extimm_l~2_combout ),
	.datad(idex_sRST1),
	.cin(gnd),
	.combout(\extimm_l~5_combout ),
	.cout());
// synopsys translate_off
defparam \extimm_l~5 .lut_mask = 16'h00EA;
defparam \extimm_l~5 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X67_Y35_N14
cycloneive_lcell_comb \rdat2_l~3 (
// Equation(s):
// \rdat2_l~3_combout  = (!idex_sRST1 & ((Selector6 & ((Mux35))) # (!Selector6 & (Mux351))))

	.dataa(Mux351),
	.datab(Selector6),
	.datac(idex_sRST1),
	.datad(Mux35),
	.cin(gnd),
	.combout(\rdat2_l~3_combout ),
	.cout());
// synopsys translate_off
defparam \rdat2_l~3 .lut_mask = 16'h0E02;
defparam \rdat2_l~3 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y32_N22
cycloneive_lcell_comb \extimm_l~6 (
// Equation(s):
// \extimm_l~6_combout  = (!idex_sRST1 & ((\extimm[30]~0_combout ) # ((plif_ifidinstr_l_11 & \extimm_l~2_combout ))))

	.dataa(plif_ifidinstr_l_11),
	.datab(idex_sRST1),
	.datac(\extimm_l~2_combout ),
	.datad(extimm_30),
	.cin(gnd),
	.combout(\extimm_l~6_combout ),
	.cout());
// synopsys translate_off
defparam \extimm_l~6 .lut_mask = 16'h3320;
defparam \extimm_l~6 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y39_N30
cycloneive_lcell_comb \rdat2_l~4 (
// Equation(s):
// \rdat2_l~4_combout  = (!idex_sRST1 & ((Selector6 & (Mux36)) # (!Selector6 & ((Mux361)))))

	.dataa(Selector6),
	.datab(Mux36),
	.datac(idex_sRST1),
	.datad(Mux361),
	.cin(gnd),
	.combout(\rdat2_l~4_combout ),
	.cout());
// synopsys translate_off
defparam \rdat2_l~4 .lut_mask = 16'h0D08;
defparam \rdat2_l~4 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y32_N24
cycloneive_lcell_comb \extimm_l~7 (
// Equation(s):
// \extimm_l~7_combout  = (!idex_sRST1 & ((\extimm[30]~0_combout ) # ((plif_ifidinstr_l_10 & \extimm_l~2_combout ))))

	.dataa(plif_ifidinstr_l_10),
	.datab(idex_sRST1),
	.datac(\extimm_l~2_combout ),
	.datad(extimm_30),
	.cin(gnd),
	.combout(\extimm_l~7_combout ),
	.cout());
// synopsys translate_off
defparam \extimm_l~7 .lut_mask = 16'h3320;
defparam \extimm_l~7 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y32_N22
cycloneive_lcell_comb \rdat2_l~5 (
// Equation(s):
// \rdat2_l~5_combout  = (!idex_sRST1 & ((Selector6 & ((Mux37))) # (!Selector6 & (Mux371))))

	.dataa(Selector6),
	.datab(idex_sRST1),
	.datac(Mux371),
	.datad(Mux37),
	.cin(gnd),
	.combout(\rdat2_l~5_combout ),
	.cout());
// synopsys translate_off
defparam \rdat2_l~5 .lut_mask = 16'h3210;
defparam \rdat2_l~5 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y32_N10
cycloneive_lcell_comb \extimm_l~8 (
// Equation(s):
// \extimm_l~8_combout  = (!idex_sRST1 & ((\extimm[30]~0_combout ) # ((plif_ifidinstr_l_9 & \extimm_l~2_combout ))))

	.dataa(plif_ifidinstr_l_9),
	.datab(idex_sRST1),
	.datac(\extimm_l~2_combout ),
	.datad(extimm_30),
	.cin(gnd),
	.combout(\extimm_l~8_combout ),
	.cout());
// synopsys translate_off
defparam \extimm_l~8 .lut_mask = 16'h3320;
defparam \extimm_l~8 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X65_Y32_N20
cycloneive_lcell_comb \rdat2_l~6 (
// Equation(s):
// \rdat2_l~6_combout  = (!idex_sRST1 & ((Selector6 & ((Mux38))) # (!Selector6 & (Mux381))))

	.dataa(Selector6),
	.datab(Mux381),
	.datac(idex_sRST1),
	.datad(Mux38),
	.cin(gnd),
	.combout(\rdat2_l~6_combout ),
	.cout());
// synopsys translate_off
defparam \rdat2_l~6 .lut_mask = 16'h0E04;
defparam \rdat2_l~6 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y32_N8
cycloneive_lcell_comb \extimm_l~9 (
// Equation(s):
// \extimm_l~9_combout  = (!idex_sRST1 & ((\extimm[30]~0_combout ) # ((plif_ifidinstr_l_8 & \extimm_l~2_combout ))))

	.dataa(plif_ifidinstr_l_8),
	.datab(idex_sRST1),
	.datac(\extimm_l~2_combout ),
	.datad(extimm_30),
	.cin(gnd),
	.combout(\extimm_l~9_combout ),
	.cout());
// synopsys translate_off
defparam \extimm_l~9 .lut_mask = 16'h3320;
defparam \extimm_l~9 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X65_Y32_N30
cycloneive_lcell_comb \rdat2_l~7 (
// Equation(s):
// \rdat2_l~7_combout  = (!idex_sRST1 & ((Selector6 & ((Mux39))) # (!Selector6 & (Mux391))))

	.dataa(idex_sRST1),
	.datab(Mux391),
	.datac(Selector6),
	.datad(Mux39),
	.cin(gnd),
	.combout(\rdat2_l~7_combout ),
	.cout());
// synopsys translate_off
defparam \rdat2_l~7 .lut_mask = 16'h5404;
defparam \rdat2_l~7 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y32_N6
cycloneive_lcell_comb \extimm_l~10 (
// Equation(s):
// \extimm_l~10_combout  = (!idex_sRST1 & ((\extimm[30]~0_combout ) # ((plif_ifidinstr_l_7 & \extimm_l~2_combout ))))

	.dataa(plif_ifidinstr_l_7),
	.datab(idex_sRST1),
	.datac(\extimm_l~2_combout ),
	.datad(extimm_30),
	.cin(gnd),
	.combout(\extimm_l~10_combout ),
	.cout());
// synopsys translate_off
defparam \extimm_l~10 .lut_mask = 16'h3320;
defparam \extimm_l~10 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X67_Y30_N24
cycloneive_lcell_comb \rdat2_l~8 (
// Equation(s):
// \rdat2_l~8_combout  = (!idex_sRST1 & ((Selector6 & (Mux40)) # (!Selector6 & ((Mux401)))))

	.dataa(Selector6),
	.datab(Mux40),
	.datac(idex_sRST1),
	.datad(Mux401),
	.cin(gnd),
	.combout(\rdat2_l~8_combout ),
	.cout());
// synopsys translate_off
defparam \rdat2_l~8 .lut_mask = 16'h0D08;
defparam \rdat2_l~8 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y32_N12
cycloneive_lcell_comb \extimm_l~11 (
// Equation(s):
// \extimm_l~11_combout  = (!idex_sRST1 & ((\extimm[30]~0_combout ) # ((\extimm_l~2_combout  & plif_ifidinstr_l_6))))

	.dataa(\extimm_l~2_combout ),
	.datab(idex_sRST1),
	.datac(plif_ifidinstr_l_6),
	.datad(extimm_30),
	.cin(gnd),
	.combout(\extimm_l~11_combout ),
	.cout());
// synopsys translate_off
defparam \extimm_l~11 .lut_mask = 16'h3320;
defparam \extimm_l~11 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X67_Y30_N14
cycloneive_lcell_comb \rdat2_l~9 (
// Equation(s):
// \rdat2_l~9_combout  = (!idex_sRST1 & ((Selector6 & ((Mux41))) # (!Selector6 & (Mux411))))

	.dataa(Mux411),
	.datab(Selector6),
	.datac(idex_sRST1),
	.datad(Mux41),
	.cin(gnd),
	.combout(\rdat2_l~9_combout ),
	.cout());
// synopsys translate_off
defparam \rdat2_l~9 .lut_mask = 16'h0E02;
defparam \rdat2_l~9 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y32_N2
cycloneive_lcell_comb \extimm_l~12 (
// Equation(s):
// \extimm_l~12_combout  = (!idex_sRST1 & ((\extimm[30]~0_combout ) # ((\extimm_l~2_combout  & plif_ifidinstr_l_5))))

	.dataa(\extimm_l~2_combout ),
	.datab(idex_sRST1),
	.datac(plif_ifidinstr_l_5),
	.datad(extimm_30),
	.cin(gnd),
	.combout(\extimm_l~12_combout ),
	.cout());
// synopsys translate_off
defparam \extimm_l~12 .lut_mask = 16'h3320;
defparam \extimm_l~12 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X67_Y30_N0
cycloneive_lcell_comb \rdat2_l~10 (
// Equation(s):
// \rdat2_l~10_combout  = (!idex_sRST1 & ((Selector6 & ((Mux42))) # (!Selector6 & (Mux421))))

	.dataa(idex_sRST1),
	.datab(Mux421),
	.datac(Selector6),
	.datad(Mux42),
	.cin(gnd),
	.combout(\rdat2_l~10_combout ),
	.cout());
// synopsys translate_off
defparam \rdat2_l~10 .lut_mask = 16'h5404;
defparam \rdat2_l~10 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y33_N28
cycloneive_lcell_comb \extimm_l~13 (
// Equation(s):
// \extimm_l~13_combout  = (!idex_sRST1 & ((\extimm[30]~0_combout ) # ((\Equal0~0_combout  & Selector14))))

	.dataa(Equal0),
	.datab(extimm_30),
	.datac(Selector14),
	.datad(idex_sRST1),
	.cin(gnd),
	.combout(\extimm_l~13_combout ),
	.cout());
// synopsys translate_off
defparam \extimm_l~13 .lut_mask = 16'h00EC;
defparam \extimm_l~13 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y39_N0
cycloneive_lcell_comb \rdat2_l~11 (
// Equation(s):
// \rdat2_l~11_combout  = (!idex_sRST1 & ((Selector6 & (Mux43)) # (!Selector6 & ((Mux431)))))

	.dataa(Mux43),
	.datab(Selector6),
	.datac(idex_sRST1),
	.datad(Mux431),
	.cin(gnd),
	.combout(\rdat2_l~11_combout ),
	.cout());
// synopsys translate_off
defparam \rdat2_l~11 .lut_mask = 16'h0B08;
defparam \rdat2_l~11 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y33_N26
cycloneive_lcell_comb \extimm_l~14 (
// Equation(s):
// \extimm_l~14_combout  = (!idex_sRST1 & ((\extimm[30]~0_combout ) # ((\Equal0~0_combout  & Selector15))))

	.dataa(Equal0),
	.datab(Selector15),
	.datac(idex_sRST1),
	.datad(extimm_30),
	.cin(gnd),
	.combout(\extimm_l~14_combout ),
	.cout());
// synopsys translate_off
defparam \extimm_l~14 .lut_mask = 16'h0F08;
defparam \extimm_l~14 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y39_N14
cycloneive_lcell_comb \rdat2_l~12 (
// Equation(s):
// \rdat2_l~12_combout  = (!idex_sRST1 & ((Selector6 & (Mux44)) # (!Selector6 & ((Mux441)))))

	.dataa(Selector6),
	.datab(Mux44),
	.datac(Mux441),
	.datad(idex_sRST1),
	.cin(gnd),
	.combout(\rdat2_l~12_combout ),
	.cout());
// synopsys translate_off
defparam \rdat2_l~12 .lut_mask = 16'h00D8;
defparam \rdat2_l~12 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y33_N18
cycloneive_lcell_comb \extimm_l~15 (
// Equation(s):
// \extimm_l~15_combout  = (!idex_sRST1 & ((\extimm[30]~0_combout ) # ((\Equal0~0_combout  & Selector16))))

	.dataa(extimm_30),
	.datab(Equal0),
	.datac(Selector16),
	.datad(idex_sRST1),
	.cin(gnd),
	.combout(\extimm_l~15_combout ),
	.cout());
// synopsys translate_off
defparam \extimm_l~15 .lut_mask = 16'h00EA;
defparam \extimm_l~15 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X63_Y39_N20
cycloneive_lcell_comb \rdat2_l~13 (
// Equation(s):
// \rdat2_l~13_combout  = (!idex_sRST1 & ((Selector6 & ((Mux45))) # (!Selector6 & (Mux451))))

	.dataa(Selector6),
	.datab(Mux451),
	.datac(idex_sRST1),
	.datad(Mux45),
	.cin(gnd),
	.combout(\rdat2_l~13_combout ),
	.cout());
// synopsys translate_off
defparam \rdat2_l~13 .lut_mask = 16'h0E04;
defparam \rdat2_l~13 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y31_N28
cycloneive_lcell_comb \extimm_l~16 (
// Equation(s):
// \extimm_l~16_combout  = (!idex_sRST1 & ((\extimm[30]~0_combout ) # ((\Equal0~0_combout  & Selector17))))

	.dataa(extimm_30),
	.datab(Equal0),
	.datac(Selector17),
	.datad(idex_sRST1),
	.cin(gnd),
	.combout(\extimm_l~16_combout ),
	.cout());
// synopsys translate_off
defparam \extimm_l~16 .lut_mask = 16'h00EA;
defparam \extimm_l~16 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X67_Y40_N24
cycloneive_lcell_comb \rdat2_l~14 (
// Equation(s):
// \rdat2_l~14_combout  = (!idex_sRST1 & ((Selector6 & ((Mux46))) # (!Selector6 & (Mux461))))

	.dataa(idex_sRST1),
	.datab(Selector6),
	.datac(Mux461),
	.datad(Mux46),
	.cin(gnd),
	.combout(\rdat2_l~14_combout ),
	.cout());
// synopsys translate_off
defparam \rdat2_l~14 .lut_mask = 16'h5410;
defparam \rdat2_l~14 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y31_N22
cycloneive_lcell_comb \extimm_l~17 (
// Equation(s):
// \extimm_l~17_combout  = (!idex_sRST1 & ((\extimm[30]~0_combout ) # ((\Equal0~0_combout  & Selector18))))

	.dataa(extimm_30),
	.datab(Equal0),
	.datac(Selector18),
	.datad(idex_sRST1),
	.cin(gnd),
	.combout(\extimm_l~17_combout ),
	.cout());
// synopsys translate_off
defparam \extimm_l~17 .lut_mask = 16'h00EA;
defparam \extimm_l~17 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X67_Y40_N2
cycloneive_lcell_comb \rdat2_l~15 (
// Equation(s):
// \rdat2_l~15_combout  = (!idex_sRST1 & ((Selector6 & ((Mux47))) # (!Selector6 & (Mux471))))

	.dataa(idex_sRST1),
	.datab(Selector6),
	.datac(Mux471),
	.datad(Mux47),
	.cin(gnd),
	.combout(\rdat2_l~15_combout ),
	.cout());
// synopsys translate_off
defparam \rdat2_l~15 .lut_mask = 16'h5410;
defparam \rdat2_l~15 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y30_N4
cycloneive_lcell_comb \extimm_l~18 (
// Equation(s):
// \extimm_l~18_combout  = (!idex_sRST & (!idex_sRST2 & (!WideOr151 & !\Equal0~0_combout )))

	.dataa(idex_sRST),
	.datab(idex_sRST2),
	.datac(WideOr15),
	.datad(Equal0),
	.cin(gnd),
	.combout(\extimm_l~18_combout ),
	.cout());
// synopsys translate_off
defparam \extimm_l~18 .lut_mask = 16'h0001;
defparam \extimm_l~18 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y30_N16
cycloneive_lcell_comb \extimm_l~19 (
// Equation(s):
// \extimm_l~19_combout  = (\extimm_l~18_combout  & plif_ifidinstr_l_15)

	.dataa(gnd),
	.datab(gnd),
	.datac(\extimm_l~18_combout ),
	.datad(plif_ifidinstr_l_15),
	.cin(gnd),
	.combout(\extimm_l~19_combout ),
	.cout());
// synopsys translate_off
defparam \extimm_l~19 .lut_mask = 16'hF000;
defparam \extimm_l~19 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X70_Y35_N24
cycloneive_lcell_comb \rdat2_l~16 (
// Equation(s):
// \rdat2_l~16_combout  = (!idex_sRST1 & ((Selector6 & ((Mux48))) # (!Selector6 & (Mux481))))

	.dataa(idex_sRST1),
	.datab(Selector6),
	.datac(Mux481),
	.datad(Mux48),
	.cin(gnd),
	.combout(\rdat2_l~16_combout ),
	.cout());
// synopsys translate_off
defparam \rdat2_l~16 .lut_mask = 16'h5410;
defparam \rdat2_l~16 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X66_Y30_N20
cycloneive_lcell_comb \rdat2_l~17 (
// Equation(s):
// \rdat2_l~17_combout  = (!idex_sRST1 & ((Selector6 & ((Mux49))) # (!Selector6 & (Mux491))))

	.dataa(Mux491),
	.datab(Selector6),
	.datac(Mux49),
	.datad(idex_sRST1),
	.cin(gnd),
	.combout(\rdat2_l~17_combout ),
	.cout());
// synopsys translate_off
defparam \rdat2_l~17 .lut_mask = 16'h00E2;
defparam \rdat2_l~17 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y30_N14
cycloneive_lcell_comb \extimm_l~20 (
// Equation(s):
// \extimm_l~20_combout  = (plif_ifidinstr_l_14 & \extimm_l~18_combout )

	.dataa(plif_ifidinstr_l_14),
	.datab(gnd),
	.datac(\extimm_l~18_combout ),
	.datad(gnd),
	.cin(gnd),
	.combout(\extimm_l~20_combout ),
	.cout());
// synopsys translate_off
defparam \extimm_l~20 .lut_mask = 16'hA0A0;
defparam \extimm_l~20 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y30_N8
cycloneive_lcell_comb \extimm_l~21 (
// Equation(s):
// \extimm_l~21_combout  = (\extimm_l~18_combout  & plif_ifidinstr_l_13)

	.dataa(gnd),
	.datab(gnd),
	.datac(\extimm_l~18_combout ),
	.datad(plif_ifidinstr_l_13),
	.cin(gnd),
	.combout(\extimm_l~21_combout ),
	.cout());
// synopsys translate_off
defparam \extimm_l~21 .lut_mask = 16'hF000;
defparam \extimm_l~21 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y38_N10
cycloneive_lcell_comb \rdat2_l~18 (
// Equation(s):
// \rdat2_l~18_combout  = (!idex_sRST1 & ((Selector6 & ((Mux50))) # (!Selector6 & (Mux501))))

	.dataa(idex_sRST1),
	.datab(Selector6),
	.datac(Mux501),
	.datad(Mux50),
	.cin(gnd),
	.combout(\rdat2_l~18_combout ),
	.cout());
// synopsys translate_off
defparam \rdat2_l~18 .lut_mask = 16'h5410;
defparam \rdat2_l~18 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y30_N24
cycloneive_lcell_comb \rdat2_l~19 (
// Equation(s):
// \rdat2_l~19_combout  = (!idex_sRST1 & ((Selector6 & ((Mux51))) # (!Selector6 & (Mux511))))

	.dataa(Mux511),
	.datab(idex_sRST1),
	.datac(Selector6),
	.datad(Mux51),
	.cin(gnd),
	.combout(\rdat2_l~19_combout ),
	.cout());
// synopsys translate_off
defparam \rdat2_l~19 .lut_mask = 16'h3202;
defparam \rdat2_l~19 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y30_N18
cycloneive_lcell_comb \extimm_l~22 (
// Equation(s):
// \extimm_l~22_combout  = (\extimm_l~18_combout  & plif_ifidinstr_l_12)

	.dataa(gnd),
	.datab(gnd),
	.datac(\extimm_l~18_combout ),
	.datad(plif_ifidinstr_l_12),
	.cin(gnd),
	.combout(\extimm_l~22_combout ),
	.cout());
// synopsys translate_off
defparam \extimm_l~22 .lut_mask = 16'hF000;
defparam \extimm_l~22 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y30_N24
cycloneive_lcell_comb \extimm_l~23 (
// Equation(s):
// \extimm_l~23_combout  = (\extimm_l~18_combout  & plif_ifidinstr_l_11)

	.dataa(gnd),
	.datab(gnd),
	.datac(\extimm_l~18_combout ),
	.datad(plif_ifidinstr_l_11),
	.cin(gnd),
	.combout(\extimm_l~23_combout ),
	.cout());
// synopsys translate_off
defparam \extimm_l~23 .lut_mask = 16'hF000;
defparam \extimm_l~23 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y38_N2
cycloneive_lcell_comb \rdat2_l~20 (
// Equation(s):
// \rdat2_l~20_combout  = (!idex_sRST1 & ((Selector6 & (Mux52)) # (!Selector6 & ((Mux521)))))

	.dataa(Selector6),
	.datab(idex_sRST1),
	.datac(Mux52),
	.datad(Mux521),
	.cin(gnd),
	.combout(\rdat2_l~20_combout ),
	.cout());
// synopsys translate_off
defparam \rdat2_l~20 .lut_mask = 16'h3120;
defparam \rdat2_l~20 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X68_Y40_N20
cycloneive_lcell_comb \rdat2_l~21 (
// Equation(s):
// \rdat2_l~21_combout  = (!idex_sRST1 & ((Selector6 & ((Mux53))) # (!Selector6 & (Mux531))))

	.dataa(Mux531),
	.datab(Selector6),
	.datac(Mux53),
	.datad(idex_sRST1),
	.cin(gnd),
	.combout(\rdat2_l~21_combout ),
	.cout());
// synopsys translate_off
defparam \rdat2_l~21 .lut_mask = 16'h00E2;
defparam \rdat2_l~21 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y30_N6
cycloneive_lcell_comb \extimm_l~24 (
// Equation(s):
// \extimm_l~24_combout  = (\extimm_l~18_combout  & plif_ifidinstr_l_10)

	.dataa(gnd),
	.datab(gnd),
	.datac(\extimm_l~18_combout ),
	.datad(plif_ifidinstr_l_10),
	.cin(gnd),
	.combout(\extimm_l~24_combout ),
	.cout());
// synopsys translate_off
defparam \extimm_l~24 .lut_mask = 16'hF000;
defparam \extimm_l~24 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y30_N20
cycloneive_lcell_comb \extimm_l~25 (
// Equation(s):
// \extimm_l~25_combout  = (plif_ifidinstr_l_9 & \extimm_l~18_combout )

	.dataa(gnd),
	.datab(plif_ifidinstr_l_9),
	.datac(\extimm_l~18_combout ),
	.datad(gnd),
	.cin(gnd),
	.combout(\extimm_l~25_combout ),
	.cout());
// synopsys translate_off
defparam \extimm_l~25 .lut_mask = 16'hC0C0;
defparam \extimm_l~25 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X68_Y40_N30
cycloneive_lcell_comb \rdat2_l~22 (
// Equation(s):
// \rdat2_l~22_combout  = (!idex_sRST1 & ((Selector6 & ((Mux54))) # (!Selector6 & (Mux541))))

	.dataa(Selector6),
	.datab(idex_sRST1),
	.datac(Mux541),
	.datad(Mux54),
	.cin(gnd),
	.combout(\rdat2_l~22_combout ),
	.cout());
// synopsys translate_off
defparam \rdat2_l~22 .lut_mask = 16'h3210;
defparam \rdat2_l~22 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y36_N24
cycloneive_lcell_comb \rdat2_l~23 (
// Equation(s):
// \rdat2_l~23_combout  = (!idex_sRST1 & ((Selector6 & (Mux55)) # (!Selector6 & ((Mux551)))))

	.dataa(Selector6),
	.datab(idex_sRST1),
	.datac(Mux55),
	.datad(Mux551),
	.cin(gnd),
	.combout(\rdat2_l~23_combout ),
	.cout());
// synopsys translate_off
defparam \rdat2_l~23 .lut_mask = 16'h3120;
defparam \rdat2_l~23 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y30_N22
cycloneive_lcell_comb \extimm_l~26 (
// Equation(s):
// \extimm_l~26_combout  = (plif_ifidinstr_l_8 & \extimm_l~18_combout )

	.dataa(plif_ifidinstr_l_8),
	.datab(gnd),
	.datac(\extimm_l~18_combout ),
	.datad(gnd),
	.cin(gnd),
	.combout(\extimm_l~26_combout ),
	.cout());
// synopsys translate_off
defparam \extimm_l~26 .lut_mask = 16'hA0A0;
defparam \extimm_l~26 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y30_N0
cycloneive_lcell_comb \extimm_l~27 (
// Equation(s):
// \extimm_l~27_combout  = (plif_ifidinstr_l_7 & \extimm_l~18_combout )

	.dataa(plif_ifidinstr_l_7),
	.datab(gnd),
	.datac(\extimm_l~18_combout ),
	.datad(gnd),
	.cin(gnd),
	.combout(\extimm_l~27_combout ),
	.cout());
// synopsys translate_off
defparam \extimm_l~27 .lut_mask = 16'hA0A0;
defparam \extimm_l~27 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y38_N22
cycloneive_lcell_comb \rdat2_l~24 (
// Equation(s):
// \rdat2_l~24_combout  = (!idex_sRST1 & ((Selector6 & (Mux56)) # (!Selector6 & ((Mux561)))))

	.dataa(Selector6),
	.datab(idex_sRST1),
	.datac(Mux56),
	.datad(Mux561),
	.cin(gnd),
	.combout(\rdat2_l~24_combout ),
	.cout());
// synopsys translate_off
defparam \rdat2_l~24 .lut_mask = 16'h3120;
defparam \rdat2_l~24 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X65_Y30_N20
cycloneive_lcell_comb \rdat2_l~25 (
// Equation(s):
// \rdat2_l~25_combout  = (!idex_sRST1 & ((Selector6 & ((Mux57))) # (!Selector6 & (Mux571))))

	.dataa(Mux571),
	.datab(Selector6),
	.datac(idex_sRST1),
	.datad(Mux57),
	.cin(gnd),
	.combout(\rdat2_l~25_combout ),
	.cout());
// synopsys translate_off
defparam \rdat2_l~25 .lut_mask = 16'h0E02;
defparam \rdat2_l~25 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y30_N2
cycloneive_lcell_comb \extimm_l~28 (
// Equation(s):
// \extimm_l~28_combout  = (plif_ifidinstr_l_6 & \extimm_l~18_combout )

	.dataa(gnd),
	.datab(plif_ifidinstr_l_6),
	.datac(\extimm_l~18_combout ),
	.datad(gnd),
	.cin(gnd),
	.combout(\extimm_l~28_combout ),
	.cout());
// synopsys translate_off
defparam \extimm_l~28 .lut_mask = 16'hC0C0;
defparam \extimm_l~28 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y30_N28
cycloneive_lcell_comb \extimm_l~29 (
// Equation(s):
// \extimm_l~29_combout  = (plif_ifidinstr_l_5 & \extimm_l~18_combout )

	.dataa(plif_ifidinstr_l_5),
	.datab(gnd),
	.datac(\extimm_l~18_combout ),
	.datad(gnd),
	.cin(gnd),
	.combout(\extimm_l~29_combout ),
	.cout());
// synopsys translate_off
defparam \extimm_l~29 .lut_mask = 16'hA0A0;
defparam \extimm_l~29 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X65_Y30_N22
cycloneive_lcell_comb \rdat2_l~26 (
// Equation(s):
// \rdat2_l~26_combout  = (!idex_sRST1 & ((Selector6 & ((Mux58))) # (!Selector6 & (Mux581))))

	.dataa(Mux581),
	.datab(Selector6),
	.datac(idex_sRST1),
	.datad(Mux58),
	.cin(gnd),
	.combout(\rdat2_l~26_combout ),
	.cout());
// synopsys translate_off
defparam \rdat2_l~26 .lut_mask = 16'h0E02;
defparam \rdat2_l~26 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y37_N12
cycloneive_lcell_comb \rsel1_l~10 (
// Equation(s):
// \rsel1_l~10_combout  = (plif_ifidinstr_l_25 & (!idex_sRST2 & (Selector4 & !idex_sRST)))

	.dataa(plif_ifidinstr_l_25),
	.datab(idex_sRST2),
	.datac(Selector4),
	.datad(idex_sRST),
	.cin(gnd),
	.combout(\rsel1_l~10_combout ),
	.cout());
// synopsys translate_off
defparam \rsel1_l~10 .lut_mask = 16'h0020;
defparam \rsel1_l~10 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y37_N8
cycloneive_lcell_comb \rsel1_l~11 (
// Equation(s):
// \rsel1_l~11_combout  = (plif_ifidinstr_l_22 & (!idex_sRST2 & (Selector4 & !idex_sRST)))

	.dataa(plif_ifidinstr_l_22),
	.datab(idex_sRST2),
	.datac(Selector4),
	.datad(idex_sRST),
	.cin(gnd),
	.combout(\rsel1_l~11_combout ),
	.cout());
// synopsys translate_off
defparam \rsel1_l~11 .lut_mask = 16'h0020;
defparam \rsel1_l~11 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y37_N6
cycloneive_lcell_comb \rsel1_l~12 (
// Equation(s):
// \rsel1_l~12_combout  = (Selector4 & (!idex_sRST2 & (plif_ifidinstr_l_21 & !idex_sRST)))

	.dataa(Selector4),
	.datab(idex_sRST2),
	.datac(plif_ifidinstr_l_21),
	.datad(idex_sRST),
	.cin(gnd),
	.combout(\rsel1_l~12_combout ),
	.cout());
// synopsys translate_off
defparam \rsel1_l~12 .lut_mask = 16'h0020;
defparam \rsel1_l~12 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y37_N18
cycloneive_lcell_comb \rsel1_l~13 (
// Equation(s):
// \rsel1_l~13_combout  = (plif_ifidinstr_l_23 & (!idex_sRST2 & (Selector4 & !idex_sRST)))

	.dataa(plif_ifidinstr_l_23),
	.datab(idex_sRST2),
	.datac(Selector4),
	.datad(idex_sRST),
	.cin(gnd),
	.combout(\rsel1_l~13_combout ),
	.cout());
// synopsys translate_off
defparam \rsel1_l~13 .lut_mask = 16'h0020;
defparam \rsel1_l~13 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y37_N24
cycloneive_lcell_comb \rsel1_l~14 (
// Equation(s):
// \rsel1_l~14_combout  = (Selector4 & (!idex_sRST & (!idex_sRST2 & plif_ifidinstr_l_24)))

	.dataa(Selector4),
	.datab(idex_sRST),
	.datac(idex_sRST2),
	.datad(plif_ifidinstr_l_24),
	.cin(gnd),
	.combout(\rsel1_l~14_combout ),
	.cout());
// synopsys translate_off
defparam \rsel1_l~14 .lut_mask = 16'h0200;
defparam \rsel1_l~14 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X63_Y32_N4
cycloneive_lcell_comb \rdat1_l~0 (
// Equation(s):
// \rdat1_l~0_combout  = (!idex_sRST1 & ((Selector1 & (Mux29)) # (!Selector1 & ((Mux291)))))

	.dataa(Selector1),
	.datab(Mux29),
	.datac(Mux291),
	.datad(idex_sRST1),
	.cin(gnd),
	.combout(\rdat1_l~0_combout ),
	.cout());
// synopsys translate_off
defparam \rdat1_l~0 .lut_mask = 16'h00D8;
defparam \rdat1_l~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X65_Y31_N24
cycloneive_lcell_comb \rdat1_l~1 (
// Equation(s):
// \rdat1_l~1_combout  = (!idex_sRST1 & ((Selector1 & (Mux30)) # (!Selector1 & ((Mux301)))))

	.dataa(Selector1),
	.datab(Mux30),
	.datac(Mux301),
	.datad(idex_sRST1),
	.cin(gnd),
	.combout(\rdat1_l~1_combout ),
	.cout());
// synopsys translate_off
defparam \rdat1_l~1 .lut_mask = 16'h00D8;
defparam \rdat1_l~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y35_N24
cycloneive_lcell_comb \rdat2_l~27 (
// Equation(s):
// \rdat2_l~27_combout  = (!idex_sRST1 & ((Selector6 & ((Mux63))) # (!Selector6 & (Mux631))))

	.dataa(idex_sRST1),
	.datab(Selector6),
	.datac(Mux631),
	.datad(Mux63),
	.cin(gnd),
	.combout(\rdat2_l~27_combout ),
	.cout());
// synopsys translate_off
defparam \rdat2_l~27 .lut_mask = 16'h5410;
defparam \rdat2_l~27 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y33_N8
cycloneive_lcell_comb \extimm_l~30 (
// Equation(s):
// \extimm_l~30_combout  = (!idex_sRST & (!\Equal0~0_combout  & (Selector18 & !idex_sRST2)))

	.dataa(idex_sRST),
	.datab(Equal0),
	.datac(Selector18),
	.datad(idex_sRST2),
	.cin(gnd),
	.combout(\extimm_l~30_combout ),
	.cout());
// synopsys translate_off
defparam \extimm_l~30 .lut_mask = 16'h0010;
defparam \extimm_l~30 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y37_N20
cycloneive_lcell_comb \extimm_l~31 (
// Equation(s):
// \extimm_l~31_combout  = (!\Equal0~0_combout  & (Selector17 & (!idex_sRST & !idex_sRST2)))

	.dataa(Equal0),
	.datab(Selector17),
	.datac(idex_sRST),
	.datad(idex_sRST2),
	.cin(gnd),
	.combout(\extimm_l~31_combout ),
	.cout());
// synopsys translate_off
defparam \extimm_l~31 .lut_mask = 16'h0004;
defparam \extimm_l~31 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y35_N10
cycloneive_lcell_comb \rdat2_l~28 (
// Equation(s):
// \rdat2_l~28_combout  = (!idex_sRST1 & ((Selector6 & ((Mux62))) # (!Selector6 & (Mux621))))

	.dataa(idex_sRST1),
	.datab(Selector6),
	.datac(Mux621),
	.datad(Mux62),
	.cin(gnd),
	.combout(\rdat2_l~28_combout ),
	.cout());
// synopsys translate_off
defparam \rdat2_l~28 .lut_mask = 16'h5410;
defparam \rdat2_l~28 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y34_N0
cycloneive_lcell_comb \rdat1_l~2 (
// Equation(s):
// \rdat1_l~2_combout  = (!idex_sRST1 & ((Selector1 & ((Mux27))) # (!Selector1 & (Mux271))))

	.dataa(Mux271),
	.datab(Selector1),
	.datac(idex_sRST1),
	.datad(Mux27),
	.cin(gnd),
	.combout(\rdat1_l~2_combout ),
	.cout());
// synopsys translate_off
defparam \rdat1_l~2 .lut_mask = 16'h0E02;
defparam \rdat1_l~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X70_Y37_N24
cycloneive_lcell_comb \rdat1_l~3 (
// Equation(s):
// \rdat1_l~3_combout  = (!idex_sRST1 & ((Selector1 & ((Mux28))) # (!Selector1 & (Mux281))))

	.dataa(Mux281),
	.datab(Selector1),
	.datac(Mux28),
	.datad(idex_sRST1),
	.cin(gnd),
	.combout(\rdat1_l~3_combout ),
	.cout());
// synopsys translate_off
defparam \rdat1_l~3 .lut_mask = 16'h00E2;
defparam \rdat1_l~3 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y35_N28
cycloneive_lcell_comb \rdat2_l~29 (
// Equation(s):
// \rdat2_l~29_combout  = (!idex_sRST1 & ((Selector6 & (Mux61)) # (!Selector6 & ((Mux611)))))

	.dataa(idex_sRST1),
	.datab(Selector6),
	.datac(Mux61),
	.datad(Mux611),
	.cin(gnd),
	.combout(\rdat2_l~29_combout ),
	.cout());
// synopsys translate_off
defparam \rdat2_l~29 .lut_mask = 16'h5140;
defparam \rdat2_l~29 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y36_N10
cycloneive_lcell_comb \extimm_l~32 (
// Equation(s):
// \extimm_l~32_combout  = (Selector16 & (!idex_sRST2 & (!\Equal0~0_combout  & !idex_sRST)))

	.dataa(Selector16),
	.datab(idex_sRST2),
	.datac(Equal0),
	.datad(idex_sRST),
	.cin(gnd),
	.combout(\extimm_l~32_combout ),
	.cout());
// synopsys translate_off
defparam \extimm_l~32 .lut_mask = 16'h0002;
defparam \extimm_l~32 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X68_Y36_N20
cycloneive_lcell_comb \rdat1_l~4 (
// Equation(s):
// \rdat1_l~4_combout  = (!idex_sRST1 & ((Selector1 & ((Mux23))) # (!Selector1 & (Mux231))))

	.dataa(idex_sRST1),
	.datab(Selector1),
	.datac(Mux231),
	.datad(Mux23),
	.cin(gnd),
	.combout(\rdat1_l~4_combout ),
	.cout());
// synopsys translate_off
defparam \rdat1_l~4 .lut_mask = 16'h5410;
defparam \rdat1_l~4 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y40_N28
cycloneive_lcell_comb \rdat1_l~5 (
// Equation(s):
// \rdat1_l~5_combout  = (!idex_sRST1 & ((Selector1 & ((Mux24))) # (!Selector1 & (Mux241))))

	.dataa(Selector1),
	.datab(idex_sRST1),
	.datac(Mux241),
	.datad(Mux24),
	.cin(gnd),
	.combout(\rdat1_l~5_combout ),
	.cout());
// synopsys translate_off
defparam \rdat1_l~5 .lut_mask = 16'h3210;
defparam \rdat1_l~5 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X67_Y36_N16
cycloneive_lcell_comb \rdat1_l~6 (
// Equation(s):
// \rdat1_l~6_combout  = (!idex_sRST1 & ((Selector1 & (Mux25)) # (!Selector1 & ((Mux251)))))

	.dataa(Selector1),
	.datab(idex_sRST1),
	.datac(Mux25),
	.datad(Mux251),
	.cin(gnd),
	.combout(\rdat1_l~6_combout ),
	.cout());
// synopsys translate_off
defparam \rdat1_l~6 .lut_mask = 16'h3120;
defparam \rdat1_l~6 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X67_Y36_N26
cycloneive_lcell_comb \rdat1_l~7 (
// Equation(s):
// \rdat1_l~7_combout  = (!idex_sRST1 & ((Selector1 & (Mux26)) # (!Selector1 & ((Mux261)))))

	.dataa(Selector1),
	.datab(idex_sRST1),
	.datac(Mux26),
	.datad(Mux261),
	.cin(gnd),
	.combout(\rdat1_l~7_combout ),
	.cout());
// synopsys translate_off
defparam \rdat1_l~7 .lut_mask = 16'h3120;
defparam \rdat1_l~7 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y36_N28
cycloneive_lcell_comb \extimm_l~33 (
// Equation(s):
// \extimm_l~33_combout  = (Selector15 & (!idex_sRST2 & (!\Equal0~0_combout  & !idex_sRST)))

	.dataa(Selector15),
	.datab(idex_sRST2),
	.datac(Equal0),
	.datad(idex_sRST),
	.cin(gnd),
	.combout(\extimm_l~33_combout ),
	.cout());
// synopsys translate_off
defparam \extimm_l~33 .lut_mask = 16'h0002;
defparam \extimm_l~33 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y36_N2
cycloneive_lcell_comb \rdat2_l~30 (
// Equation(s):
// \rdat2_l~30_combout  = (!idex_sRST1 & ((Selector6 & ((Mux60))) # (!Selector6 & (Mux601))))

	.dataa(Mux601),
	.datab(idex_sRST1),
	.datac(Selector6),
	.datad(Mux60),
	.cin(gnd),
	.combout(\rdat2_l~30_combout ),
	.cout());
// synopsys translate_off
defparam \rdat2_l~30 .lut_mask = 16'h3202;
defparam \rdat2_l~30 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X63_Y36_N0
cycloneive_lcell_comb \rdat1_l~8 (
// Equation(s):
// \rdat1_l~8_combout  = (!idex_sRST1 & ((Selector1 & (Mux15)) # (!Selector1 & ((Mux151)))))

	.dataa(idex_sRST1),
	.datab(Mux15),
	.datac(Selector1),
	.datad(Mux151),
	.cin(gnd),
	.combout(\rdat1_l~8_combout ),
	.cout());
// synopsys translate_off
defparam \rdat1_l~8 .lut_mask = 16'h4540;
defparam \rdat1_l~8 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y40_N22
cycloneive_lcell_comb \rdat1_l~9 (
// Equation(s):
// \rdat1_l~9_combout  = (!idex_sRST1 & ((Selector1 & (Mux16)) # (!Selector1 & ((Mux161)))))

	.dataa(idex_sRST1),
	.datab(Selector1),
	.datac(Mux16),
	.datad(Mux161),
	.cin(gnd),
	.combout(\rdat1_l~9_combout ),
	.cout());
// synopsys translate_off
defparam \rdat1_l~9 .lut_mask = 16'h5140;
defparam \rdat1_l~9 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X66_Y30_N14
cycloneive_lcell_comb \rdat1_l~10 (
// Equation(s):
// \rdat1_l~10_combout  = (!idex_sRST1 & ((Selector1 & (Mux17)) # (!Selector1 & ((Mux171)))))

	.dataa(idex_sRST1),
	.datab(Selector1),
	.datac(Mux17),
	.datad(Mux171),
	.cin(gnd),
	.combout(\rdat1_l~10_combout ),
	.cout());
// synopsys translate_off
defparam \rdat1_l~10 .lut_mask = 16'h5140;
defparam \rdat1_l~10 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X63_Y38_N4
cycloneive_lcell_comb \rdat1_l~11 (
// Equation(s):
// \rdat1_l~11_combout  = (!idex_sRST1 & ((Selector1 & ((Mux18))) # (!Selector1 & (Mux181))))

	.dataa(Mux181),
	.datab(Selector1),
	.datac(idex_sRST1),
	.datad(Mux18),
	.cin(gnd),
	.combout(\rdat1_l~11_combout ),
	.cout());
// synopsys translate_off
defparam \rdat1_l~11 .lut_mask = 16'h0E02;
defparam \rdat1_l~11 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y30_N2
cycloneive_lcell_comb \rdat1_l~12 (
// Equation(s):
// \rdat1_l~12_combout  = (!idex_sRST1 & ((Selector1 & ((Mux19))) # (!Selector1 & (Mux191))))

	.dataa(Selector1),
	.datab(idex_sRST1),
	.datac(Mux191),
	.datad(Mux19),
	.cin(gnd),
	.combout(\rdat1_l~12_combout ),
	.cout());
// synopsys translate_off
defparam \rdat1_l~12 .lut_mask = 16'h3210;
defparam \rdat1_l~12 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X63_Y38_N18
cycloneive_lcell_comb \rdat1_l~13 (
// Equation(s):
// \rdat1_l~13_combout  = (!idex_sRST1 & ((Selector1 & ((Mux20))) # (!Selector1 & (Mux201))))

	.dataa(Mux201),
	.datab(Selector1),
	.datac(idex_sRST1),
	.datad(Mux20),
	.cin(gnd),
	.combout(\rdat1_l~13_combout ),
	.cout());
// synopsys translate_off
defparam \rdat1_l~13 .lut_mask = 16'h0E02;
defparam \rdat1_l~13 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X70_Y36_N4
cycloneive_lcell_comb \rdat1_l~14 (
// Equation(s):
// \rdat1_l~14_combout  = (!idex_sRST1 & ((Selector1 & ((Mux21))) # (!Selector1 & (Mux211))))

	.dataa(Selector1),
	.datab(Mux211),
	.datac(Mux21),
	.datad(idex_sRST1),
	.cin(gnd),
	.combout(\rdat1_l~14_combout ),
	.cout());
// synopsys translate_off
defparam \rdat1_l~14 .lut_mask = 16'h00E4;
defparam \rdat1_l~14 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y41_N12
cycloneive_lcell_comb \rdat1_l~15 (
// Equation(s):
// \rdat1_l~15_combout  = (!idex_sRST1 & ((Selector1 & ((Mux22))) # (!Selector1 & (Mux221))))

	.dataa(Selector1),
	.datab(idex_sRST1),
	.datac(Mux221),
	.datad(Mux22),
	.cin(gnd),
	.combout(\rdat1_l~15_combout ),
	.cout());
// synopsys translate_off
defparam \rdat1_l~15 .lut_mask = 16'h3210;
defparam \rdat1_l~15 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y41_N14
cycloneive_lcell_comb \rdat2_l~31 (
// Equation(s):
// \rdat2_l~31_combout  = (!idex_sRST1 & ((Selector6 & ((Mux59))) # (!Selector6 & (Mux591))))

	.dataa(Selector6),
	.datab(idex_sRST1),
	.datac(Mux591),
	.datad(Mux59),
	.cin(gnd),
	.combout(\rdat2_l~31_combout ),
	.cout());
// synopsys translate_off
defparam \rdat2_l~31 .lut_mask = 16'h3210;
defparam \rdat2_l~31 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y41_N4
cycloneive_lcell_comb \extimm_l~34 (
// Equation(s):
// \extimm_l~34_combout  = (!\Equal0~0_combout  & (Selector14 & (!idex_sRST2 & !idex_sRST)))

	.dataa(Equal0),
	.datab(Selector14),
	.datac(idex_sRST2),
	.datad(idex_sRST),
	.cin(gnd),
	.combout(\extimm_l~34_combout ),
	.cout());
// synopsys translate_off
defparam \extimm_l~34 .lut_mask = 16'h0004;
defparam \extimm_l~34 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y41_N20
cycloneive_lcell_comb \plif_idex.extimm_l[4]~feeder (
// Equation(s):
// \plif_idex.extimm_l[4]~feeder_combout  = \extimm_l~34_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(\extimm_l~34_combout ),
	.cin(gnd),
	.combout(\plif_idex.extimm_l[4]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \plif_idex.extimm_l[4]~feeder .lut_mask = 16'hFF00;
defparam \plif_idex.extimm_l[4]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y33_N24
cycloneive_lcell_comb \rdat1_l~16 (
// Equation(s):
// \rdat1_l~16_combout  = (!idex_sRST1 & ((Selector1 & ((Mux0))) # (!Selector1 & (Mux01))))

	.dataa(Selector1),
	.datab(idex_sRST1),
	.datac(Mux01),
	.datad(Mux0),
	.cin(gnd),
	.combout(\rdat1_l~16_combout ),
	.cout());
// synopsys translate_off
defparam \rdat1_l~16 .lut_mask = 16'h3210;
defparam \rdat1_l~16 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y33_N2
cycloneive_lcell_comb \rdat1_l~17 (
// Equation(s):
// \rdat1_l~17_combout  = (!idex_sRST1 & ((Selector1 & (Mux2)) # (!Selector1 & ((Mux210)))))

	.dataa(Selector1),
	.datab(Mux2),
	.datac(idex_sRST1),
	.datad(Mux210),
	.cin(gnd),
	.combout(\rdat1_l~17_combout ),
	.cout());
// synopsys translate_off
defparam \rdat1_l~17 .lut_mask = 16'h0D08;
defparam \rdat1_l~17 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y33_N8
cycloneive_lcell_comb \rdat1_l~18 (
// Equation(s):
// \rdat1_l~18_combout  = (!idex_sRST1 & ((Selector1 & (Mux1)) # (!Selector1 & ((Mux11)))))

	.dataa(Selector1),
	.datab(idex_sRST1),
	.datac(Mux1),
	.datad(Mux11),
	.cin(gnd),
	.combout(\rdat1_l~18_combout ),
	.cout());
// synopsys translate_off
defparam \rdat1_l~18 .lut_mask = 16'h3120;
defparam \rdat1_l~18 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X63_Y39_N26
cycloneive_lcell_comb \rdat1_l~19 (
// Equation(s):
// \rdat1_l~19_combout  = (!idex_sRST1 & ((Selector1 & ((Mux3))) # (!Selector1 & (Mux31))))

	.dataa(Selector1),
	.datab(idex_sRST1),
	.datac(Mux31),
	.datad(Mux3),
	.cin(gnd),
	.combout(\rdat1_l~19_combout ),
	.cout());
// synopsys translate_off
defparam \rdat1_l~19 .lut_mask = 16'h3210;
defparam \rdat1_l~19 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X63_Y39_N4
cycloneive_lcell_comb \rdat1_l~20 (
// Equation(s):
// \rdat1_l~20_combout  = (!idex_sRST1 & ((Selector1 & (Mux4)) # (!Selector1 & ((Mux410)))))

	.dataa(Selector1),
	.datab(Mux4),
	.datac(idex_sRST1),
	.datad(Mux410),
	.cin(gnd),
	.combout(\rdat1_l~20_combout ),
	.cout());
// synopsys translate_off
defparam \rdat1_l~20 .lut_mask = 16'h0D08;
defparam \rdat1_l~20 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X63_Y32_N6
cycloneive_lcell_comb \rdat1_l~21 (
// Equation(s):
// \rdat1_l~21_combout  = (!idex_sRST1 & ((Selector1 & (Mux5)) # (!Selector1 & ((Mux510)))))

	.dataa(Selector1),
	.datab(Mux5),
	.datac(Mux510),
	.datad(idex_sRST1),
	.cin(gnd),
	.combout(\rdat1_l~21_combout ),
	.cout());
// synopsys translate_off
defparam \rdat1_l~21 .lut_mask = 16'h00D8;
defparam \rdat1_l~21 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X65_Y31_N14
cycloneive_lcell_comb \rdat1_l~22 (
// Equation(s):
// \rdat1_l~22_combout  = (!idex_sRST1 & ((Selector1 & ((Mux6))) # (!Selector1 & (Mux64))))

	.dataa(Selector1),
	.datab(idex_sRST1),
	.datac(Mux64),
	.datad(Mux6),
	.cin(gnd),
	.combout(\rdat1_l~22_combout ),
	.cout());
// synopsys translate_off
defparam \rdat1_l~22 .lut_mask = 16'h3210;
defparam \rdat1_l~22 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y34_N22
cycloneive_lcell_comb \rdat1_l~23 (
// Equation(s):
// \rdat1_l~23_combout  = (!idex_sRST1 & ((Selector1 & ((Mux7))) # (!Selector1 & (Mux71))))

	.dataa(idex_sRST1),
	.datab(Selector1),
	.datac(Mux71),
	.datad(Mux7),
	.cin(gnd),
	.combout(\rdat1_l~23_combout ),
	.cout());
// synopsys translate_off
defparam \rdat1_l~23 .lut_mask = 16'h5410;
defparam \rdat1_l~23 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X70_Y37_N10
cycloneive_lcell_comb \rdat1_l~24 (
// Equation(s):
// \rdat1_l~24_combout  = (!idex_sRST1 & ((Selector1 & (Mux8)) # (!Selector1 & ((Mux81)))))

	.dataa(Mux8),
	.datab(Selector1),
	.datac(Mux81),
	.datad(idex_sRST1),
	.cin(gnd),
	.combout(\rdat1_l~24_combout ),
	.cout());
// synopsys translate_off
defparam \rdat1_l~24 .lut_mask = 16'h00B8;
defparam \rdat1_l~24 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X68_Y36_N14
cycloneive_lcell_comb \rdat1_l~25 (
// Equation(s):
// \rdat1_l~25_combout  = (!idex_sRST1 & ((Selector1 & ((Mux9))) # (!Selector1 & (Mux91))))

	.dataa(idex_sRST1),
	.datab(Selector1),
	.datac(Mux91),
	.datad(Mux9),
	.cin(gnd),
	.combout(\rdat1_l~25_combout ),
	.cout());
// synopsys translate_off
defparam \rdat1_l~25 .lut_mask = 16'h5410;
defparam \rdat1_l~25 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y38_N18
cycloneive_lcell_comb \rdat1_l~26 (
// Equation(s):
// \rdat1_l~26_combout  = (!idex_sRST1 & ((Selector1 & (Mux10)) # (!Selector1 & ((Mux101)))))

	.dataa(idex_sRST1),
	.datab(Selector1),
	.datac(Mux10),
	.datad(Mux101),
	.cin(gnd),
	.combout(\rdat1_l~26_combout ),
	.cout());
// synopsys translate_off
defparam \rdat1_l~26 .lut_mask = 16'h5140;
defparam \rdat1_l~26 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y40_N30
cycloneive_lcell_comb \rdat1_l~27 (
// Equation(s):
// \rdat1_l~27_combout  = (!idex_sRST1 & ((Selector1 & ((Mux111))) # (!Selector1 & (Mux112))))

	.dataa(Selector1),
	.datab(idex_sRST1),
	.datac(Mux112),
	.datad(Mux111),
	.cin(gnd),
	.combout(\rdat1_l~27_combout ),
	.cout());
// synopsys translate_off
defparam \rdat1_l~27 .lut_mask = 16'h3210;
defparam \rdat1_l~27 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X67_Y36_N12
cycloneive_lcell_comb \rdat1_l~28 (
// Equation(s):
// \rdat1_l~28_combout  = (!idex_sRST1 & ((Selector1 & ((Mux12))) # (!Selector1 & (Mux121))))

	.dataa(Selector1),
	.datab(idex_sRST1),
	.datac(Mux121),
	.datad(Mux12),
	.cin(gnd),
	.combout(\rdat1_l~28_combout ),
	.cout());
// synopsys translate_off
defparam \rdat1_l~28 .lut_mask = 16'h3210;
defparam \rdat1_l~28 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X63_Y36_N10
cycloneive_lcell_comb \rdat1_l~29 (
// Equation(s):
// \rdat1_l~29_combout  = (!idex_sRST1 & ((Selector1 & ((Mux13))) # (!Selector1 & (Mux131))))

	.dataa(idex_sRST1),
	.datab(Mux131),
	.datac(Selector1),
	.datad(Mux13),
	.cin(gnd),
	.combout(\rdat1_l~29_combout ),
	.cout());
// synopsys translate_off
defparam \rdat1_l~29 .lut_mask = 16'h5404;
defparam \rdat1_l~29 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y40_N16
cycloneive_lcell_comb \rdat1_l~30 (
// Equation(s):
// \rdat1_l~30_combout  = (!idex_sRST1 & ((Selector1 & ((Mux14))) # (!Selector1 & (Mux141))))

	.dataa(Selector1),
	.datab(idex_sRST1),
	.datac(Mux141),
	.datad(Mux14),
	.cin(gnd),
	.combout(\rdat1_l~30_combout ),
	.cout());
// synopsys translate_off
defparam \rdat1_l~30 .lut_mask = 16'h3210;
defparam \rdat1_l~30 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y40_N16
cycloneive_lcell_comb \rdat1_l~31 (
// Equation(s):
// \rdat1_l~31_combout  = (!idex_sRST1 & ((Selector1 & ((Mux311))) # (!Selector1 & (Mux312))))

	.dataa(Mux312),
	.datab(Selector1),
	.datac(idex_sRST1),
	.datad(Mux311),
	.cin(gnd),
	.combout(\rdat1_l~31_combout ),
	.cout());
// synopsys translate_off
defparam \rdat1_l~31 .lut_mask = 16'h0E02;
defparam \rdat1_l~31 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y33_N22
cycloneive_lcell_comb \dmemREN_l~0 (
// Equation(s):
// \dmemREN_l~0_combout  = (!idex_sRST & (Equal21 & !idex_sRST2))

	.dataa(idex_sRST),
	.datab(Equal21),
	.datac(gnd),
	.datad(idex_sRST2),
	.cin(gnd),
	.combout(\dmemREN_l~0_combout ),
	.cout());
// synopsys translate_off
defparam \dmemREN_l~0 .lut_mask = 16'h0044;
defparam \dmemREN_l~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y32_N18
cycloneive_lcell_comb \wsel_l~1 (
// Equation(s):
// \wsel_l~1_combout  = (!Equal26 & ((\wsel_l~0_combout ) # ((Selector24 & plif_ifidinstr_l_16))))

	.dataa(\wsel_l~0_combout ),
	.datab(Equal26),
	.datac(Selector24),
	.datad(plif_ifidinstr_l_16),
	.cin(gnd),
	.combout(\wsel_l~1_combout ),
	.cout());
// synopsys translate_off
defparam \wsel_l~1 .lut_mask = 16'h3222;
defparam \wsel_l~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y32_N8
cycloneive_lcell_comb \wsel_l~2 (
// Equation(s):
// \wsel_l~2_combout  = (!idex_sRST1 & ((\wsel_l~1_combout ) # ((plif_ifidinstr_l_11 & Selector11))))

	.dataa(plif_ifidinstr_l_11),
	.datab(idex_sRST1),
	.datac(Selector11),
	.datad(\wsel_l~1_combout ),
	.cin(gnd),
	.combout(\wsel_l~2_combout ),
	.cout());
// synopsys translate_off
defparam \wsel_l~2 .lut_mask = 16'h3320;
defparam \wsel_l~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y29_N12
cycloneive_lcell_comb \wsel_l~0 (
// Equation(s):
// \wsel_l~0_combout  = (!plif_ifidinstr_l_31 & (!plif_ifidinstr_l_29 & (!plif_ifidinstr_l_30 & Equal16)))

	.dataa(plif_ifidinstr_l_31),
	.datab(plif_ifidinstr_l_29),
	.datac(plif_ifidinstr_l_30),
	.datad(Equal16),
	.cin(gnd),
	.combout(\wsel_l~0_combout ),
	.cout());
// synopsys translate_off
defparam \wsel_l~0 .lut_mask = 16'h0100;
defparam \wsel_l~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y31_N24
cycloneive_lcell_comb \wsel_l~3 (
// Equation(s):
// \wsel_l~3_combout  = (!Equal26 & ((\wsel_l~0_combout ) # ((plif_ifidinstr_l_17 & Selector24))))

	.dataa(plif_ifidinstr_l_17),
	.datab(Selector24),
	.datac(\wsel_l~0_combout ),
	.datad(Equal26),
	.cin(gnd),
	.combout(\wsel_l~3_combout ),
	.cout());
// synopsys translate_off
defparam \wsel_l~3 .lut_mask = 16'h00F8;
defparam \wsel_l~3 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y32_N22
cycloneive_lcell_comb \wsel_l~4 (
// Equation(s):
// \wsel_l~4_combout  = (!idex_sRST1 & ((\wsel_l~3_combout ) # ((Selector11 & plif_ifidinstr_l_12))))

	.dataa(\wsel_l~3_combout ),
	.datab(idex_sRST1),
	.datac(Selector11),
	.datad(plif_ifidinstr_l_12),
	.cin(gnd),
	.combout(\wsel_l~4_combout ),
	.cout());
// synopsys translate_off
defparam \wsel_l~4 .lut_mask = 16'h3222;
defparam \wsel_l~4 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y31_N6
cycloneive_lcell_comb \wsel_l~5 (
// Equation(s):
// \wsel_l~5_combout  = (!Equal26 & ((\wsel_l~0_combout ) # ((Selector24 & plif_ifidinstr_l_18))))

	.dataa(Equal26),
	.datab(Selector24),
	.datac(\wsel_l~0_combout ),
	.datad(plif_ifidinstr_l_18),
	.cin(gnd),
	.combout(\wsel_l~5_combout ),
	.cout());
// synopsys translate_off
defparam \wsel_l~5 .lut_mask = 16'h5450;
defparam \wsel_l~5 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y32_N26
cycloneive_lcell_comb \wsel_l~6 (
// Equation(s):
// \wsel_l~6_combout  = (!idex_sRST1 & ((\wsel_l~5_combout ) # ((plif_ifidinstr_l_13 & Selector11))))

	.dataa(plif_ifidinstr_l_13),
	.datab(idex_sRST1),
	.datac(Selector11),
	.datad(\wsel_l~5_combout ),
	.cin(gnd),
	.combout(\wsel_l~6_combout ),
	.cout());
// synopsys translate_off
defparam \wsel_l~6 .lut_mask = 16'h3320;
defparam \wsel_l~6 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y32_N20
cycloneive_lcell_comb \wsel_l~7 (
// Equation(s):
// \wsel_l~7_combout  = (!Equal26 & ((\wsel_l~0_combout ) # ((Selector24 & plif_ifidinstr_l_19))))

	.dataa(\wsel_l~0_combout ),
	.datab(Equal26),
	.datac(Selector24),
	.datad(plif_ifidinstr_l_19),
	.cin(gnd),
	.combout(\wsel_l~7_combout ),
	.cout());
// synopsys translate_off
defparam \wsel_l~7 .lut_mask = 16'h3222;
defparam \wsel_l~7 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y32_N24
cycloneive_lcell_comb \wsel_l~8 (
// Equation(s):
// \wsel_l~8_combout  = (!idex_sRST1 & ((\wsel_l~7_combout ) # ((plif_ifidinstr_l_14 & Selector11))))

	.dataa(plif_ifidinstr_l_14),
	.datab(idex_sRST1),
	.datac(Selector11),
	.datad(\wsel_l~7_combout ),
	.cin(gnd),
	.combout(\wsel_l~8_combout ),
	.cout());
// synopsys translate_off
defparam \wsel_l~8 .lut_mask = 16'h3320;
defparam \wsel_l~8 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y32_N2
cycloneive_lcell_comb \wsel_l~9 (
// Equation(s):
// \wsel_l~9_combout  = (!Equal26 & ((\wsel_l~0_combout ) # ((Selector24 & plif_ifidinstr_l_20))))

	.dataa(\wsel_l~0_combout ),
	.datab(Equal26),
	.datac(Selector24),
	.datad(plif_ifidinstr_l_20),
	.cin(gnd),
	.combout(\wsel_l~9_combout ),
	.cout());
// synopsys translate_off
defparam \wsel_l~9 .lut_mask = 16'h3222;
defparam \wsel_l~9 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y32_N4
cycloneive_lcell_comb \wsel_l~10 (
// Equation(s):
// \wsel_l~10_combout  = (!idex_sRST1 & ((\wsel_l~9_combout ) # ((plif_ifidinstr_l_15 & Selector11))))

	.dataa(plif_ifidinstr_l_15),
	.datab(idex_sRST1),
	.datac(Selector11),
	.datad(\wsel_l~9_combout ),
	.cin(gnd),
	.combout(\wsel_l~10_combout ),
	.cout());
// synopsys translate_off
defparam \wsel_l~10 .lut_mask = 16'h3320;
defparam \wsel_l~10 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y30_N26
cycloneive_lcell_comb \dmemWEN_l~0 (
// Equation(s):
// \dmemWEN_l~0_combout  = (!idex_sRST & (Equal22 & !idex_sRST2))

	.dataa(idex_sRST),
	.datab(gnd),
	.datac(Equal22),
	.datad(idex_sRST2),
	.cin(gnd),
	.combout(\dmemWEN_l~0_combout ),
	.cout());
// synopsys translate_off
defparam \dmemWEN_l~0 .lut_mask = 16'h0050;
defparam \dmemWEN_l~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y32_N0
cycloneive_lcell_comb \regen_l~0 (
// Equation(s):
// \regen_l~0_combout  = (!idex_sRST1 & ((Equal25) # ((Selector11) # (!WideOr161))))

	.dataa(Equal25),
	.datab(idex_sRST1),
	.datac(Selector11),
	.datad(WideOr16),
	.cin(gnd),
	.combout(\regen_l~0_combout ),
	.cout());
// synopsys translate_off
defparam \regen_l~0 .lut_mask = 16'h3233;
defparam \regen_l~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y32_N20
cycloneive_lcell_comb \regsrc_l~0 (
// Equation(s):
// \regsrc_l~0_combout  = (!idex_sRST2 & (!idex_sRST & ((Equal22) # (Equal21))))

	.dataa(Equal22),
	.datab(idex_sRST2),
	.datac(idex_sRST),
	.datad(Equal21),
	.cin(gnd),
	.combout(\regsrc_l~0_combout ),
	.cout());
// synopsys translate_off
defparam \regsrc_l~0 .lut_mask = 16'h0302;
defparam \regsrc_l~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y33_N20
cycloneive_lcell_comb \regsrc_l~1 (
// Equation(s):
// \regsrc_l~1_combout  = (!idex_sRST & (Equal25 & !idex_sRST2))

	.dataa(idex_sRST),
	.datab(gnd),
	.datac(Equal25),
	.datad(idex_sRST2),
	.cin(gnd),
	.combout(\regsrc_l~1_combout ),
	.cout());
// synopsys translate_off
defparam \regsrc_l~1 .lut_mask = 16'h0050;
defparam \regsrc_l~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y31_N26
cycloneive_lcell_comb \rtnaddr_l~0 (
// Equation(s):
// \rtnaddr_l~0_combout  = (!idex_sRST & (!idex_sRST2 & plif_ifidrtnaddr_l_31))

	.dataa(gnd),
	.datab(idex_sRST),
	.datac(idex_sRST2),
	.datad(plif_ifidrtnaddr_l_31),
	.cin(gnd),
	.combout(\rtnaddr_l~0_combout ),
	.cout());
// synopsys translate_off
defparam \rtnaddr_l~0 .lut_mask = 16'h0300;
defparam \rtnaddr_l~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y31_N16
cycloneive_lcell_comb \rtnaddr_l~1 (
// Equation(s):
// \rtnaddr_l~1_combout  = (!idex_sRST & (!idex_sRST2 & plif_ifidrtnaddr_l_30))

	.dataa(gnd),
	.datab(idex_sRST),
	.datac(idex_sRST2),
	.datad(plif_ifidrtnaddr_l_30),
	.cin(gnd),
	.combout(\rtnaddr_l~1_combout ),
	.cout());
// synopsys translate_off
defparam \rtnaddr_l~1 .lut_mask = 16'h0300;
defparam \rtnaddr_l~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y31_N14
cycloneive_lcell_comb \rtnaddr_l~2 (
// Equation(s):
// \rtnaddr_l~2_combout  = (!idex_sRST & (!idex_sRST2 & plif_ifidrtnaddr_l_29))

	.dataa(gnd),
	.datab(idex_sRST),
	.datac(idex_sRST2),
	.datad(plif_ifidrtnaddr_l_29),
	.cin(gnd),
	.combout(\rtnaddr_l~2_combout ),
	.cout());
// synopsys translate_off
defparam \rtnaddr_l~2 .lut_mask = 16'h0300;
defparam \rtnaddr_l~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y31_N10
cycloneive_lcell_comb \rtnaddr_l~3 (
// Equation(s):
// \rtnaddr_l~3_combout  = (!idex_sRST & (!idex_sRST2 & plif_ifidrtnaddr_l_28))

	.dataa(idex_sRST),
	.datab(gnd),
	.datac(idex_sRST2),
	.datad(plif_ifidrtnaddr_l_28),
	.cin(gnd),
	.combout(\rtnaddr_l~3_combout ),
	.cout());
// synopsys translate_off
defparam \rtnaddr_l~3 .lut_mask = 16'h0500;
defparam \rtnaddr_l~3 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X52_Y31_N12
cycloneive_lcell_comb \rtnaddr_l~4 (
// Equation(s):
// \rtnaddr_l~4_combout  = (!idex_sRST2 & (!idex_sRST & plif_ifidrtnaddr_l_27))

	.dataa(idex_sRST2),
	.datab(idex_sRST),
	.datac(plif_ifidrtnaddr_l_27),
	.datad(gnd),
	.cin(gnd),
	.combout(\rtnaddr_l~4_combout ),
	.cout());
// synopsys translate_off
defparam \rtnaddr_l~4 .lut_mask = 16'h1010;
defparam \rtnaddr_l~4 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X52_Y31_N10
cycloneive_lcell_comb \rtnaddr_l~5 (
// Equation(s):
// \rtnaddr_l~5_combout  = (!idex_sRST2 & (!idex_sRST & plif_ifidrtnaddr_l_26))

	.dataa(idex_sRST2),
	.datab(idex_sRST),
	.datac(plif_ifidrtnaddr_l_26),
	.datad(gnd),
	.cin(gnd),
	.combout(\rtnaddr_l~5_combout ),
	.cout());
// synopsys translate_off
defparam \rtnaddr_l~5 .lut_mask = 16'h1010;
defparam \rtnaddr_l~5 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X52_Y31_N20
cycloneive_lcell_comb \rtnaddr_l~6 (
// Equation(s):
// \rtnaddr_l~6_combout  = (!idex_sRST2 & (!idex_sRST & plif_ifidrtnaddr_l_25))

	.dataa(idex_sRST2),
	.datab(idex_sRST),
	.datac(plif_ifidrtnaddr_l_25),
	.datad(gnd),
	.cin(gnd),
	.combout(\rtnaddr_l~6_combout ),
	.cout());
// synopsys translate_off
defparam \rtnaddr_l~6 .lut_mask = 16'h1010;
defparam \rtnaddr_l~6 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X52_Y31_N2
cycloneive_lcell_comb \rtnaddr_l~7 (
// Equation(s):
// \rtnaddr_l~7_combout  = (!idex_sRST2 & (!idex_sRST & plif_ifidrtnaddr_l_24))

	.dataa(idex_sRST2),
	.datab(idex_sRST),
	.datac(plif_ifidrtnaddr_l_24),
	.datad(gnd),
	.cin(gnd),
	.combout(\rtnaddr_l~7_combout ),
	.cout());
// synopsys translate_off
defparam \rtnaddr_l~7 .lut_mask = 16'h1010;
defparam \rtnaddr_l~7 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X52_Y31_N24
cycloneive_lcell_comb \rtnaddr_l~8 (
// Equation(s):
// \rtnaddr_l~8_combout  = (!idex_sRST2 & (!idex_sRST & plif_ifidrtnaddr_l_23))

	.dataa(idex_sRST2),
	.datab(idex_sRST),
	.datac(plif_ifidrtnaddr_l_23),
	.datad(gnd),
	.cin(gnd),
	.combout(\rtnaddr_l~8_combout ),
	.cout());
// synopsys translate_off
defparam \rtnaddr_l~8 .lut_mask = 16'h1010;
defparam \rtnaddr_l~8 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X52_Y31_N6
cycloneive_lcell_comb \rtnaddr_l~9 (
// Equation(s):
// \rtnaddr_l~9_combout  = (!idex_sRST2 & (plif_ifidrtnaddr_l_22 & !idex_sRST))

	.dataa(idex_sRST2),
	.datab(plif_ifidrtnaddr_l_22),
	.datac(idex_sRST),
	.datad(gnd),
	.cin(gnd),
	.combout(\rtnaddr_l~9_combout ),
	.cout());
// synopsys translate_off
defparam \rtnaddr_l~9 .lut_mask = 16'h0404;
defparam \rtnaddr_l~9 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y30_N0
cycloneive_lcell_comb \rtnaddr_l~10 (
// Equation(s):
// \rtnaddr_l~10_combout  = (!idex_sRST2 & (!idex_sRST & plif_ifidrtnaddr_l_21))

	.dataa(idex_sRST2),
	.datab(gnd),
	.datac(idex_sRST),
	.datad(plif_ifidrtnaddr_l_21),
	.cin(gnd),
	.combout(\rtnaddr_l~10_combout ),
	.cout());
// synopsys translate_off
defparam \rtnaddr_l~10 .lut_mask = 16'h0500;
defparam \rtnaddr_l~10 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y30_N2
cycloneive_lcell_comb \rtnaddr_l~11 (
// Equation(s):
// \rtnaddr_l~11_combout  = (!idex_sRST2 & (!idex_sRST & plif_ifidrtnaddr_l_20))

	.dataa(idex_sRST2),
	.datab(gnd),
	.datac(idex_sRST),
	.datad(plif_ifidrtnaddr_l_20),
	.cin(gnd),
	.combout(\rtnaddr_l~11_combout ),
	.cout());
// synopsys translate_off
defparam \rtnaddr_l~11 .lut_mask = 16'h0500;
defparam \rtnaddr_l~11 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y30_N24
cycloneive_lcell_comb \rtnaddr_l~12 (
// Equation(s):
// \rtnaddr_l~12_combout  = (!idex_sRST2 & (!idex_sRST & plif_ifidrtnaddr_l_19))

	.dataa(idex_sRST2),
	.datab(gnd),
	.datac(idex_sRST),
	.datad(plif_ifidrtnaddr_l_19),
	.cin(gnd),
	.combout(\rtnaddr_l~12_combout ),
	.cout());
// synopsys translate_off
defparam \rtnaddr_l~12 .lut_mask = 16'h0500;
defparam \rtnaddr_l~12 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y30_N26
cycloneive_lcell_comb \rtnaddr_l~13 (
// Equation(s):
// \rtnaddr_l~13_combout  = (!idex_sRST2 & (!idex_sRST & plif_ifidrtnaddr_l_18))

	.dataa(idex_sRST2),
	.datab(gnd),
	.datac(idex_sRST),
	.datad(plif_ifidrtnaddr_l_18),
	.cin(gnd),
	.combout(\rtnaddr_l~13_combout ),
	.cout());
// synopsys translate_off
defparam \rtnaddr_l~13 .lut_mask = 16'h0500;
defparam \rtnaddr_l~13 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y30_N16
cycloneive_lcell_comb \rtnaddr_l~14 (
// Equation(s):
// \rtnaddr_l~14_combout  = (!idex_sRST2 & (!idex_sRST & plif_ifidrtnaddr_l_17))

	.dataa(idex_sRST2),
	.datab(idex_sRST),
	.datac(plif_ifidrtnaddr_l_17),
	.datad(gnd),
	.cin(gnd),
	.combout(\rtnaddr_l~14_combout ),
	.cout());
// synopsys translate_off
defparam \rtnaddr_l~14 .lut_mask = 16'h1010;
defparam \rtnaddr_l~14 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y30_N22
cycloneive_lcell_comb \rtnaddr_l~15 (
// Equation(s):
// \rtnaddr_l~15_combout  = (plif_ifidrtnaddr_l_16 & (!idex_sRST & !idex_sRST2))

	.dataa(plif_ifidrtnaddr_l_16),
	.datab(gnd),
	.datac(idex_sRST),
	.datad(idex_sRST2),
	.cin(gnd),
	.combout(\rtnaddr_l~15_combout ),
	.cout());
// synopsys translate_off
defparam \rtnaddr_l~15 .lut_mask = 16'h000A;
defparam \rtnaddr_l~15 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y30_N20
cycloneive_lcell_comb \rtnaddr_l~16 (
// Equation(s):
// \rtnaddr_l~16_combout  = (!idex_sRST2 & (!idex_sRST & plif_ifidrtnaddr_l_15))

	.dataa(idex_sRST2),
	.datab(gnd),
	.datac(idex_sRST),
	.datad(plif_ifidrtnaddr_l_15),
	.cin(gnd),
	.combout(\rtnaddr_l~16_combout ),
	.cout());
// synopsys translate_off
defparam \rtnaddr_l~16 .lut_mask = 16'h0500;
defparam \rtnaddr_l~16 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y30_N30
cycloneive_lcell_comb \rtnaddr_l~17 (
// Equation(s):
// \rtnaddr_l~17_combout  = (!idex_sRST2 & (!idex_sRST & plif_ifidrtnaddr_l_14))

	.dataa(idex_sRST2),
	.datab(gnd),
	.datac(idex_sRST),
	.datad(plif_ifidrtnaddr_l_14),
	.cin(gnd),
	.combout(\rtnaddr_l~17_combout ),
	.cout());
// synopsys translate_off
defparam \rtnaddr_l~17 .lut_mask = 16'h0500;
defparam \rtnaddr_l~17 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y31_N20
cycloneive_lcell_comb \rtnaddr_l~18 (
// Equation(s):
// \rtnaddr_l~18_combout  = (!idex_sRST & (!idex_sRST2 & plif_ifidrtnaddr_l_13))

	.dataa(idex_sRST),
	.datab(gnd),
	.datac(idex_sRST2),
	.datad(plif_ifidrtnaddr_l_13),
	.cin(gnd),
	.combout(\rtnaddr_l~18_combout ),
	.cout());
// synopsys translate_off
defparam \rtnaddr_l~18 .lut_mask = 16'h0500;
defparam \rtnaddr_l~18 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y31_N14
cycloneive_lcell_comb \rtnaddr_l~19 (
// Equation(s):
// \rtnaddr_l~19_combout  = (!idex_sRST & (!idex_sRST2 & plif_ifidrtnaddr_l_12))

	.dataa(idex_sRST),
	.datab(gnd),
	.datac(idex_sRST2),
	.datad(plif_ifidrtnaddr_l_12),
	.cin(gnd),
	.combout(\rtnaddr_l~19_combout ),
	.cout());
// synopsys translate_off
defparam \rtnaddr_l~19 .lut_mask = 16'h0500;
defparam \rtnaddr_l~19 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y31_N28
cycloneive_lcell_comb \rtnaddr_l~20 (
// Equation(s):
// \rtnaddr_l~20_combout  = (!idex_sRST & (!idex_sRST2 & plif_ifidrtnaddr_l_11))

	.dataa(idex_sRST),
	.datab(gnd),
	.datac(idex_sRST2),
	.datad(plif_ifidrtnaddr_l_11),
	.cin(gnd),
	.combout(\rtnaddr_l~20_combout ),
	.cout());
// synopsys translate_off
defparam \rtnaddr_l~20 .lut_mask = 16'h0500;
defparam \rtnaddr_l~20 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y31_N30
cycloneive_lcell_comb \rtnaddr_l~21 (
// Equation(s):
// \rtnaddr_l~21_combout  = (!idex_sRST & (!idex_sRST2 & plif_ifidrtnaddr_l_10))

	.dataa(idex_sRST),
	.datab(gnd),
	.datac(idex_sRST2),
	.datad(plif_ifidrtnaddr_l_10),
	.cin(gnd),
	.combout(\rtnaddr_l~21_combout ),
	.cout());
// synopsys translate_off
defparam \rtnaddr_l~21 .lut_mask = 16'h0500;
defparam \rtnaddr_l~21 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y31_N24
cycloneive_lcell_comb \rtnaddr_l~22 (
// Equation(s):
// \rtnaddr_l~22_combout  = (!idex_sRST & (plif_ifidrtnaddr_l_9 & !idex_sRST2))

	.dataa(idex_sRST),
	.datab(plif_ifidrtnaddr_l_9),
	.datac(idex_sRST2),
	.datad(gnd),
	.cin(gnd),
	.combout(\rtnaddr_l~22_combout ),
	.cout());
// synopsys translate_off
defparam \rtnaddr_l~22 .lut_mask = 16'h0404;
defparam \rtnaddr_l~22 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y31_N2
cycloneive_lcell_comb \rtnaddr_l~23 (
// Equation(s):
// \rtnaddr_l~23_combout  = (!idex_sRST & (!idex_sRST2 & plif_ifidrtnaddr_l_8))

	.dataa(idex_sRST),
	.datab(gnd),
	.datac(idex_sRST2),
	.datad(plif_ifidrtnaddr_l_8),
	.cin(gnd),
	.combout(\rtnaddr_l~23_combout ),
	.cout());
// synopsys translate_off
defparam \rtnaddr_l~23 .lut_mask = 16'h0500;
defparam \rtnaddr_l~23 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y31_N0
cycloneive_lcell_comb \rtnaddr_l~24 (
// Equation(s):
// \rtnaddr_l~24_combout  = (!idex_sRST & (!idex_sRST2 & plif_ifidrtnaddr_l_7))

	.dataa(idex_sRST),
	.datab(gnd),
	.datac(idex_sRST2),
	.datad(plif_ifidrtnaddr_l_7),
	.cin(gnd),
	.combout(\rtnaddr_l~24_combout ),
	.cout());
// synopsys translate_off
defparam \rtnaddr_l~24 .lut_mask = 16'h0500;
defparam \rtnaddr_l~24 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y31_N20
cycloneive_lcell_comb \rtnaddr_l~25 (
// Equation(s):
// \rtnaddr_l~25_combout  = (!idex_sRST & (!idex_sRST2 & plif_ifidrtnaddr_l_6))

	.dataa(gnd),
	.datab(idex_sRST),
	.datac(idex_sRST2),
	.datad(plif_ifidrtnaddr_l_6),
	.cin(gnd),
	.combout(\rtnaddr_l~25_combout ),
	.cout());
// synopsys translate_off
defparam \rtnaddr_l~25 .lut_mask = 16'h0300;
defparam \rtnaddr_l~25 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y31_N6
cycloneive_lcell_comb \rtnaddr_l~26 (
// Equation(s):
// \rtnaddr_l~26_combout  = (!idex_sRST & (!idex_sRST2 & plif_ifidrtnaddr_l_5))

	.dataa(idex_sRST),
	.datab(gnd),
	.datac(idex_sRST2),
	.datad(plif_ifidrtnaddr_l_5),
	.cin(gnd),
	.combout(\rtnaddr_l~26_combout ),
	.cout());
// synopsys translate_off
defparam \rtnaddr_l~26 .lut_mask = 16'h0500;
defparam \rtnaddr_l~26 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X50_Y41_N0
cycloneive_lcell_comb \rtnaddr_l~27 (
// Equation(s):
// \rtnaddr_l~27_combout  = (plif_ifidrtnaddr_l_2 & (!idex_sRST2 & !idex_sRST))

	.dataa(plif_ifidrtnaddr_l_2),
	.datab(idex_sRST2),
	.datac(gnd),
	.datad(idex_sRST),
	.cin(gnd),
	.combout(\rtnaddr_l~27_combout ),
	.cout());
// synopsys translate_off
defparam \rtnaddr_l~27 .lut_mask = 16'h0022;
defparam \rtnaddr_l~27 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X52_Y31_N16
cycloneive_lcell_comb \rtnaddr_l~28 (
// Equation(s):
// \rtnaddr_l~28_combout  = (!idex_sRST2 & (plif_ifidrtnaddr_l_1 & !idex_sRST))

	.dataa(idex_sRST2),
	.datab(plif_ifidrtnaddr_l_1),
	.datac(idex_sRST),
	.datad(gnd),
	.cin(gnd),
	.combout(\rtnaddr_l~28_combout ),
	.cout());
// synopsys translate_off
defparam \rtnaddr_l~28 .lut_mask = 16'h0404;
defparam \rtnaddr_l~28 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X50_Y41_N22
cycloneive_lcell_comb \rtnaddr_l~29 (
// Equation(s):
// \rtnaddr_l~29_combout  = (!idex_sRST2 & (plif_ifidrtnaddr_l_0 & !idex_sRST))

	.dataa(gnd),
	.datab(idex_sRST2),
	.datac(plif_ifidrtnaddr_l_0),
	.datad(idex_sRST),
	.cin(gnd),
	.combout(\rtnaddr_l~29_combout ),
	.cout());
// synopsys translate_off
defparam \rtnaddr_l~29 .lut_mask = 16'h0030;
defparam \rtnaddr_l~29 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X50_Y41_N28
cycloneive_lcell_comb \rtnaddr_l~30 (
// Equation(s):
// \rtnaddr_l~30_combout  = (plif_ifidrtnaddr_l_4 & (!idex_sRST2 & !idex_sRST))

	.dataa(plif_ifidrtnaddr_l_4),
	.datab(idex_sRST2),
	.datac(gnd),
	.datad(idex_sRST),
	.cin(gnd),
	.combout(\rtnaddr_l~30_combout ),
	.cout());
// synopsys translate_off
defparam \rtnaddr_l~30 .lut_mask = 16'h0022;
defparam \rtnaddr_l~30 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X50_Y41_N10
cycloneive_lcell_comb \rtnaddr_l~31 (
// Equation(s):
// \rtnaddr_l~31_combout  = (plif_ifidrtnaddr_l_3 & (!idex_sRST2 & !idex_sRST))

	.dataa(plif_ifidrtnaddr_l_3),
	.datab(idex_sRST2),
	.datac(gnd),
	.datad(idex_sRST),
	.cin(gnd),
	.combout(\rtnaddr_l~31_combout ),
	.cout());
// synopsys translate_off
defparam \rtnaddr_l~31 .lut_mask = 16'h0022;
defparam \rtnaddr_l~31 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y30_N12
cycloneive_lcell_comb \btype_l~0 (
// Equation(s):
// \btype_l~0_combout  = (!idex_sRST & (!idex_sRST2 & (Equal11 & Equal121)))

	.dataa(idex_sRST),
	.datab(idex_sRST2),
	.datac(Equal11),
	.datad(Equal121),
	.cin(gnd),
	.combout(\btype_l~0_combout ),
	.cout());
// synopsys translate_off
defparam \btype_l~0 .lut_mask = 16'h1000;
defparam \btype_l~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y30_N30
cycloneive_lcell_comb \jaddr_l~0 (
// Equation(s):
// \jaddr_l~0_combout  = (!pcsrc & (!idex_sRST & (plif_ifidinstr_l_1 & !idex_sRST2)))

	.dataa(pcsrc),
	.datab(idex_sRST),
	.datac(plif_ifidinstr_l_1),
	.datad(idex_sRST2),
	.cin(gnd),
	.combout(\jaddr_l~0_combout ),
	.cout());
// synopsys translate_off
defparam \jaddr_l~0 .lut_mask = 16'h0010;
defparam \jaddr_l~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y33_N26
cycloneive_lcell_comb \jaddr_l~1 (
// Equation(s):
// \jaddr_l~1_combout  = (!idex_sRST & (plif_ifidinstr_l_0 & (!pcsrc & !idex_sRST2)))

	.dataa(idex_sRST),
	.datab(plif_ifidinstr_l_0),
	.datac(pcsrc),
	.datad(idex_sRST2),
	.cin(gnd),
	.combout(\jaddr_l~1_combout ),
	.cout());
// synopsys translate_off
defparam \jaddr_l~1 .lut_mask = 16'h0004;
defparam \jaddr_l~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y33_N0
cycloneive_lcell_comb \jaddr_l~2 (
// Equation(s):
// \jaddr_l~2_combout  = (!idex_sRST & (plif_ifidinstr_l_3 & (!pcsrc & !idex_sRST2)))

	.dataa(idex_sRST),
	.datab(plif_ifidinstr_l_3),
	.datac(pcsrc),
	.datad(idex_sRST2),
	.cin(gnd),
	.combout(\jaddr_l~2_combout ),
	.cout());
// synopsys translate_off
defparam \jaddr_l~2 .lut_mask = 16'h0004;
defparam \jaddr_l~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y33_N14
cycloneive_lcell_comb \jaddr_l~3 (
// Equation(s):
// \jaddr_l~3_combout  = (!idex_sRST & (plif_ifidinstr_l_2 & (!pcsrc & !idex_sRST2)))

	.dataa(idex_sRST),
	.datab(plif_ifidinstr_l_2),
	.datac(pcsrc),
	.datad(idex_sRST2),
	.cin(gnd),
	.combout(\jaddr_l~3_combout ),
	.cout());
// synopsys translate_off
defparam \jaddr_l~3 .lut_mask = 16'h0004;
defparam \jaddr_l~3 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y30_N12
cycloneive_lcell_comb \jaddr_l~4 (
// Equation(s):
// \jaddr_l~4_combout  = (!pcsrc & (!idex_sRST & (plif_ifidinstr_l_5 & !idex_sRST2)))

	.dataa(pcsrc),
	.datab(idex_sRST),
	.datac(plif_ifidinstr_l_5),
	.datad(idex_sRST2),
	.cin(gnd),
	.combout(\jaddr_l~4_combout ),
	.cout());
// synopsys translate_off
defparam \jaddr_l~4 .lut_mask = 16'h0010;
defparam \jaddr_l~4 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y33_N12
cycloneive_lcell_comb \jaddr_l~5 (
// Equation(s):
// \jaddr_l~5_combout  = (!idex_sRST & (plif_ifidinstr_l_4 & (!pcsrc & !idex_sRST2)))

	.dataa(idex_sRST),
	.datab(plif_ifidinstr_l_4),
	.datac(pcsrc),
	.datad(idex_sRST2),
	.cin(gnd),
	.combout(\jaddr_l~5_combout ),
	.cout());
// synopsys translate_off
defparam \jaddr_l~5 .lut_mask = 16'h0004;
defparam \jaddr_l~5 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y32_N14
cycloneive_lcell_comb \jaddr_l~6 (
// Equation(s):
// \jaddr_l~6_combout  = (plif_ifidinstr_l_7 & (!idex_sRST2 & (!idex_sRST & !pcsrc)))

	.dataa(plif_ifidinstr_l_7),
	.datab(idex_sRST2),
	.datac(idex_sRST),
	.datad(pcsrc),
	.cin(gnd),
	.combout(\jaddr_l~6_combout ),
	.cout());
// synopsys translate_off
defparam \jaddr_l~6 .lut_mask = 16'h0002;
defparam \jaddr_l~6 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y33_N30
cycloneive_lcell_comb \jaddr_l~7 (
// Equation(s):
// \jaddr_l~7_combout  = (!idex_sRST & (plif_ifidinstr_l_6 & (!pcsrc & !idex_sRST2)))

	.dataa(idex_sRST),
	.datab(plif_ifidinstr_l_6),
	.datac(pcsrc),
	.datad(idex_sRST2),
	.cin(gnd),
	.combout(\jaddr_l~7_combout ),
	.cout());
// synopsys translate_off
defparam \jaddr_l~7 .lut_mask = 16'h0004;
defparam \jaddr_l~7 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y33_N24
cycloneive_lcell_comb \jaddr_l~8 (
// Equation(s):
// \jaddr_l~8_combout  = (!idex_sRST & (plif_ifidinstr_l_9 & (!pcsrc & !idex_sRST2)))

	.dataa(idex_sRST),
	.datab(plif_ifidinstr_l_9),
	.datac(pcsrc),
	.datad(idex_sRST2),
	.cin(gnd),
	.combout(\jaddr_l~8_combout ),
	.cout());
// synopsys translate_off
defparam \jaddr_l~8 .lut_mask = 16'h0004;
defparam \jaddr_l~8 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y33_N6
cycloneive_lcell_comb \jaddr_l~9 (
// Equation(s):
// \jaddr_l~9_combout  = (!idex_sRST & (plif_ifidinstr_l_8 & (!pcsrc & !idex_sRST2)))

	.dataa(idex_sRST),
	.datab(plif_ifidinstr_l_8),
	.datac(pcsrc),
	.datad(idex_sRST2),
	.cin(gnd),
	.combout(\jaddr_l~9_combout ),
	.cout());
// synopsys translate_off
defparam \jaddr_l~9 .lut_mask = 16'h0004;
defparam \jaddr_l~9 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y33_N4
cycloneive_lcell_comb \jaddr_l~10 (
// Equation(s):
// \jaddr_l~10_combout  = (!idex_sRST & (plif_ifidinstr_l_11 & (!pcsrc & !idex_sRST2)))

	.dataa(idex_sRST),
	.datab(plif_ifidinstr_l_11),
	.datac(pcsrc),
	.datad(idex_sRST2),
	.cin(gnd),
	.combout(\jaddr_l~10_combout ),
	.cout());
// synopsys translate_off
defparam \jaddr_l~10 .lut_mask = 16'h0004;
defparam \jaddr_l~10 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y33_N2
cycloneive_lcell_comb \jaddr_l~11 (
// Equation(s):
// \jaddr_l~11_combout  = (!idex_sRST & (plif_ifidinstr_l_10 & (!pcsrc & !idex_sRST2)))

	.dataa(idex_sRST),
	.datab(plif_ifidinstr_l_10),
	.datac(pcsrc),
	.datad(idex_sRST2),
	.cin(gnd),
	.combout(\jaddr_l~11_combout ),
	.cout());
// synopsys translate_off
defparam \jaddr_l~11 .lut_mask = 16'h0004;
defparam \jaddr_l~11 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y32_N28
cycloneive_lcell_comb \jaddr_l~12 (
// Equation(s):
// \jaddr_l~12_combout  = (plif_ifidinstr_l_13 & (!idex_sRST & (!idex_sRST2 & !pcsrc)))

	.dataa(plif_ifidinstr_l_13),
	.datab(idex_sRST),
	.datac(idex_sRST2),
	.datad(pcsrc),
	.cin(gnd),
	.combout(\jaddr_l~12_combout ),
	.cout());
// synopsys translate_off
defparam \jaddr_l~12 .lut_mask = 16'h0002;
defparam \jaddr_l~12 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y31_N2
cycloneive_lcell_comb \jaddr_l~13 (
// Equation(s):
// \jaddr_l~13_combout  = (!idex_sRST2 & (!idex_sRST & (plif_ifidinstr_l_12 & !pcsrc)))

	.dataa(idex_sRST2),
	.datab(idex_sRST),
	.datac(plif_ifidinstr_l_12),
	.datad(pcsrc),
	.cin(gnd),
	.combout(\jaddr_l~13_combout ),
	.cout());
// synopsys translate_off
defparam \jaddr_l~13 .lut_mask = 16'h0010;
defparam \jaddr_l~13 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y31_N24
cycloneive_lcell_comb \jaddr_l~14 (
// Equation(s):
// \jaddr_l~14_combout  = (!idex_sRST2 & (!idex_sRST & (plif_ifidinstr_l_15 & !pcsrc)))

	.dataa(idex_sRST2),
	.datab(idex_sRST),
	.datac(plif_ifidinstr_l_15),
	.datad(pcsrc),
	.cin(gnd),
	.combout(\jaddr_l~14_combout ),
	.cout());
// synopsys translate_off
defparam \jaddr_l~14 .lut_mask = 16'h0010;
defparam \jaddr_l~14 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y30_N26
cycloneive_lcell_comb \jaddr_l~15 (
// Equation(s):
// \jaddr_l~15_combout  = (plif_ifidinstr_l_14 & (!pcsrc & (!idex_sRST & !idex_sRST2)))

	.dataa(plif_ifidinstr_l_14),
	.datab(pcsrc),
	.datac(idex_sRST),
	.datad(idex_sRST2),
	.cin(gnd),
	.combout(\jaddr_l~15_combout ),
	.cout());
// synopsys translate_off
defparam \jaddr_l~15 .lut_mask = 16'h0002;
defparam \jaddr_l~15 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y31_N18
cycloneive_lcell_comb \jaddr_l~16 (
// Equation(s):
// \jaddr_l~16_combout  = (plif_ifidinstr_l_17 & (!idex_sRST & (!idex_sRST2 & !pcsrc)))

	.dataa(plif_ifidinstr_l_17),
	.datab(idex_sRST),
	.datac(idex_sRST2),
	.datad(pcsrc),
	.cin(gnd),
	.combout(\jaddr_l~16_combout ),
	.cout());
// synopsys translate_off
defparam \jaddr_l~16 .lut_mask = 16'h0002;
defparam \jaddr_l~16 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y33_N16
cycloneive_lcell_comb \jaddr_l~17 (
// Equation(s):
// \jaddr_l~17_combout  = (!idex_sRST & (plif_ifidinstr_l_16 & (!pcsrc & !idex_sRST2)))

	.dataa(idex_sRST),
	.datab(plif_ifidinstr_l_16),
	.datac(pcsrc),
	.datad(idex_sRST2),
	.cin(gnd),
	.combout(\jaddr_l~17_combout ),
	.cout());
// synopsys translate_off
defparam \jaddr_l~17 .lut_mask = 16'h0004;
defparam \jaddr_l~17 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y37_N10
cycloneive_lcell_comb \jaddr_l~18 (
// Equation(s):
// \jaddr_l~18_combout  = (!pcsrc & (!idex_sRST2 & (!idex_sRST & plif_ifidinstr_l_19)))

	.dataa(pcsrc),
	.datab(idex_sRST2),
	.datac(idex_sRST),
	.datad(plif_ifidinstr_l_19),
	.cin(gnd),
	.combout(\jaddr_l~18_combout ),
	.cout());
// synopsys translate_off
defparam \jaddr_l~18 .lut_mask = 16'h0100;
defparam \jaddr_l~18 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y37_N8
cycloneive_lcell_comb \jaddr_l~19 (
// Equation(s):
// \jaddr_l~19_combout  = (!pcsrc & (!idex_sRST2 & (!idex_sRST & plif_ifidinstr_l_18)))

	.dataa(pcsrc),
	.datab(idex_sRST2),
	.datac(idex_sRST),
	.datad(plif_ifidinstr_l_18),
	.cin(gnd),
	.combout(\jaddr_l~19_combout ),
	.cout());
// synopsys translate_off
defparam \jaddr_l~19 .lut_mask = 16'h0100;
defparam \jaddr_l~19 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y37_N14
cycloneive_lcell_comb \jaddr_l~20 (
// Equation(s):
// \jaddr_l~20_combout  = (!idex_sRST2 & (!pcsrc & (!idex_sRST & plif_ifidinstr_l_21)))

	.dataa(idex_sRST2),
	.datab(pcsrc),
	.datac(idex_sRST),
	.datad(plif_ifidinstr_l_21),
	.cin(gnd),
	.combout(\jaddr_l~20_combout ),
	.cout());
// synopsys translate_off
defparam \jaddr_l~20 .lut_mask = 16'h0100;
defparam \jaddr_l~20 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y37_N18
cycloneive_lcell_comb \jaddr_l~21 (
// Equation(s):
// \jaddr_l~21_combout  = (!pcsrc & (!idex_sRST2 & (!idex_sRST & plif_ifidinstr_l_20)))

	.dataa(pcsrc),
	.datab(idex_sRST2),
	.datac(idex_sRST),
	.datad(plif_ifidinstr_l_20),
	.cin(gnd),
	.combout(\jaddr_l~21_combout ),
	.cout());
// synopsys translate_off
defparam \jaddr_l~21 .lut_mask = 16'h0100;
defparam \jaddr_l~21 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y37_N24
cycloneive_lcell_comb \jaddr_l~22 (
// Equation(s):
// \jaddr_l~22_combout  = (!pcsrc & (plif_ifidinstr_l_23 & (!idex_sRST & !idex_sRST2)))

	.dataa(pcsrc),
	.datab(plif_ifidinstr_l_23),
	.datac(idex_sRST),
	.datad(idex_sRST2),
	.cin(gnd),
	.combout(\jaddr_l~22_combout ),
	.cout());
// synopsys translate_off
defparam \jaddr_l~22 .lut_mask = 16'h0004;
defparam \jaddr_l~22 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y33_N10
cycloneive_lcell_comb \jaddr_l~23 (
// Equation(s):
// \jaddr_l~23_combout  = (!idex_sRST & (plif_ifidinstr_l_22 & (!pcsrc & !idex_sRST2)))

	.dataa(idex_sRST),
	.datab(plif_ifidinstr_l_22),
	.datac(pcsrc),
	.datad(idex_sRST2),
	.cin(gnd),
	.combout(\jaddr_l~23_combout ),
	.cout());
// synopsys translate_off
defparam \jaddr_l~23 .lut_mask = 16'h0004;
defparam \jaddr_l~23 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y37_N14
cycloneive_lcell_comb \jaddr_l~24 (
// Equation(s):
// \jaddr_l~24_combout  = (!pcsrc & (!idex_sRST2 & (!idex_sRST & plif_ifidinstr_l_25)))

	.dataa(pcsrc),
	.datab(idex_sRST2),
	.datac(idex_sRST),
	.datad(plif_ifidinstr_l_25),
	.cin(gnd),
	.combout(\jaddr_l~24_combout ),
	.cout());
// synopsys translate_off
defparam \jaddr_l~24 .lut_mask = 16'h0100;
defparam \jaddr_l~24 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y37_N28
cycloneive_lcell_comb \jaddr_l~25 (
// Equation(s):
// \jaddr_l~25_combout  = (!pcsrc & (!idex_sRST2 & (!idex_sRST & plif_ifidinstr_l_24)))

	.dataa(pcsrc),
	.datab(idex_sRST2),
	.datac(idex_sRST),
	.datad(plif_ifidinstr_l_24),
	.cin(gnd),
	.combout(\jaddr_l~25_combout ),
	.cout());
// synopsys translate_off
defparam \jaddr_l~25 .lut_mask = 16'h0100;
defparam \jaddr_l~25 .sum_lutc_input = "datac";
// synopsys translate_on

endmodule

module pipeline_ifid (
	PCreg_1,
	PCreg_0,
	pcifrtnaddr_2,
	pcifrtnaddr_3,
	pcifrtnaddr_4,
	pcifrtnaddr_5,
	pcifrtnaddr_6,
	pcifrtnaddr_7,
	pcifrtnaddr_8,
	pcifrtnaddr_9,
	pcifrtnaddr_10,
	pcifrtnaddr_11,
	pcifrtnaddr_12,
	pcifrtnaddr_13,
	pcifrtnaddr_14,
	pcifrtnaddr_15,
	pcifrtnaddr_16,
	pcifrtnaddr_17,
	pcifrtnaddr_18,
	pcifrtnaddr_19,
	pcifrtnaddr_20,
	pcifrtnaddr_21,
	pcifrtnaddr_22,
	pcifrtnaddr_23,
	pcifrtnaddr_24,
	pcifrtnaddr_25,
	pcifrtnaddr_26,
	pcifrtnaddr_27,
	pcifrtnaddr_28,
	pcifrtnaddr_29,
	pcifrtnaddr_30,
	pcifrtnaddr_31,
	ramiframload_0,
	ramiframload_1,
	ramiframload_2,
	ramiframload_3,
	ramiframload_4,
	ramiframload_5,
	ramiframload_6,
	ramiframload_7,
	ramiframload_8,
	ramiframload_9,
	ramiframload_10,
	ramiframload_11,
	ramiframload_12,
	ramiframload_13,
	ramiframload_14,
	ramiframload_15,
	ramiframload_16,
	ramiframload_17,
	ramiframload_18,
	ramiframload_19,
	ramiframload_20,
	ramiframload_21,
	ramiframload_22,
	ramiframload_23,
	ramiframload_24,
	ramiframload_25,
	ramiframload_26,
	ramiframload_27,
	ramiframload_28,
	ramiframload_29,
	ramiframload_30,
	ramiframload_31,
	plif_ifidinstr_l_31,
	plif_ifidinstr_l_29,
	plif_ifidinstr_l_27,
	plif_ifidinstr_l_26,
	plif_ifidinstr_l_28,
	plif_ifidinstr_l_30,
	plif_ifidinstr_l_5,
	plif_ifidinstr_l_1,
	plif_ifidinstr_l_0,
	plif_ifidinstr_l_2,
	plif_ifidinstr_l_3,
	plif_ifidinstr_l_4,
	plif_ifidinstr_l_22,
	plif_ifidinstr_l_21,
	plif_ifidinstr_l_24,
	plif_ifidinstr_l_23,
	plif_ifidinstr_l_25,
	plif_ifidinstr_l_17,
	plif_ifidinstr_l_16,
	plif_ifidinstr_l_19,
	plif_ifidinstr_l_18,
	plif_ifidinstr_l_20,
	ifid_en,
	plif_ifidinstr_l_15,
	plif_ifidinstr_l_14,
	plif_ifidinstr_l_13,
	plif_ifidinstr_l_12,
	plif_ifidinstr_l_11,
	plif_ifidinstr_l_10,
	plif_ifidinstr_l_9,
	plif_ifidinstr_l_8,
	plif_ifidinstr_l_7,
	plif_ifidinstr_l_6,
	instr_31,
	instr_29,
	instr_27,
	instr_26,
	instr_28,
	instr_30,
	instr_5,
	instr_1,
	instr_0,
	instr_2,
	instr_3,
	instr_4,
	instr_22,
	instr_21,
	instr_24,
	instr_23,
	instr_25,
	instr_17,
	instr_16,
	instr_19,
	instr_18,
	instr_20,
	instr_15,
	instr_14,
	instr_13,
	instr_12,
	instr_11,
	instr_10,
	instr_9,
	instr_8,
	instr_7,
	instr_6,
	plif_ifidrtnaddr_l_31,
	plif_ifidrtnaddr_l_30,
	plif_ifidrtnaddr_l_29,
	plif_ifidrtnaddr_l_28,
	plif_ifidrtnaddr_l_27,
	plif_ifidrtnaddr_l_26,
	plif_ifidrtnaddr_l_25,
	plif_ifidrtnaddr_l_24,
	plif_ifidrtnaddr_l_23,
	plif_ifidrtnaddr_l_22,
	plif_ifidrtnaddr_l_21,
	plif_ifidrtnaddr_l_20,
	plif_ifidrtnaddr_l_19,
	plif_ifidrtnaddr_l_18,
	plif_ifidrtnaddr_l_17,
	plif_ifidrtnaddr_l_16,
	plif_ifidrtnaddr_l_15,
	plif_ifidrtnaddr_l_14,
	plif_ifidrtnaddr_l_13,
	plif_ifidrtnaddr_l_12,
	plif_ifidrtnaddr_l_11,
	plif_ifidrtnaddr_l_10,
	plif_ifidrtnaddr_l_9,
	plif_ifidrtnaddr_l_8,
	plif_ifidrtnaddr_l_7,
	plif_ifidrtnaddr_l_6,
	plif_ifidrtnaddr_l_5,
	plif_ifidrtnaddr_l_2,
	plif_ifidrtnaddr_l_1,
	plif_ifidrtnaddr_l_0,
	plif_ifidrtnaddr_l_4,
	plif_ifidrtnaddr_l_3,
	ccifiwait_0,
	ifid_sRST,
	CPUCLK,
	nRST,
	devpor,
	devclrn,
	devoe);
input 	PCreg_1;
input 	PCreg_0;
input 	pcifrtnaddr_2;
input 	pcifrtnaddr_3;
input 	pcifrtnaddr_4;
input 	pcifrtnaddr_5;
input 	pcifrtnaddr_6;
input 	pcifrtnaddr_7;
input 	pcifrtnaddr_8;
input 	pcifrtnaddr_9;
input 	pcifrtnaddr_10;
input 	pcifrtnaddr_11;
input 	pcifrtnaddr_12;
input 	pcifrtnaddr_13;
input 	pcifrtnaddr_14;
input 	pcifrtnaddr_15;
input 	pcifrtnaddr_16;
input 	pcifrtnaddr_17;
input 	pcifrtnaddr_18;
input 	pcifrtnaddr_19;
input 	pcifrtnaddr_20;
input 	pcifrtnaddr_21;
input 	pcifrtnaddr_22;
input 	pcifrtnaddr_23;
input 	pcifrtnaddr_24;
input 	pcifrtnaddr_25;
input 	pcifrtnaddr_26;
input 	pcifrtnaddr_27;
input 	pcifrtnaddr_28;
input 	pcifrtnaddr_29;
input 	pcifrtnaddr_30;
input 	pcifrtnaddr_31;
input 	ramiframload_0;
input 	ramiframload_1;
input 	ramiframload_2;
input 	ramiframload_3;
input 	ramiframload_4;
input 	ramiframload_5;
input 	ramiframload_6;
input 	ramiframload_7;
input 	ramiframload_8;
input 	ramiframload_9;
input 	ramiframload_10;
input 	ramiframload_11;
input 	ramiframload_12;
input 	ramiframload_13;
input 	ramiframload_14;
input 	ramiframload_15;
input 	ramiframload_16;
input 	ramiframload_17;
input 	ramiframload_18;
input 	ramiframload_19;
input 	ramiframload_20;
input 	ramiframload_21;
input 	ramiframload_22;
input 	ramiframload_23;
input 	ramiframload_24;
input 	ramiframload_25;
input 	ramiframload_26;
input 	ramiframload_27;
input 	ramiframload_28;
input 	ramiframload_29;
input 	ramiframload_30;
input 	ramiframload_31;
output 	plif_ifidinstr_l_31;
output 	plif_ifidinstr_l_29;
output 	plif_ifidinstr_l_27;
output 	plif_ifidinstr_l_26;
output 	plif_ifidinstr_l_28;
output 	plif_ifidinstr_l_30;
output 	plif_ifidinstr_l_5;
output 	plif_ifidinstr_l_1;
output 	plif_ifidinstr_l_0;
output 	plif_ifidinstr_l_2;
output 	plif_ifidinstr_l_3;
output 	plif_ifidinstr_l_4;
output 	plif_ifidinstr_l_22;
output 	plif_ifidinstr_l_21;
output 	plif_ifidinstr_l_24;
output 	plif_ifidinstr_l_23;
output 	plif_ifidinstr_l_25;
output 	plif_ifidinstr_l_17;
output 	plif_ifidinstr_l_16;
output 	plif_ifidinstr_l_19;
output 	plif_ifidinstr_l_18;
output 	plif_ifidinstr_l_20;
input 	ifid_en;
output 	plif_ifidinstr_l_15;
output 	plif_ifidinstr_l_14;
output 	plif_ifidinstr_l_13;
output 	plif_ifidinstr_l_12;
output 	plif_ifidinstr_l_11;
output 	plif_ifidinstr_l_10;
output 	plif_ifidinstr_l_9;
output 	plif_ifidinstr_l_8;
output 	plif_ifidinstr_l_7;
output 	plif_ifidinstr_l_6;
input 	instr_31;
input 	instr_29;
input 	instr_27;
input 	instr_26;
input 	instr_28;
input 	instr_30;
input 	instr_5;
input 	instr_1;
input 	instr_0;
input 	instr_2;
input 	instr_3;
input 	instr_4;
input 	instr_22;
input 	instr_21;
input 	instr_24;
input 	instr_23;
input 	instr_25;
input 	instr_17;
input 	instr_16;
input 	instr_19;
input 	instr_18;
input 	instr_20;
input 	instr_15;
input 	instr_14;
input 	instr_13;
input 	instr_12;
input 	instr_11;
input 	instr_10;
input 	instr_9;
input 	instr_8;
input 	instr_7;
input 	instr_6;
output 	plif_ifidrtnaddr_l_31;
output 	plif_ifidrtnaddr_l_30;
output 	plif_ifidrtnaddr_l_29;
output 	plif_ifidrtnaddr_l_28;
output 	plif_ifidrtnaddr_l_27;
output 	plif_ifidrtnaddr_l_26;
output 	plif_ifidrtnaddr_l_25;
output 	plif_ifidrtnaddr_l_24;
output 	plif_ifidrtnaddr_l_23;
output 	plif_ifidrtnaddr_l_22;
output 	plif_ifidrtnaddr_l_21;
output 	plif_ifidrtnaddr_l_20;
output 	plif_ifidrtnaddr_l_19;
output 	plif_ifidrtnaddr_l_18;
output 	plif_ifidrtnaddr_l_17;
output 	plif_ifidrtnaddr_l_16;
output 	plif_ifidrtnaddr_l_15;
output 	plif_ifidrtnaddr_l_14;
output 	plif_ifidrtnaddr_l_13;
output 	plif_ifidrtnaddr_l_12;
output 	plif_ifidrtnaddr_l_11;
output 	plif_ifidrtnaddr_l_10;
output 	plif_ifidrtnaddr_l_9;
output 	plif_ifidrtnaddr_l_8;
output 	plif_ifidrtnaddr_l_7;
output 	plif_ifidrtnaddr_l_6;
output 	plif_ifidrtnaddr_l_5;
output 	plif_ifidrtnaddr_l_2;
output 	plif_ifidrtnaddr_l_1;
output 	plif_ifidrtnaddr_l_0;
output 	plif_ifidrtnaddr_l_4;
output 	plif_ifidrtnaddr_l_3;
input 	ccifiwait_0;
input 	ifid_sRST;
input 	CPUCLK;
input 	nRST;

// Design Ports Information

input 	devpor;
input 	devclrn;
input 	devoe;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
assign unknown = 1'bx;

wire \instr_l~0_combout ;
wire \plif_ifid.rtnaddr_l[24]~0_combout ;
wire \instr_l~1_combout ;
wire \instr_l~2_combout ;
wire \instr_l~3_combout ;
wire \instr_l~4_combout ;
wire \instr_l~5_combout ;
wire \instr_l~6_combout ;
wire \instr_l~7_combout ;
wire \instr_l~8_combout ;
wire \instr_l~9_combout ;
wire \instr_l~10_combout ;
wire \instr_l~11_combout ;
wire \instr_l~12_combout ;
wire \instr_l~13_combout ;
wire \instr_l~14_combout ;
wire \instr_l~15_combout ;
wire \instr_l~16_combout ;
wire \instr_l~17_combout ;
wire \instr_l~18_combout ;
wire \instr_l~19_combout ;
wire \instr_l~20_combout ;
wire \instr_l~21_combout ;
wire \instr_l~22_combout ;
wire \instr_l~23_combout ;
wire \instr_l~24_combout ;
wire \instr_l~25_combout ;
wire \instr_l~26_combout ;
wire \instr_l~27_combout ;
wire \instr_l~28_combout ;
wire \instr_l~29_combout ;
wire \instr_l~30_combout ;
wire \instr_l~31_combout ;
wire \rtnaddr_l~0_combout ;
wire \rtnaddr_l~1_combout ;
wire \rtnaddr_l~2_combout ;
wire \rtnaddr_l~3_combout ;
wire \rtnaddr_l~4_combout ;
wire \rtnaddr_l~5_combout ;
wire \rtnaddr_l~6_combout ;
wire \rtnaddr_l~7_combout ;
wire \rtnaddr_l~8_combout ;
wire \rtnaddr_l~9_combout ;
wire \rtnaddr_l~10_combout ;
wire \rtnaddr_l~11_combout ;
wire \rtnaddr_l~12_combout ;
wire \rtnaddr_l~13_combout ;
wire \rtnaddr_l~14_combout ;
wire \rtnaddr_l~15_combout ;
wire \rtnaddr_l~16_combout ;
wire \rtnaddr_l~17_combout ;
wire \rtnaddr_l~18_combout ;
wire \rtnaddr_l~19_combout ;
wire \rtnaddr_l~20_combout ;
wire \rtnaddr_l~21_combout ;
wire \rtnaddr_l~22_combout ;
wire \rtnaddr_l~23_combout ;
wire \rtnaddr_l~24_combout ;
wire \rtnaddr_l~25_combout ;
wire \rtnaddr_l~26_combout ;
wire \rtnaddr_l~27_combout ;
wire \rtnaddr_l~28_combout ;
wire \rtnaddr_l~29_combout ;
wire \rtnaddr_l~30_combout ;
wire \rtnaddr_l~31_combout ;


// Location: FF_X59_Y30_N11
dffeas \plif_ifid.instr_l[31] (
	.clk(CPUCLK),
	.d(\instr_l~0_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\plif_ifid.rtnaddr_l[24]~0_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(plif_ifidinstr_l_31),
	.prn(vcc));
// synopsys translate_off
defparam \plif_ifid.instr_l[31] .is_wysiwyg = "true";
defparam \plif_ifid.instr_l[31] .power_up = "low";
// synopsys translate_on

// Location: FF_X59_Y30_N9
dffeas \plif_ifid.instr_l[29] (
	.clk(CPUCLK),
	.d(\instr_l~1_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\plif_ifid.rtnaddr_l[24]~0_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(plif_ifidinstr_l_29),
	.prn(vcc));
// synopsys translate_off
defparam \plif_ifid.instr_l[29] .is_wysiwyg = "true";
defparam \plif_ifid.instr_l[29] .power_up = "low";
// synopsys translate_on

// Location: FF_X59_Y30_N7
dffeas \plif_ifid.instr_l[27] (
	.clk(CPUCLK),
	.d(\instr_l~2_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\plif_ifid.rtnaddr_l[24]~0_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(plif_ifidinstr_l_27),
	.prn(vcc));
// synopsys translate_off
defparam \plif_ifid.instr_l[27] .is_wysiwyg = "true";
defparam \plif_ifid.instr_l[27] .power_up = "low";
// synopsys translate_on

// Location: FF_X58_Y30_N25
dffeas \plif_ifid.instr_l[26] (
	.clk(CPUCLK),
	.d(\instr_l~3_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\plif_ifid.rtnaddr_l[24]~0_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(plif_ifidinstr_l_26),
	.prn(vcc));
// synopsys translate_off
defparam \plif_ifid.instr_l[26] .is_wysiwyg = "true";
defparam \plif_ifid.instr_l[26] .power_up = "low";
// synopsys translate_on

// Location: FF_X58_Y30_N7
dffeas \plif_ifid.instr_l[28] (
	.clk(CPUCLK),
	.d(\instr_l~4_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\plif_ifid.rtnaddr_l[24]~0_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(plif_ifidinstr_l_28),
	.prn(vcc));
// synopsys translate_off
defparam \plif_ifid.instr_l[28] .is_wysiwyg = "true";
defparam \plif_ifid.instr_l[28] .power_up = "low";
// synopsys translate_on

// Location: FF_X59_Y30_N31
dffeas \plif_ifid.instr_l[30] (
	.clk(CPUCLK),
	.d(\instr_l~5_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\plif_ifid.rtnaddr_l[24]~0_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(plif_ifidinstr_l_30),
	.prn(vcc));
// synopsys translate_off
defparam \plif_ifid.instr_l[30] .is_wysiwyg = "true";
defparam \plif_ifid.instr_l[30] .power_up = "low";
// synopsys translate_on

// Location: FF_X58_Y30_N29
dffeas \plif_ifid.instr_l[5] (
	.clk(CPUCLK),
	.d(\instr_l~6_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\plif_ifid.rtnaddr_l[24]~0_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(plif_ifidinstr_l_5),
	.prn(vcc));
// synopsys translate_off
defparam \plif_ifid.instr_l[5] .is_wysiwyg = "true";
defparam \plif_ifid.instr_l[5] .power_up = "low";
// synopsys translate_on

// Location: FF_X55_Y30_N29
dffeas \plif_ifid.instr_l[1] (
	.clk(CPUCLK),
	.d(\instr_l~7_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\plif_ifid.rtnaddr_l[24]~0_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(plif_ifidinstr_l_1),
	.prn(vcc));
// synopsys translate_off
defparam \plif_ifid.instr_l[1] .is_wysiwyg = "true";
defparam \plif_ifid.instr_l[1] .power_up = "low";
// synopsys translate_on

// Location: FF_X56_Y33_N9
dffeas \plif_ifid.instr_l[0] (
	.clk(CPUCLK),
	.d(\instr_l~8_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\plif_ifid.rtnaddr_l[24]~0_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(plif_ifidinstr_l_0),
	.prn(vcc));
// synopsys translate_off
defparam \plif_ifid.instr_l[0] .is_wysiwyg = "true";
defparam \plif_ifid.instr_l[0] .power_up = "low";
// synopsys translate_on

// Location: FF_X60_Y30_N29
dffeas \plif_ifid.instr_l[2] (
	.clk(CPUCLK),
	.d(\instr_l~9_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\plif_ifid.rtnaddr_l[24]~0_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(plif_ifidinstr_l_2),
	.prn(vcc));
// synopsys translate_off
defparam \plif_ifid.instr_l[2] .is_wysiwyg = "true";
defparam \plif_ifid.instr_l[2] .power_up = "low";
// synopsys translate_on

// Location: FF_X55_Y30_N3
dffeas \plif_ifid.instr_l[3] (
	.clk(CPUCLK),
	.d(\instr_l~10_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\plif_ifid.rtnaddr_l[24]~0_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(plif_ifidinstr_l_3),
	.prn(vcc));
// synopsys translate_off
defparam \plif_ifid.instr_l[3] .is_wysiwyg = "true";
defparam \plif_ifid.instr_l[3] .power_up = "low";
// synopsys translate_on

// Location: FF_X56_Y33_N31
dffeas \plif_ifid.instr_l[4] (
	.clk(CPUCLK),
	.d(\instr_l~11_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\plif_ifid.rtnaddr_l[24]~0_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(plif_ifidinstr_l_4),
	.prn(vcc));
// synopsys translate_off
defparam \plif_ifid.instr_l[4] .is_wysiwyg = "true";
defparam \plif_ifid.instr_l[4] .power_up = "low";
// synopsys translate_on

// Location: FF_X59_Y32_N1
dffeas \plif_ifid.instr_l[22] (
	.clk(CPUCLK),
	.d(\instr_l~12_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\plif_ifid.rtnaddr_l[24]~0_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(plif_ifidinstr_l_22),
	.prn(vcc));
// synopsys translate_off
defparam \plif_ifid.instr_l[22] .is_wysiwyg = "true";
defparam \plif_ifid.instr_l[22] .power_up = "low";
// synopsys translate_on

// Location: FF_X59_Y32_N19
dffeas \plif_ifid.instr_l[21] (
	.clk(CPUCLK),
	.d(\instr_l~13_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\plif_ifid.rtnaddr_l[24]~0_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(plif_ifidinstr_l_21),
	.prn(vcc));
// synopsys translate_off
defparam \plif_ifid.instr_l[21] .is_wysiwyg = "true";
defparam \plif_ifid.instr_l[21] .power_up = "low";
// synopsys translate_on

// Location: FF_X59_Y32_N21
dffeas \plif_ifid.instr_l[24] (
	.clk(CPUCLK),
	.d(\instr_l~14_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\plif_ifid.rtnaddr_l[24]~0_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(plif_ifidinstr_l_24),
	.prn(vcc));
// synopsys translate_off
defparam \plif_ifid.instr_l[24] .is_wysiwyg = "true";
defparam \plif_ifid.instr_l[24] .power_up = "low";
// synopsys translate_on

// Location: FF_X59_Y32_N11
dffeas \plif_ifid.instr_l[23] (
	.clk(CPUCLK),
	.d(\instr_l~15_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\plif_ifid.rtnaddr_l[24]~0_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(plif_ifidinstr_l_23),
	.prn(vcc));
// synopsys translate_off
defparam \plif_ifid.instr_l[23] .is_wysiwyg = "true";
defparam \plif_ifid.instr_l[23] .power_up = "low";
// synopsys translate_on

// Location: FF_X59_Y33_N21
dffeas \plif_ifid.instr_l[25] (
	.clk(CPUCLK),
	.d(\instr_l~16_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\plif_ifid.rtnaddr_l[24]~0_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(plif_ifidinstr_l_25),
	.prn(vcc));
// synopsys translate_off
defparam \plif_ifid.instr_l[25] .is_wysiwyg = "true";
defparam \plif_ifid.instr_l[25] .power_up = "low";
// synopsys translate_on

// Location: FF_X59_Y31_N31
dffeas \plif_ifid.instr_l[17] (
	.clk(CPUCLK),
	.d(\instr_l~17_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\plif_ifid.rtnaddr_l[24]~0_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(plif_ifidinstr_l_17),
	.prn(vcc));
// synopsys translate_off
defparam \plif_ifid.instr_l[17] .is_wysiwyg = "true";
defparam \plif_ifid.instr_l[17] .power_up = "low";
// synopsys translate_on

// Location: FF_X59_Y31_N21
dffeas \plif_ifid.instr_l[16] (
	.clk(CPUCLK),
	.d(\instr_l~18_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\plif_ifid.rtnaddr_l[24]~0_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(plif_ifidinstr_l_16),
	.prn(vcc));
// synopsys translate_off
defparam \plif_ifid.instr_l[16] .is_wysiwyg = "true";
defparam \plif_ifid.instr_l[16] .power_up = "low";
// synopsys translate_on

// Location: FF_X59_Y33_N31
dffeas \plif_ifid.instr_l[19] (
	.clk(CPUCLK),
	.d(\instr_l~19_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\plif_ifid.rtnaddr_l[24]~0_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(plif_ifidinstr_l_19),
	.prn(vcc));
// synopsys translate_off
defparam \plif_ifid.instr_l[19] .is_wysiwyg = "true";
defparam \plif_ifid.instr_l[19] .power_up = "low";
// synopsys translate_on

// Location: FF_X59_Y31_N11
dffeas \plif_ifid.instr_l[18] (
	.clk(CPUCLK),
	.d(\instr_l~20_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\plif_ifid.rtnaddr_l[24]~0_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(plif_ifidinstr_l_18),
	.prn(vcc));
// synopsys translate_off
defparam \plif_ifid.instr_l[18] .is_wysiwyg = "true";
defparam \plif_ifid.instr_l[18] .power_up = "low";
// synopsys translate_on

// Location: FF_X59_Y33_N13
dffeas \plif_ifid.instr_l[20] (
	.clk(CPUCLK),
	.d(\instr_l~21_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\plif_ifid.rtnaddr_l[24]~0_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(plif_ifidinstr_l_20),
	.prn(vcc));
// synopsys translate_off
defparam \plif_ifid.instr_l[20] .is_wysiwyg = "true";
defparam \plif_ifid.instr_l[20] .power_up = "low";
// synopsys translate_on

// Location: FF_X59_Y33_N7
dffeas \plif_ifid.instr_l[15] (
	.clk(CPUCLK),
	.d(\instr_l~22_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\plif_ifid.rtnaddr_l[24]~0_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(plif_ifidinstr_l_15),
	.prn(vcc));
// synopsys translate_off
defparam \plif_ifid.instr_l[15] .is_wysiwyg = "true";
defparam \plif_ifid.instr_l[15] .power_up = "low";
// synopsys translate_on

// Location: FF_X57_Y31_N5
dffeas \plif_ifid.instr_l[14] (
	.clk(CPUCLK),
	.d(\instr_l~23_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\plif_ifid.rtnaddr_l[24]~0_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(plif_ifidinstr_l_14),
	.prn(vcc));
// synopsys translate_off
defparam \plif_ifid.instr_l[14] .is_wysiwyg = "true";
defparam \plif_ifid.instr_l[14] .power_up = "low";
// synopsys translate_on

// Location: FF_X56_Y33_N7
dffeas \plif_ifid.instr_l[13] (
	.clk(CPUCLK),
	.d(\instr_l~24_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\plif_ifid.rtnaddr_l[24]~0_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(plif_ifidinstr_l_13),
	.prn(vcc));
// synopsys translate_off
defparam \plif_ifid.instr_l[13] .is_wysiwyg = "true";
defparam \plif_ifid.instr_l[13] .power_up = "low";
// synopsys translate_on

// Location: FF_X57_Y31_N7
dffeas \plif_ifid.instr_l[12] (
	.clk(CPUCLK),
	.d(\instr_l~25_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\plif_ifid.rtnaddr_l[24]~0_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(plif_ifidinstr_l_12),
	.prn(vcc));
// synopsys translate_off
defparam \plif_ifid.instr_l[12] .is_wysiwyg = "true";
defparam \plif_ifid.instr_l[12] .power_up = "low";
// synopsys translate_on

// Location: FF_X56_Y29_N29
dffeas \plif_ifid.instr_l[11] (
	.clk(CPUCLK),
	.d(\instr_l~26_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\plif_ifid.rtnaddr_l[24]~0_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(plif_ifidinstr_l_11),
	.prn(vcc));
// synopsys translate_off
defparam \plif_ifid.instr_l[11] .is_wysiwyg = "true";
defparam \plif_ifid.instr_l[11] .power_up = "low";
// synopsys translate_on

// Location: FF_X58_Y30_N19
dffeas \plif_ifid.instr_l[10] (
	.clk(CPUCLK),
	.d(\instr_l~27_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\plif_ifid.rtnaddr_l[24]~0_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(plif_ifidinstr_l_10),
	.prn(vcc));
// synopsys translate_off
defparam \plif_ifid.instr_l[10] .is_wysiwyg = "true";
defparam \plif_ifid.instr_l[10] .power_up = "low";
// synopsys translate_on

// Location: FF_X57_Y31_N17
dffeas \plif_ifid.instr_l[9] (
	.clk(CPUCLK),
	.d(\instr_l~28_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\plif_ifid.rtnaddr_l[24]~0_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(plif_ifidinstr_l_9),
	.prn(vcc));
// synopsys translate_off
defparam \plif_ifid.instr_l[9] .is_wysiwyg = "true";
defparam \plif_ifid.instr_l[9] .power_up = "low";
// synopsys translate_on

// Location: FF_X56_Y29_N11
dffeas \plif_ifid.instr_l[8] (
	.clk(CPUCLK),
	.d(\instr_l~29_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\plif_ifid.rtnaddr_l[24]~0_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(plif_ifidinstr_l_8),
	.prn(vcc));
// synopsys translate_off
defparam \plif_ifid.instr_l[8] .is_wysiwyg = "true";
defparam \plif_ifid.instr_l[8] .power_up = "low";
// synopsys translate_on

// Location: FF_X55_Y30_N17
dffeas \plif_ifid.instr_l[7] (
	.clk(CPUCLK),
	.d(\instr_l~30_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\plif_ifid.rtnaddr_l[24]~0_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(plif_ifidinstr_l_7),
	.prn(vcc));
// synopsys translate_off
defparam \plif_ifid.instr_l[7] .is_wysiwyg = "true";
defparam \plif_ifid.instr_l[7] .power_up = "low";
// synopsys translate_on

// Location: FF_X55_Y30_N11
dffeas \plif_ifid.instr_l[6] (
	.clk(CPUCLK),
	.d(\instr_l~31_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\plif_ifid.rtnaddr_l[24]~0_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(plif_ifidinstr_l_6),
	.prn(vcc));
// synopsys translate_off
defparam \plif_ifid.instr_l[6] .is_wysiwyg = "true";
defparam \plif_ifid.instr_l[6] .power_up = "low";
// synopsys translate_on

// Location: FF_X53_Y31_N17
dffeas \plif_ifid.rtnaddr_l[31] (
	.clk(CPUCLK),
	.d(\rtnaddr_l~0_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\plif_ifid.rtnaddr_l[24]~0_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(plif_ifidrtnaddr_l_31),
	.prn(vcc));
// synopsys translate_off
defparam \plif_ifid.rtnaddr_l[31] .is_wysiwyg = "true";
defparam \plif_ifid.rtnaddr_l[31] .power_up = "low";
// synopsys translate_on

// Location: FF_X57_Y31_N29
dffeas \plif_ifid.rtnaddr_l[30] (
	.clk(CPUCLK),
	.d(\rtnaddr_l~1_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\plif_ifid.rtnaddr_l[24]~0_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(plif_ifidrtnaddr_l_30),
	.prn(vcc));
// synopsys translate_off
defparam \plif_ifid.rtnaddr_l[30] .is_wysiwyg = "true";
defparam \plif_ifid.rtnaddr_l[30] .power_up = "low";
// synopsys translate_on

// Location: FF_X57_Y31_N25
dffeas \plif_ifid.rtnaddr_l[29] (
	.clk(CPUCLK),
	.d(\rtnaddr_l~2_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\plif_ifid.rtnaddr_l[24]~0_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(plif_ifidrtnaddr_l_29),
	.prn(vcc));
// synopsys translate_off
defparam \plif_ifid.rtnaddr_l[29] .is_wysiwyg = "true";
defparam \plif_ifid.rtnaddr_l[29] .power_up = "low";
// synopsys translate_on

// Location: FF_X52_Y30_N1
dffeas \plif_ifid.rtnaddr_l[28] (
	.clk(CPUCLK),
	.d(\rtnaddr_l~3_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\plif_ifid.rtnaddr_l[24]~0_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(plif_ifidrtnaddr_l_28),
	.prn(vcc));
// synopsys translate_off
defparam \plif_ifid.rtnaddr_l[28] .is_wysiwyg = "true";
defparam \plif_ifid.rtnaddr_l[28] .power_up = "low";
// synopsys translate_on

// Location: FF_X52_Y31_N23
dffeas \plif_ifid.rtnaddr_l[27] (
	.clk(CPUCLK),
	.d(\rtnaddr_l~4_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\plif_ifid.rtnaddr_l[24]~0_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(plif_ifidrtnaddr_l_27),
	.prn(vcc));
// synopsys translate_off
defparam \plif_ifid.rtnaddr_l[27] .is_wysiwyg = "true";
defparam \plif_ifid.rtnaddr_l[27] .power_up = "low";
// synopsys translate_on

// Location: FF_X52_Y31_N5
dffeas \plif_ifid.rtnaddr_l[26] (
	.clk(CPUCLK),
	.d(\rtnaddr_l~5_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\plif_ifid.rtnaddr_l[24]~0_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(plif_ifidrtnaddr_l_26),
	.prn(vcc));
// synopsys translate_off
defparam \plif_ifid.rtnaddr_l[26] .is_wysiwyg = "true";
defparam \plif_ifid.rtnaddr_l[26] .power_up = "low";
// synopsys translate_on

// Location: FF_X52_Y31_N27
dffeas \plif_ifid.rtnaddr_l[25] (
	.clk(CPUCLK),
	.d(\rtnaddr_l~6_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\plif_ifid.rtnaddr_l[24]~0_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(plif_ifidrtnaddr_l_25),
	.prn(vcc));
// synopsys translate_off
defparam \plif_ifid.rtnaddr_l[25] .is_wysiwyg = "true";
defparam \plif_ifid.rtnaddr_l[25] .power_up = "low";
// synopsys translate_on

// Location: FF_X52_Y31_N9
dffeas \plif_ifid.rtnaddr_l[24] (
	.clk(CPUCLK),
	.d(\rtnaddr_l~7_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\plif_ifid.rtnaddr_l[24]~0_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(plif_ifidrtnaddr_l_24),
	.prn(vcc));
// synopsys translate_off
defparam \plif_ifid.rtnaddr_l[24] .is_wysiwyg = "true";
defparam \plif_ifid.rtnaddr_l[24] .power_up = "low";
// synopsys translate_on

// Location: FF_X52_Y31_N31
dffeas \plif_ifid.rtnaddr_l[23] (
	.clk(CPUCLK),
	.d(\rtnaddr_l~8_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\plif_ifid.rtnaddr_l[24]~0_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(plif_ifidrtnaddr_l_23),
	.prn(vcc));
// synopsys translate_off
defparam \plif_ifid.rtnaddr_l[23] .is_wysiwyg = "true";
defparam \plif_ifid.rtnaddr_l[23] .power_up = "low";
// synopsys translate_on

// Location: FF_X52_Y31_N29
dffeas \plif_ifid.rtnaddr_l[22] (
	.clk(CPUCLK),
	.d(\rtnaddr_l~9_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\plif_ifid.rtnaddr_l[24]~0_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(plif_ifidrtnaddr_l_22),
	.prn(vcc));
// synopsys translate_off
defparam \plif_ifid.rtnaddr_l[22] .is_wysiwyg = "true";
defparam \plif_ifid.rtnaddr_l[22] .power_up = "low";
// synopsys translate_on

// Location: FF_X52_Y30_N15
dffeas \plif_ifid.rtnaddr_l[21] (
	.clk(CPUCLK),
	.d(\rtnaddr_l~10_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\plif_ifid.rtnaddr_l[24]~0_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(plif_ifidrtnaddr_l_21),
	.prn(vcc));
// synopsys translate_off
defparam \plif_ifid.rtnaddr_l[21] .is_wysiwyg = "true";
defparam \plif_ifid.rtnaddr_l[21] .power_up = "low";
// synopsys translate_on

// Location: FF_X52_Y30_N25
dffeas \plif_ifid.rtnaddr_l[20] (
	.clk(CPUCLK),
	.d(\rtnaddr_l~11_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\plif_ifid.rtnaddr_l[24]~0_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(plif_ifidrtnaddr_l_20),
	.prn(vcc));
// synopsys translate_off
defparam \plif_ifid.rtnaddr_l[20] .is_wysiwyg = "true";
defparam \plif_ifid.rtnaddr_l[20] .power_up = "low";
// synopsys translate_on

// Location: FF_X53_Y31_N27
dffeas \plif_ifid.rtnaddr_l[19] (
	.clk(CPUCLK),
	.d(\rtnaddr_l~12_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\plif_ifid.rtnaddr_l[24]~0_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(plif_ifidrtnaddr_l_19),
	.prn(vcc));
// synopsys translate_off
defparam \plif_ifid.rtnaddr_l[19] .is_wysiwyg = "true";
defparam \plif_ifid.rtnaddr_l[19] .power_up = "low";
// synopsys translate_on

// Location: FF_X53_Y31_N21
dffeas \plif_ifid.rtnaddr_l[18] (
	.clk(CPUCLK),
	.d(\rtnaddr_l~13_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\plif_ifid.rtnaddr_l[24]~0_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(plif_ifidrtnaddr_l_18),
	.prn(vcc));
// synopsys translate_off
defparam \plif_ifid.rtnaddr_l[18] .is_wysiwyg = "true";
defparam \plif_ifid.rtnaddr_l[18] .power_up = "low";
// synopsys translate_on

// Location: FF_X52_Y31_N19
dffeas \plif_ifid.rtnaddr_l[17] (
	.clk(CPUCLK),
	.d(\rtnaddr_l~14_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\plif_ifid.rtnaddr_l[24]~0_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(plif_ifidrtnaddr_l_17),
	.prn(vcc));
// synopsys translate_off
defparam \plif_ifid.rtnaddr_l[17] .is_wysiwyg = "true";
defparam \plif_ifid.rtnaddr_l[17] .power_up = "low";
// synopsys translate_on

// Location: FF_X53_Y31_N31
dffeas \plif_ifid.rtnaddr_l[16] (
	.clk(CPUCLK),
	.d(\rtnaddr_l~15_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\plif_ifid.rtnaddr_l[24]~0_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(plif_ifidrtnaddr_l_16),
	.prn(vcc));
// synopsys translate_off
defparam \plif_ifid.rtnaddr_l[16] .is_wysiwyg = "true";
defparam \plif_ifid.rtnaddr_l[16] .power_up = "low";
// synopsys translate_on

// Location: FF_X54_Y30_N5
dffeas \plif_ifid.rtnaddr_l[15] (
	.clk(CPUCLK),
	.d(\rtnaddr_l~16_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\plif_ifid.rtnaddr_l[24]~0_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(plif_ifidrtnaddr_l_15),
	.prn(vcc));
// synopsys translate_off
defparam \plif_ifid.rtnaddr_l[15] .is_wysiwyg = "true";
defparam \plif_ifid.rtnaddr_l[15] .power_up = "low";
// synopsys translate_on

// Location: FF_X53_Y29_N1
dffeas \plif_ifid.rtnaddr_l[14] (
	.clk(CPUCLK),
	.d(\rtnaddr_l~17_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\plif_ifid.rtnaddr_l[24]~0_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(plif_ifidrtnaddr_l_14),
	.prn(vcc));
// synopsys translate_off
defparam \plif_ifid.rtnaddr_l[14] .is_wysiwyg = "true";
defparam \plif_ifid.rtnaddr_l[14] .power_up = "low";
// synopsys translate_on

// Location: FF_X53_Y31_N25
dffeas \plif_ifid.rtnaddr_l[13] (
	.clk(CPUCLK),
	.d(\rtnaddr_l~18_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\plif_ifid.rtnaddr_l[24]~0_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(plif_ifidrtnaddr_l_13),
	.prn(vcc));
// synopsys translate_off
defparam \plif_ifid.rtnaddr_l[13] .is_wysiwyg = "true";
defparam \plif_ifid.rtnaddr_l[13] .power_up = "low";
// synopsys translate_on

// Location: FF_X53_Y31_N15
dffeas \plif_ifid.rtnaddr_l[12] (
	.clk(CPUCLK),
	.d(\rtnaddr_l~19_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\plif_ifid.rtnaddr_l[24]~0_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(plif_ifidrtnaddr_l_12),
	.prn(vcc));
// synopsys translate_off
defparam \plif_ifid.rtnaddr_l[12] .is_wysiwyg = "true";
defparam \plif_ifid.rtnaddr_l[12] .power_up = "low";
// synopsys translate_on

// Location: FF_X53_Y31_N13
dffeas \plif_ifid.rtnaddr_l[11] (
	.clk(CPUCLK),
	.d(\rtnaddr_l~20_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\plif_ifid.rtnaddr_l[24]~0_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(plif_ifidrtnaddr_l_11),
	.prn(vcc));
// synopsys translate_off
defparam \plif_ifid.rtnaddr_l[11] .is_wysiwyg = "true";
defparam \plif_ifid.rtnaddr_l[11] .power_up = "low";
// synopsys translate_on

// Location: FF_X53_Y31_N11
dffeas \plif_ifid.rtnaddr_l[10] (
	.clk(CPUCLK),
	.d(\rtnaddr_l~21_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\plif_ifid.rtnaddr_l[24]~0_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(plif_ifidrtnaddr_l_10),
	.prn(vcc));
// synopsys translate_off
defparam \plif_ifid.rtnaddr_l[10] .is_wysiwyg = "true";
defparam \plif_ifid.rtnaddr_l[10] .power_up = "low";
// synopsys translate_on

// Location: FF_X57_Y31_N3
dffeas \plif_ifid.rtnaddr_l[9] (
	.clk(CPUCLK),
	.d(\rtnaddr_l~22_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\plif_ifid.rtnaddr_l[24]~0_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(plif_ifidrtnaddr_l_9),
	.prn(vcc));
// synopsys translate_off
defparam \plif_ifid.rtnaddr_l[9] .is_wysiwyg = "true";
defparam \plif_ifid.rtnaddr_l[9] .power_up = "low";
// synopsys translate_on

// Location: FF_X57_Y31_N21
dffeas \plif_ifid.rtnaddr_l[8] (
	.clk(CPUCLK),
	.d(\rtnaddr_l~23_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\plif_ifid.rtnaddr_l[24]~0_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(plif_ifidrtnaddr_l_8),
	.prn(vcc));
// synopsys translate_off
defparam \plif_ifid.rtnaddr_l[8] .is_wysiwyg = "true";
defparam \plif_ifid.rtnaddr_l[8] .power_up = "low";
// synopsys translate_on

// Location: FF_X53_Y31_N9
dffeas \plif_ifid.rtnaddr_l[7] (
	.clk(CPUCLK),
	.d(\rtnaddr_l~24_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\plif_ifid.rtnaddr_l[24]~0_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(plif_ifidrtnaddr_l_7),
	.prn(vcc));
// synopsys translate_off
defparam \plif_ifid.rtnaddr_l[7] .is_wysiwyg = "true";
defparam \plif_ifid.rtnaddr_l[7] .power_up = "low";
// synopsys translate_on

// Location: FF_X57_Y31_N11
dffeas \plif_ifid.rtnaddr_l[6] (
	.clk(CPUCLK),
	.d(\rtnaddr_l~25_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\plif_ifid.rtnaddr_l[24]~0_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(plif_ifidrtnaddr_l_6),
	.prn(vcc));
// synopsys translate_off
defparam \plif_ifid.rtnaddr_l[6] .is_wysiwyg = "true";
defparam \plif_ifid.rtnaddr_l[6] .power_up = "low";
// synopsys translate_on

// Location: FF_X53_Y31_N23
dffeas \plif_ifid.rtnaddr_l[5] (
	.clk(CPUCLK),
	.d(\rtnaddr_l~26_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\plif_ifid.rtnaddr_l[24]~0_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(plif_ifidrtnaddr_l_5),
	.prn(vcc));
// synopsys translate_off
defparam \plif_ifid.rtnaddr_l[5] .is_wysiwyg = "true";
defparam \plif_ifid.rtnaddr_l[5] .power_up = "low";
// synopsys translate_on

// Location: FF_X52_Y30_N23
dffeas \plif_ifid.rtnaddr_l[2] (
	.clk(CPUCLK),
	.d(\rtnaddr_l~27_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\plif_ifid.rtnaddr_l[24]~0_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(plif_ifidrtnaddr_l_2),
	.prn(vcc));
// synopsys translate_off
defparam \plif_ifid.rtnaddr_l[2] .is_wysiwyg = "true";
defparam \plif_ifid.rtnaddr_l[2] .power_up = "low";
// synopsys translate_on

// Location: FF_X53_Y31_N29
dffeas \plif_ifid.rtnaddr_l[1] (
	.clk(CPUCLK),
	.d(\rtnaddr_l~28_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\plif_ifid.rtnaddr_l[24]~0_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(plif_ifidrtnaddr_l_1),
	.prn(vcc));
// synopsys translate_off
defparam \plif_ifid.rtnaddr_l[1] .is_wysiwyg = "true";
defparam \plif_ifid.rtnaddr_l[1] .power_up = "low";
// synopsys translate_on

// Location: FF_X53_Y31_N7
dffeas \plif_ifid.rtnaddr_l[0] (
	.clk(CPUCLK),
	.d(\rtnaddr_l~29_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\plif_ifid.rtnaddr_l[24]~0_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(plif_ifidrtnaddr_l_0),
	.prn(vcc));
// synopsys translate_off
defparam \plif_ifid.rtnaddr_l[0] .is_wysiwyg = "true";
defparam \plif_ifid.rtnaddr_l[0] .power_up = "low";
// synopsys translate_on

// Location: FF_X57_Y31_N13
dffeas \plif_ifid.rtnaddr_l[4] (
	.clk(CPUCLK),
	.d(\rtnaddr_l~30_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\plif_ifid.rtnaddr_l[24]~0_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(plif_ifidrtnaddr_l_4),
	.prn(vcc));
// synopsys translate_off
defparam \plif_ifid.rtnaddr_l[4] .is_wysiwyg = "true";
defparam \plif_ifid.rtnaddr_l[4] .power_up = "low";
// synopsys translate_on

// Location: FF_X57_Y31_N23
dffeas \plif_ifid.rtnaddr_l[3] (
	.clk(CPUCLK),
	.d(\rtnaddr_l~31_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\plif_ifid.rtnaddr_l[24]~0_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(plif_ifidrtnaddr_l_3),
	.prn(vcc));
// synopsys translate_off
defparam \plif_ifid.rtnaddr_l[3] .is_wysiwyg = "true";
defparam \plif_ifid.rtnaddr_l[3] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X59_Y30_N10
cycloneive_lcell_comb \instr_l~0 (
// Equation(s):
// \instr_l~0_combout  = (!ifid_sRST1 & ((ccifiwait_0 & (instr_31)) # (!ccifiwait_0 & ((ramiframload_31)))))

	.dataa(instr_31),
	.datab(ramiframload_31),
	.datac(ccifiwait_0),
	.datad(ifid_sRST),
	.cin(gnd),
	.combout(\instr_l~0_combout ),
	.cout());
// synopsys translate_off
defparam \instr_l~0 .lut_mask = 16'h00AC;
defparam \instr_l~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y33_N4
cycloneive_lcell_comb \plif_ifid.rtnaddr_l[24]~0 (
// Equation(s):
// \plif_ifid.rtnaddr_l[24]~0_combout  = (ifid_sRST1) # (ifid_en)

	.dataa(gnd),
	.datab(ifid_sRST),
	.datac(gnd),
	.datad(ifid_en),
	.cin(gnd),
	.combout(\plif_ifid.rtnaddr_l[24]~0_combout ),
	.cout());
// synopsys translate_off
defparam \plif_ifid.rtnaddr_l[24]~0 .lut_mask = 16'hFFCC;
defparam \plif_ifid.rtnaddr_l[24]~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y30_N8
cycloneive_lcell_comb \instr_l~1 (
// Equation(s):
// \instr_l~1_combout  = (!ifid_sRST1 & ((ccifiwait_0 & (instr_29)) # (!ccifiwait_0 & ((ramiframload_29)))))

	.dataa(instr_29),
	.datab(ifid_sRST),
	.datac(ccifiwait_0),
	.datad(ramiframload_29),
	.cin(gnd),
	.combout(\instr_l~1_combout ),
	.cout());
// synopsys translate_off
defparam \instr_l~1 .lut_mask = 16'h2320;
defparam \instr_l~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y30_N6
cycloneive_lcell_comb \instr_l~2 (
// Equation(s):
// \instr_l~2_combout  = (!ifid_sRST1 & ((ccifiwait_0 & ((instr_27))) # (!ccifiwait_0 & (ramiframload_27))))

	.dataa(ramiframload_27),
	.datab(instr_27),
	.datac(ccifiwait_0),
	.datad(ifid_sRST),
	.cin(gnd),
	.combout(\instr_l~2_combout ),
	.cout());
// synopsys translate_off
defparam \instr_l~2 .lut_mask = 16'h00CA;
defparam \instr_l~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y30_N24
cycloneive_lcell_comb \instr_l~3 (
// Equation(s):
// \instr_l~3_combout  = (!ifid_sRST1 & ((ccifiwait_0 & ((instr_26))) # (!ccifiwait_0 & (ramiframload_26))))

	.dataa(ramiframload_26),
	.datab(ccifiwait_0),
	.datac(instr_26),
	.datad(ifid_sRST),
	.cin(gnd),
	.combout(\instr_l~3_combout ),
	.cout());
// synopsys translate_off
defparam \instr_l~3 .lut_mask = 16'h00E2;
defparam \instr_l~3 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y30_N6
cycloneive_lcell_comb \instr_l~4 (
// Equation(s):
// \instr_l~4_combout  = (!ifid_sRST1 & ((ccifiwait_0 & ((instr_28))) # (!ccifiwait_0 & (ramiframload_28))))

	.dataa(ramiframload_28),
	.datab(ccifiwait_0),
	.datac(instr_28),
	.datad(ifid_sRST),
	.cin(gnd),
	.combout(\instr_l~4_combout ),
	.cout());
// synopsys translate_off
defparam \instr_l~4 .lut_mask = 16'h00E2;
defparam \instr_l~4 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y30_N30
cycloneive_lcell_comb \instr_l~5 (
// Equation(s):
// \instr_l~5_combout  = (!ifid_sRST1 & ((ccifiwait_0 & (instr_30)) # (!ccifiwait_0 & ((ramiframload_30)))))

	.dataa(instr_30),
	.datab(ifid_sRST),
	.datac(ccifiwait_0),
	.datad(ramiframload_30),
	.cin(gnd),
	.combout(\instr_l~5_combout ),
	.cout());
// synopsys translate_off
defparam \instr_l~5 .lut_mask = 16'h2320;
defparam \instr_l~5 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y30_N28
cycloneive_lcell_comb \instr_l~6 (
// Equation(s):
// \instr_l~6_combout  = (!ifid_sRST1 & ((ccifiwait_0 & ((instr_5))) # (!ccifiwait_0 & (ramiframload_5))))

	.dataa(ifid_sRST),
	.datab(ramiframload_5),
	.datac(instr_5),
	.datad(ccifiwait_0),
	.cin(gnd),
	.combout(\instr_l~6_combout ),
	.cout());
// synopsys translate_off
defparam \instr_l~6 .lut_mask = 16'h5044;
defparam \instr_l~6 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y30_N28
cycloneive_lcell_comb \instr_l~7 (
// Equation(s):
// \instr_l~7_combout  = (!ifid_sRST1 & ((ccifiwait_0 & ((instr_1))) # (!ccifiwait_0 & (ramiframload_1))))

	.dataa(ccifiwait_0),
	.datab(ramiframload_1),
	.datac(instr_1),
	.datad(ifid_sRST),
	.cin(gnd),
	.combout(\instr_l~7_combout ),
	.cout());
// synopsys translate_off
defparam \instr_l~7 .lut_mask = 16'h00E4;
defparam \instr_l~7 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y33_N8
cycloneive_lcell_comb \instr_l~8 (
// Equation(s):
// \instr_l~8_combout  = (!ifid_sRST1 & ((ccifiwait_0 & ((instr_0))) # (!ccifiwait_0 & (ramiframload_0))))

	.dataa(ccifiwait_0),
	.datab(ramiframload_0),
	.datac(instr_0),
	.datad(ifid_sRST),
	.cin(gnd),
	.combout(\instr_l~8_combout ),
	.cout());
// synopsys translate_off
defparam \instr_l~8 .lut_mask = 16'h00E4;
defparam \instr_l~8 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y30_N28
cycloneive_lcell_comb \instr_l~9 (
// Equation(s):
// \instr_l~9_combout  = (!ifid_sRST1 & ((ccifiwait_0 & ((instr_2))) # (!ccifiwait_0 & (ramiframload_2))))

	.dataa(ramiframload_2),
	.datab(ccifiwait_0),
	.datac(instr_2),
	.datad(ifid_sRST),
	.cin(gnd),
	.combout(\instr_l~9_combout ),
	.cout());
// synopsys translate_off
defparam \instr_l~9 .lut_mask = 16'h00E2;
defparam \instr_l~9 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y30_N2
cycloneive_lcell_comb \instr_l~10 (
// Equation(s):
// \instr_l~10_combout  = (!ifid_sRST1 & ((ccifiwait_0 & ((instr_3))) # (!ccifiwait_0 & (ramiframload_3))))

	.dataa(ccifiwait_0),
	.datab(ramiframload_3),
	.datac(instr_3),
	.datad(ifid_sRST),
	.cin(gnd),
	.combout(\instr_l~10_combout ),
	.cout());
// synopsys translate_off
defparam \instr_l~10 .lut_mask = 16'h00E4;
defparam \instr_l~10 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y33_N30
cycloneive_lcell_comb \instr_l~11 (
// Equation(s):
// \instr_l~11_combout  = (!ifid_sRST1 & ((ccifiwait_0 & ((instr_4))) # (!ccifiwait_0 & (ramiframload_4))))

	.dataa(ramiframload_4),
	.datab(ifid_sRST),
	.datac(ccifiwait_0),
	.datad(instr_4),
	.cin(gnd),
	.combout(\instr_l~11_combout ),
	.cout());
// synopsys translate_off
defparam \instr_l~11 .lut_mask = 16'h3202;
defparam \instr_l~11 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y32_N0
cycloneive_lcell_comb \instr_l~12 (
// Equation(s):
// \instr_l~12_combout  = (!ifid_sRST1 & ((ccifiwait_0 & ((instr_22))) # (!ccifiwait_0 & (ramiframload_22))))

	.dataa(ifid_sRST),
	.datab(ccifiwait_0),
	.datac(ramiframload_22),
	.datad(instr_22),
	.cin(gnd),
	.combout(\instr_l~12_combout ),
	.cout());
// synopsys translate_off
defparam \instr_l~12 .lut_mask = 16'h5410;
defparam \instr_l~12 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y32_N18
cycloneive_lcell_comb \instr_l~13 (
// Equation(s):
// \instr_l~13_combout  = (!ifid_sRST1 & ((ccifiwait_0 & ((instr_21))) # (!ccifiwait_0 & (ramiframload_21))))

	.dataa(ifid_sRST),
	.datab(ramiframload_21),
	.datac(instr_21),
	.datad(ccifiwait_0),
	.cin(gnd),
	.combout(\instr_l~13_combout ),
	.cout());
// synopsys translate_off
defparam \instr_l~13 .lut_mask = 16'h5044;
defparam \instr_l~13 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y32_N20
cycloneive_lcell_comb \instr_l~14 (
// Equation(s):
// \instr_l~14_combout  = (!ifid_sRST1 & ((ccifiwait_0 & ((instr_24))) # (!ccifiwait_0 & (ramiframload_24))))

	.dataa(ifid_sRST),
	.datab(ccifiwait_0),
	.datac(ramiframload_24),
	.datad(instr_24),
	.cin(gnd),
	.combout(\instr_l~14_combout ),
	.cout());
// synopsys translate_off
defparam \instr_l~14 .lut_mask = 16'h5410;
defparam \instr_l~14 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y32_N10
cycloneive_lcell_comb \instr_l~15 (
// Equation(s):
// \instr_l~15_combout  = (!ifid_sRST1 & ((ccifiwait_0 & ((instr_23))) # (!ccifiwait_0 & (ramiframload_23))))

	.dataa(ramiframload_23),
	.datab(ccifiwait_0),
	.datac(instr_23),
	.datad(ifid_sRST),
	.cin(gnd),
	.combout(\instr_l~15_combout ),
	.cout());
// synopsys translate_off
defparam \instr_l~15 .lut_mask = 16'h00E2;
defparam \instr_l~15 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y33_N20
cycloneive_lcell_comb \instr_l~16 (
// Equation(s):
// \instr_l~16_combout  = (!ifid_sRST1 & ((ccifiwait_0 & ((instr_25))) # (!ccifiwait_0 & (ramiframload_25))))

	.dataa(ramiframload_25),
	.datab(ifid_sRST),
	.datac(instr_25),
	.datad(ccifiwait_0),
	.cin(gnd),
	.combout(\instr_l~16_combout ),
	.cout());
// synopsys translate_off
defparam \instr_l~16 .lut_mask = 16'h3022;
defparam \instr_l~16 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y31_N30
cycloneive_lcell_comb \instr_l~17 (
// Equation(s):
// \instr_l~17_combout  = (!ifid_sRST1 & ((ccifiwait_0 & ((instr_17))) # (!ccifiwait_0 & (ramiframload_17))))

	.dataa(ccifiwait_0),
	.datab(ramiframload_17),
	.datac(instr_17),
	.datad(ifid_sRST),
	.cin(gnd),
	.combout(\instr_l~17_combout ),
	.cout());
// synopsys translate_off
defparam \instr_l~17 .lut_mask = 16'h00E4;
defparam \instr_l~17 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y31_N20
cycloneive_lcell_comb \instr_l~18 (
// Equation(s):
// \instr_l~18_combout  = (!ifid_sRST1 & ((ccifiwait_0 & (instr_16)) # (!ccifiwait_0 & ((ramiframload_16)))))

	.dataa(ccifiwait_0),
	.datab(ifid_sRST),
	.datac(instr_16),
	.datad(ramiframload_16),
	.cin(gnd),
	.combout(\instr_l~18_combout ),
	.cout());
// synopsys translate_off
defparam \instr_l~18 .lut_mask = 16'h3120;
defparam \instr_l~18 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y33_N30
cycloneive_lcell_comb \instr_l~19 (
// Equation(s):
// \instr_l~19_combout  = (!ifid_sRST1 & ((ccifiwait_0 & (instr_19)) # (!ccifiwait_0 & ((ramiframload_19)))))

	.dataa(instr_19),
	.datab(ifid_sRST),
	.datac(ramiframload_19),
	.datad(ccifiwait_0),
	.cin(gnd),
	.combout(\instr_l~19_combout ),
	.cout());
// synopsys translate_off
defparam \instr_l~19 .lut_mask = 16'h2230;
defparam \instr_l~19 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y31_N10
cycloneive_lcell_comb \instr_l~20 (
// Equation(s):
// \instr_l~20_combout  = (!ifid_sRST1 & ((ccifiwait_0 & ((instr_18))) # (!ccifiwait_0 & (ramiframload_18))))

	.dataa(ccifiwait_0),
	.datab(ramiframload_18),
	.datac(instr_18),
	.datad(ifid_sRST),
	.cin(gnd),
	.combout(\instr_l~20_combout ),
	.cout());
// synopsys translate_off
defparam \instr_l~20 .lut_mask = 16'h00E4;
defparam \instr_l~20 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y33_N12
cycloneive_lcell_comb \instr_l~21 (
// Equation(s):
// \instr_l~21_combout  = (!ifid_sRST1 & ((ccifiwait_0 & (instr_20)) # (!ccifiwait_0 & ((ramiframload_20)))))

	.dataa(ccifiwait_0),
	.datab(instr_20),
	.datac(ramiframload_20),
	.datad(ifid_sRST),
	.cin(gnd),
	.combout(\instr_l~21_combout ),
	.cout());
// synopsys translate_off
defparam \instr_l~21 .lut_mask = 16'h00D8;
defparam \instr_l~21 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y33_N6
cycloneive_lcell_comb \instr_l~22 (
// Equation(s):
// \instr_l~22_combout  = (!ifid_sRST1 & ((ccifiwait_0 & ((instr_15))) # (!ccifiwait_0 & (ramiframload_15))))

	.dataa(ifid_sRST),
	.datab(ramiframload_15),
	.datac(instr_15),
	.datad(ccifiwait_0),
	.cin(gnd),
	.combout(\instr_l~22_combout ),
	.cout());
// synopsys translate_off
defparam \instr_l~22 .lut_mask = 16'h5044;
defparam \instr_l~22 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y31_N4
cycloneive_lcell_comb \instr_l~23 (
// Equation(s):
// \instr_l~23_combout  = (!ifid_sRST1 & ((ccifiwait_0 & ((instr_14))) # (!ccifiwait_0 & (ramiframload_14))))

	.dataa(ccifiwait_0),
	.datab(ramiframload_14),
	.datac(instr_14),
	.datad(ifid_sRST),
	.cin(gnd),
	.combout(\instr_l~23_combout ),
	.cout());
// synopsys translate_off
defparam \instr_l~23 .lut_mask = 16'h00E4;
defparam \instr_l~23 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y33_N6
cycloneive_lcell_comb \instr_l~24 (
// Equation(s):
// \instr_l~24_combout  = (!ifid_sRST1 & ((ccifiwait_0 & ((instr_13))) # (!ccifiwait_0 & (ramiframload_13))))

	.dataa(ccifiwait_0),
	.datab(ramiframload_13),
	.datac(instr_13),
	.datad(ifid_sRST),
	.cin(gnd),
	.combout(\instr_l~24_combout ),
	.cout());
// synopsys translate_off
defparam \instr_l~24 .lut_mask = 16'h00E4;
defparam \instr_l~24 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y31_N6
cycloneive_lcell_comb \instr_l~25 (
// Equation(s):
// \instr_l~25_combout  = (!ifid_sRST1 & ((ccifiwait_0 & ((instr_12))) # (!ccifiwait_0 & (ramiframload_12))))

	.dataa(ccifiwait_0),
	.datab(ramiframload_12),
	.datac(instr_12),
	.datad(ifid_sRST),
	.cin(gnd),
	.combout(\instr_l~25_combout ),
	.cout());
// synopsys translate_off
defparam \instr_l~25 .lut_mask = 16'h00E4;
defparam \instr_l~25 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y29_N28
cycloneive_lcell_comb \instr_l~26 (
// Equation(s):
// \instr_l~26_combout  = (!ifid_sRST1 & ((ccifiwait_0 & ((instr_11))) # (!ccifiwait_0 & (ramiframload_11))))

	.dataa(ramiframload_11),
	.datab(ifid_sRST),
	.datac(instr_11),
	.datad(ccifiwait_0),
	.cin(gnd),
	.combout(\instr_l~26_combout ),
	.cout());
// synopsys translate_off
defparam \instr_l~26 .lut_mask = 16'h3022;
defparam \instr_l~26 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y30_N18
cycloneive_lcell_comb \instr_l~27 (
// Equation(s):
// \instr_l~27_combout  = (!ifid_sRST1 & ((ccifiwait_0 & ((instr_10))) # (!ccifiwait_0 & (ramiframload_10))))

	.dataa(ramiframload_10),
	.datab(ccifiwait_0),
	.datac(instr_10),
	.datad(ifid_sRST),
	.cin(gnd),
	.combout(\instr_l~27_combout ),
	.cout());
// synopsys translate_off
defparam \instr_l~27 .lut_mask = 16'h00E2;
defparam \instr_l~27 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y31_N16
cycloneive_lcell_comb \instr_l~28 (
// Equation(s):
// \instr_l~28_combout  = (!ifid_sRST1 & ((ccifiwait_0 & (instr_9)) # (!ccifiwait_0 & ((ramiframload_9)))))

	.dataa(ifid_sRST),
	.datab(ccifiwait_0),
	.datac(instr_9),
	.datad(ramiframload_9),
	.cin(gnd),
	.combout(\instr_l~28_combout ),
	.cout());
// synopsys translate_off
defparam \instr_l~28 .lut_mask = 16'h5140;
defparam \instr_l~28 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y29_N10
cycloneive_lcell_comb \instr_l~29 (
// Equation(s):
// \instr_l~29_combout  = (!ifid_sRST1 & ((ccifiwait_0 & ((instr_8))) # (!ccifiwait_0 & (ramiframload_8))))

	.dataa(ramiframload_8),
	.datab(ifid_sRST),
	.datac(instr_8),
	.datad(ccifiwait_0),
	.cin(gnd),
	.combout(\instr_l~29_combout ),
	.cout());
// synopsys translate_off
defparam \instr_l~29 .lut_mask = 16'h3022;
defparam \instr_l~29 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y30_N16
cycloneive_lcell_comb \instr_l~30 (
// Equation(s):
// \instr_l~30_combout  = (!ifid_sRST1 & ((ccifiwait_0 & (instr_7)) # (!ccifiwait_0 & ((ramiframload_7)))))

	.dataa(ifid_sRST),
	.datab(ccifiwait_0),
	.datac(instr_7),
	.datad(ramiframload_7),
	.cin(gnd),
	.combout(\instr_l~30_combout ),
	.cout());
// synopsys translate_off
defparam \instr_l~30 .lut_mask = 16'h5140;
defparam \instr_l~30 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y30_N10
cycloneive_lcell_comb \instr_l~31 (
// Equation(s):
// \instr_l~31_combout  = (!ifid_sRST1 & ((ccifiwait_0 & ((instr_6))) # (!ccifiwait_0 & (ramiframload_6))))

	.dataa(ccifiwait_0),
	.datab(ramiframload_6),
	.datac(instr_6),
	.datad(ifid_sRST),
	.cin(gnd),
	.combout(\instr_l~31_combout ),
	.cout());
// synopsys translate_off
defparam \instr_l~31 .lut_mask = 16'h00E4;
defparam \instr_l~31 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y31_N16
cycloneive_lcell_comb \rtnaddr_l~0 (
// Equation(s):
// \rtnaddr_l~0_combout  = (!ifid_sRST1 & pcifrtnaddr_31)

	.dataa(gnd),
	.datab(gnd),
	.datac(ifid_sRST),
	.datad(pcifrtnaddr_31),
	.cin(gnd),
	.combout(\rtnaddr_l~0_combout ),
	.cout());
// synopsys translate_off
defparam \rtnaddr_l~0 .lut_mask = 16'h0F00;
defparam \rtnaddr_l~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y31_N28
cycloneive_lcell_comb \rtnaddr_l~1 (
// Equation(s):
// \rtnaddr_l~1_combout  = (!ifid_sRST1 & pcifrtnaddr_30)

	.dataa(ifid_sRST),
	.datab(gnd),
	.datac(gnd),
	.datad(pcifrtnaddr_30),
	.cin(gnd),
	.combout(\rtnaddr_l~1_combout ),
	.cout());
// synopsys translate_off
defparam \rtnaddr_l~1 .lut_mask = 16'h5500;
defparam \rtnaddr_l~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y31_N24
cycloneive_lcell_comb \rtnaddr_l~2 (
// Equation(s):
// \rtnaddr_l~2_combout  = (pcifrtnaddr_29 & !ifid_sRST1)

	.dataa(gnd),
	.datab(pcifrtnaddr_29),
	.datac(gnd),
	.datad(ifid_sRST),
	.cin(gnd),
	.combout(\rtnaddr_l~2_combout ),
	.cout());
// synopsys translate_off
defparam \rtnaddr_l~2 .lut_mask = 16'h00CC;
defparam \rtnaddr_l~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X52_Y30_N0
cycloneive_lcell_comb \rtnaddr_l~3 (
// Equation(s):
// \rtnaddr_l~3_combout  = (!ifid_sRST1 & pcifrtnaddr_28)

	.dataa(ifid_sRST),
	.datab(gnd),
	.datac(gnd),
	.datad(pcifrtnaddr_28),
	.cin(gnd),
	.combout(\rtnaddr_l~3_combout ),
	.cout());
// synopsys translate_off
defparam \rtnaddr_l~3 .lut_mask = 16'h5500;
defparam \rtnaddr_l~3 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X52_Y31_N22
cycloneive_lcell_comb \rtnaddr_l~4 (
// Equation(s):
// \rtnaddr_l~4_combout  = (pcifrtnaddr_27 & !ifid_sRST1)

	.dataa(gnd),
	.datab(gnd),
	.datac(pcifrtnaddr_27),
	.datad(ifid_sRST),
	.cin(gnd),
	.combout(\rtnaddr_l~4_combout ),
	.cout());
// synopsys translate_off
defparam \rtnaddr_l~4 .lut_mask = 16'h00F0;
defparam \rtnaddr_l~4 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X52_Y31_N4
cycloneive_lcell_comb \rtnaddr_l~5 (
// Equation(s):
// \rtnaddr_l~5_combout  = (pcifrtnaddr_26 & !ifid_sRST1)

	.dataa(gnd),
	.datab(gnd),
	.datac(pcifrtnaddr_26),
	.datad(ifid_sRST),
	.cin(gnd),
	.combout(\rtnaddr_l~5_combout ),
	.cout());
// synopsys translate_off
defparam \rtnaddr_l~5 .lut_mask = 16'h00F0;
defparam \rtnaddr_l~5 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X52_Y31_N26
cycloneive_lcell_comb \rtnaddr_l~6 (
// Equation(s):
// \rtnaddr_l~6_combout  = (!ifid_sRST1 & pcifrtnaddr_25)

	.dataa(gnd),
	.datab(ifid_sRST),
	.datac(gnd),
	.datad(pcifrtnaddr_25),
	.cin(gnd),
	.combout(\rtnaddr_l~6_combout ),
	.cout());
// synopsys translate_off
defparam \rtnaddr_l~6 .lut_mask = 16'h3300;
defparam \rtnaddr_l~6 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X52_Y31_N8
cycloneive_lcell_comb \rtnaddr_l~7 (
// Equation(s):
// \rtnaddr_l~7_combout  = (!ifid_sRST1 & pcifrtnaddr_24)

	.dataa(gnd),
	.datab(ifid_sRST),
	.datac(gnd),
	.datad(pcifrtnaddr_24),
	.cin(gnd),
	.combout(\rtnaddr_l~7_combout ),
	.cout());
// synopsys translate_off
defparam \rtnaddr_l~7 .lut_mask = 16'h3300;
defparam \rtnaddr_l~7 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X52_Y31_N30
cycloneive_lcell_comb \rtnaddr_l~8 (
// Equation(s):
// \rtnaddr_l~8_combout  = (pcifrtnaddr_23 & !ifid_sRST1)

	.dataa(gnd),
	.datab(gnd),
	.datac(pcifrtnaddr_23),
	.datad(ifid_sRST),
	.cin(gnd),
	.combout(\rtnaddr_l~8_combout ),
	.cout());
// synopsys translate_off
defparam \rtnaddr_l~8 .lut_mask = 16'h00F0;
defparam \rtnaddr_l~8 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X52_Y31_N28
cycloneive_lcell_comb \rtnaddr_l~9 (
// Equation(s):
// \rtnaddr_l~9_combout  = (pcifrtnaddr_22 & !ifid_sRST1)

	.dataa(gnd),
	.datab(gnd),
	.datac(pcifrtnaddr_22),
	.datad(ifid_sRST),
	.cin(gnd),
	.combout(\rtnaddr_l~9_combout ),
	.cout());
// synopsys translate_off
defparam \rtnaddr_l~9 .lut_mask = 16'h00F0;
defparam \rtnaddr_l~9 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X52_Y30_N14
cycloneive_lcell_comb \rtnaddr_l~10 (
// Equation(s):
// \rtnaddr_l~10_combout  = (!ifid_sRST1 & pcifrtnaddr_21)

	.dataa(ifid_sRST),
	.datab(gnd),
	.datac(gnd),
	.datad(pcifrtnaddr_21),
	.cin(gnd),
	.combout(\rtnaddr_l~10_combout ),
	.cout());
// synopsys translate_off
defparam \rtnaddr_l~10 .lut_mask = 16'h5500;
defparam \rtnaddr_l~10 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X52_Y30_N24
cycloneive_lcell_comb \rtnaddr_l~11 (
// Equation(s):
// \rtnaddr_l~11_combout  = (!ifid_sRST1 & pcifrtnaddr_20)

	.dataa(ifid_sRST),
	.datab(gnd),
	.datac(gnd),
	.datad(pcifrtnaddr_20),
	.cin(gnd),
	.combout(\rtnaddr_l~11_combout ),
	.cout());
// synopsys translate_off
defparam \rtnaddr_l~11 .lut_mask = 16'h5500;
defparam \rtnaddr_l~11 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y31_N26
cycloneive_lcell_comb \rtnaddr_l~12 (
// Equation(s):
// \rtnaddr_l~12_combout  = (!ifid_sRST1 & pcifrtnaddr_19)

	.dataa(gnd),
	.datab(gnd),
	.datac(ifid_sRST),
	.datad(pcifrtnaddr_19),
	.cin(gnd),
	.combout(\rtnaddr_l~12_combout ),
	.cout());
// synopsys translate_off
defparam \rtnaddr_l~12 .lut_mask = 16'h0F00;
defparam \rtnaddr_l~12 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y31_N20
cycloneive_lcell_comb \rtnaddr_l~13 (
// Equation(s):
// \rtnaddr_l~13_combout  = (!ifid_sRST1 & pcifrtnaddr_18)

	.dataa(ifid_sRST),
	.datab(gnd),
	.datac(pcifrtnaddr_18),
	.datad(gnd),
	.cin(gnd),
	.combout(\rtnaddr_l~13_combout ),
	.cout());
// synopsys translate_off
defparam \rtnaddr_l~13 .lut_mask = 16'h5050;
defparam \rtnaddr_l~13 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X52_Y31_N18
cycloneive_lcell_comb \rtnaddr_l~14 (
// Equation(s):
// \rtnaddr_l~14_combout  = (pcifrtnaddr_17 & !ifid_sRST1)

	.dataa(gnd),
	.datab(gnd),
	.datac(pcifrtnaddr_17),
	.datad(ifid_sRST),
	.cin(gnd),
	.combout(\rtnaddr_l~14_combout ),
	.cout());
// synopsys translate_off
defparam \rtnaddr_l~14 .lut_mask = 16'h00F0;
defparam \rtnaddr_l~14 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y31_N30
cycloneive_lcell_comb \rtnaddr_l~15 (
// Equation(s):
// \rtnaddr_l~15_combout  = (!ifid_sRST1 & pcifrtnaddr_16)

	.dataa(gnd),
	.datab(gnd),
	.datac(ifid_sRST),
	.datad(pcifrtnaddr_16),
	.cin(gnd),
	.combout(\rtnaddr_l~15_combout ),
	.cout());
// synopsys translate_off
defparam \rtnaddr_l~15 .lut_mask = 16'h0F00;
defparam \rtnaddr_l~15 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y30_N4
cycloneive_lcell_comb \rtnaddr_l~16 (
// Equation(s):
// \rtnaddr_l~16_combout  = (pcifrtnaddr_15 & !ifid_sRST1)

	.dataa(pcifrtnaddr_15),
	.datab(gnd),
	.datac(ifid_sRST),
	.datad(gnd),
	.cin(gnd),
	.combout(\rtnaddr_l~16_combout ),
	.cout());
// synopsys translate_off
defparam \rtnaddr_l~16 .lut_mask = 16'h0A0A;
defparam \rtnaddr_l~16 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y29_N0
cycloneive_lcell_comb \rtnaddr_l~17 (
// Equation(s):
// \rtnaddr_l~17_combout  = (pcifrtnaddr_14 & !ifid_sRST1)

	.dataa(gnd),
	.datab(gnd),
	.datac(pcifrtnaddr_14),
	.datad(ifid_sRST),
	.cin(gnd),
	.combout(\rtnaddr_l~17_combout ),
	.cout());
// synopsys translate_off
defparam \rtnaddr_l~17 .lut_mask = 16'h00F0;
defparam \rtnaddr_l~17 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y31_N24
cycloneive_lcell_comb \rtnaddr_l~18 (
// Equation(s):
// \rtnaddr_l~18_combout  = (!ifid_sRST1 & pcifrtnaddr_13)

	.dataa(ifid_sRST),
	.datab(gnd),
	.datac(pcifrtnaddr_13),
	.datad(gnd),
	.cin(gnd),
	.combout(\rtnaddr_l~18_combout ),
	.cout());
// synopsys translate_off
defparam \rtnaddr_l~18 .lut_mask = 16'h5050;
defparam \rtnaddr_l~18 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y31_N14
cycloneive_lcell_comb \rtnaddr_l~19 (
// Equation(s):
// \rtnaddr_l~19_combout  = (!ifid_sRST1 & pcifrtnaddr_12)

	.dataa(ifid_sRST),
	.datab(gnd),
	.datac(pcifrtnaddr_12),
	.datad(gnd),
	.cin(gnd),
	.combout(\rtnaddr_l~19_combout ),
	.cout());
// synopsys translate_off
defparam \rtnaddr_l~19 .lut_mask = 16'h5050;
defparam \rtnaddr_l~19 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y31_N12
cycloneive_lcell_comb \rtnaddr_l~20 (
// Equation(s):
// \rtnaddr_l~20_combout  = (!ifid_sRST1 & pcifrtnaddr_11)

	.dataa(gnd),
	.datab(gnd),
	.datac(ifid_sRST),
	.datad(pcifrtnaddr_11),
	.cin(gnd),
	.combout(\rtnaddr_l~20_combout ),
	.cout());
// synopsys translate_off
defparam \rtnaddr_l~20 .lut_mask = 16'h0F00;
defparam \rtnaddr_l~20 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y31_N10
cycloneive_lcell_comb \rtnaddr_l~21 (
// Equation(s):
// \rtnaddr_l~21_combout  = (!ifid_sRST1 & pcifrtnaddr_10)

	.dataa(gnd),
	.datab(gnd),
	.datac(ifid_sRST),
	.datad(pcifrtnaddr_10),
	.cin(gnd),
	.combout(\rtnaddr_l~21_combout ),
	.cout());
// synopsys translate_off
defparam \rtnaddr_l~21 .lut_mask = 16'h0F00;
defparam \rtnaddr_l~21 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y31_N2
cycloneive_lcell_comb \rtnaddr_l~22 (
// Equation(s):
// \rtnaddr_l~22_combout  = (pcifrtnaddr_9 & !ifid_sRST1)

	.dataa(gnd),
	.datab(gnd),
	.datac(pcifrtnaddr_9),
	.datad(ifid_sRST),
	.cin(gnd),
	.combout(\rtnaddr_l~22_combout ),
	.cout());
// synopsys translate_off
defparam \rtnaddr_l~22 .lut_mask = 16'h00F0;
defparam \rtnaddr_l~22 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y31_N20
cycloneive_lcell_comb \rtnaddr_l~23 (
// Equation(s):
// \rtnaddr_l~23_combout  = (pcifrtnaddr_8 & !ifid_sRST1)

	.dataa(gnd),
	.datab(gnd),
	.datac(pcifrtnaddr_8),
	.datad(ifid_sRST),
	.cin(gnd),
	.combout(\rtnaddr_l~23_combout ),
	.cout());
// synopsys translate_off
defparam \rtnaddr_l~23 .lut_mask = 16'h00F0;
defparam \rtnaddr_l~23 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y31_N8
cycloneive_lcell_comb \rtnaddr_l~24 (
// Equation(s):
// \rtnaddr_l~24_combout  = (!ifid_sRST1 & pcifrtnaddr_7)

	.dataa(gnd),
	.datab(gnd),
	.datac(ifid_sRST),
	.datad(pcifrtnaddr_7),
	.cin(gnd),
	.combout(\rtnaddr_l~24_combout ),
	.cout());
// synopsys translate_off
defparam \rtnaddr_l~24 .lut_mask = 16'h0F00;
defparam \rtnaddr_l~24 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y31_N10
cycloneive_lcell_comb \rtnaddr_l~25 (
// Equation(s):
// \rtnaddr_l~25_combout  = (!ifid_sRST1 & pcifrtnaddr_6)

	.dataa(ifid_sRST),
	.datab(gnd),
	.datac(gnd),
	.datad(pcifrtnaddr_6),
	.cin(gnd),
	.combout(\rtnaddr_l~25_combout ),
	.cout());
// synopsys translate_off
defparam \rtnaddr_l~25 .lut_mask = 16'h5500;
defparam \rtnaddr_l~25 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y31_N22
cycloneive_lcell_comb \rtnaddr_l~26 (
// Equation(s):
// \rtnaddr_l~26_combout  = (pcifrtnaddr_5 & !ifid_sRST1)

	.dataa(pcifrtnaddr_5),
	.datab(gnd),
	.datac(ifid_sRST),
	.datad(gnd),
	.cin(gnd),
	.combout(\rtnaddr_l~26_combout ),
	.cout());
// synopsys translate_off
defparam \rtnaddr_l~26 .lut_mask = 16'h0A0A;
defparam \rtnaddr_l~26 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X52_Y30_N22
cycloneive_lcell_comb \rtnaddr_l~27 (
// Equation(s):
// \rtnaddr_l~27_combout  = (pcifrtnaddr_2 & !ifid_sRST1)

	.dataa(gnd),
	.datab(gnd),
	.datac(pcifrtnaddr_2),
	.datad(ifid_sRST),
	.cin(gnd),
	.combout(\rtnaddr_l~27_combout ),
	.cout());
// synopsys translate_off
defparam \rtnaddr_l~27 .lut_mask = 16'h00F0;
defparam \rtnaddr_l~27 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y31_N28
cycloneive_lcell_comb \rtnaddr_l~28 (
// Equation(s):
// \rtnaddr_l~28_combout  = (PCreg_1 & !ifid_sRST1)

	.dataa(gnd),
	.datab(PCreg_1),
	.datac(ifid_sRST),
	.datad(gnd),
	.cin(gnd),
	.combout(\rtnaddr_l~28_combout ),
	.cout());
// synopsys translate_off
defparam \rtnaddr_l~28 .lut_mask = 16'h0C0C;
defparam \rtnaddr_l~28 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y31_N6
cycloneive_lcell_comb \rtnaddr_l~29 (
// Equation(s):
// \rtnaddr_l~29_combout  = (!ifid_sRST1 & PCreg_0)

	.dataa(gnd),
	.datab(gnd),
	.datac(ifid_sRST),
	.datad(PCreg_0),
	.cin(gnd),
	.combout(\rtnaddr_l~29_combout ),
	.cout());
// synopsys translate_off
defparam \rtnaddr_l~29 .lut_mask = 16'h0F00;
defparam \rtnaddr_l~29 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y31_N12
cycloneive_lcell_comb \rtnaddr_l~30 (
// Equation(s):
// \rtnaddr_l~30_combout  = (!ifid_sRST1 & pcifrtnaddr_4)

	.dataa(ifid_sRST),
	.datab(gnd),
	.datac(gnd),
	.datad(pcifrtnaddr_4),
	.cin(gnd),
	.combout(\rtnaddr_l~30_combout ),
	.cout());
// synopsys translate_off
defparam \rtnaddr_l~30 .lut_mask = 16'h5500;
defparam \rtnaddr_l~30 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y31_N22
cycloneive_lcell_comb \rtnaddr_l~31 (
// Equation(s):
// \rtnaddr_l~31_combout  = (!ifid_sRST1 & pcifrtnaddr_3)

	.dataa(ifid_sRST),
	.datab(gnd),
	.datac(gnd),
	.datad(pcifrtnaddr_3),
	.cin(gnd),
	.combout(\rtnaddr_l~31_combout ),
	.cout());
// synopsys translate_off
defparam \rtnaddr_l~31 .lut_mask = 16'h5500;
defparam \rtnaddr_l~31 .sum_lutc_input = "datac";
// synopsys translate_on

endmodule

module pipeline_memwb (
	plif_exmemporto_l_1,
	plif_exmemporto_l_0,
	plif_exmemporto_l_3,
	plif_exmemporto_l_2,
	plif_exmemporto_l_5,
	plif_exmemporto_l_4,
	plif_exmemporto_l_7,
	plif_exmemporto_l_6,
	plif_exmemporto_l_9,
	plif_exmemporto_l_8,
	plif_exmemporto_l_11,
	plif_exmemporto_l_10,
	plif_exmemporto_l_13,
	plif_exmemporto_l_12,
	plif_exmemporto_l_15,
	plif_exmemporto_l_14,
	plif_exmemporto_l_17,
	plif_exmemporto_l_16,
	plif_exmemporto_l_19,
	plif_exmemporto_l_18,
	plif_exmemporto_l_21,
	plif_exmemporto_l_20,
	plif_exmemporto_l_23,
	plif_exmemporto_l_22,
	plif_exmemporto_l_25,
	plif_exmemporto_l_24,
	plif_exmemporto_l_27,
	plif_exmemporto_l_26,
	plif_exmemporto_l_29,
	plif_exmemporto_l_28,
	plif_exmemporto_l_31,
	plif_exmemporto_l_30,
	ramiframload_0,
	ramiframload_1,
	ramiframload_2,
	ramiframload_3,
	ramiframload_4,
	ramiframload_5,
	ramiframload_6,
	ramiframload_7,
	ramiframload_8,
	ramiframload_9,
	ramiframload_10,
	ramiframload_11,
	ramiframload_12,
	ramiframload_13,
	ramiframload_14,
	ramiframload_15,
	ramiframload_16,
	ramiframload_17,
	ramiframload_18,
	ramiframload_19,
	ramiframload_20,
	ramiframload_21,
	ramiframload_22,
	ramiframload_23,
	ramiframload_24,
	ramiframload_25,
	ramiframload_26,
	ramiframload_27,
	ramiframload_28,
	ramiframload_29,
	ramiframload_30,
	ramiframload_31,
	plif_memwbpcsrc_l_1,
	plif_memwbpcsrc_l_0,
	plif_exmempcsrc_l_1,
	plif_exmempcsrc_l_0,
	plif_exmemregen_l,
	plif_exmemwsel_l_0,
	plif_exmemwsel_l_1,
	plif_exmemwsel_l_4,
	plif_exmemwsel_l_3,
	plif_exmemwsel_l_2,
	plif_memwbdmemload_l_31,
	plif_memwbporto_l_31,
	plif_memwbregsrc_l_0,
	plif_memwbregsrc_l_1,
	plif_memwbrtnaddr_l_31,
	plif_memwbwsel_l_4,
	plif_memwbwsel_l_3,
	plif_memwbwsel_l_0,
	plif_memwbwsel_l_2,
	plif_memwbwsel_l_1,
	plif_memwbregen_l,
	plif_memwbdmemload_l_30,
	plif_memwbporto_l_30,
	plif_memwbrtnaddr_l_30,
	plif_memwbdmemload_l_29,
	plif_memwbporto_l_29,
	plif_memwbrtnaddr_l_29,
	plif_memwbdmemload_l_28,
	plif_memwbporto_l_28,
	plif_memwbrtnaddr_l_28,
	plif_memwbdmemload_l_27,
	plif_memwbporto_l_27,
	plif_memwbrtnaddr_l_27,
	plif_memwbdmemload_l_26,
	plif_memwbporto_l_26,
	plif_memwbrtnaddr_l_26,
	plif_memwbdmemload_l_25,
	plif_memwbporto_l_25,
	plif_memwbrtnaddr_l_25,
	plif_memwbdmemload_l_24,
	plif_memwbporto_l_24,
	plif_memwbrtnaddr_l_24,
	plif_memwbdmemload_l_23,
	plif_memwbporto_l_23,
	plif_memwbrtnaddr_l_23,
	plif_memwbdmemload_l_22,
	plif_memwbporto_l_22,
	plif_memwbrtnaddr_l_22,
	plif_memwbdmemload_l_21,
	plif_memwbporto_l_21,
	plif_memwbrtnaddr_l_21,
	plif_memwbdmemload_l_20,
	plif_memwbporto_l_20,
	plif_memwbrtnaddr_l_20,
	plif_memwbdmemload_l_19,
	plif_memwbporto_l_19,
	plif_memwbrtnaddr_l_19,
	plif_memwbdmemload_l_18,
	plif_memwbporto_l_18,
	plif_memwbrtnaddr_l_18,
	plif_memwbdmemload_l_17,
	plif_memwbporto_l_17,
	plif_memwbrtnaddr_l_17,
	plif_memwbdmemload_l_16,
	plif_memwbporto_l_16,
	plif_memwbrtnaddr_l_16,
	plif_memwbdmemload_l_15,
	plif_memwbporto_l_15,
	plif_memwbrtnaddr_l_15,
	plif_memwbdmemload_l_14,
	plif_memwbporto_l_14,
	plif_memwbrtnaddr_l_14,
	plif_memwbdmemload_l_13,
	plif_memwbporto_l_13,
	plif_memwbrtnaddr_l_13,
	plif_memwbdmemload_l_12,
	plif_memwbporto_l_12,
	plif_memwbrtnaddr_l_12,
	plif_memwbdmemload_l_11,
	plif_memwbporto_l_11,
	plif_memwbrtnaddr_l_11,
	plif_memwbdmemload_l_10,
	plif_memwbporto_l_10,
	plif_memwbrtnaddr_l_10,
	plif_memwbdmemload_l_9,
	plif_memwbporto_l_9,
	plif_memwbrtnaddr_l_9,
	plif_memwbdmemload_l_8,
	plif_memwbporto_l_8,
	plif_memwbrtnaddr_l_8,
	plif_memwbdmemload_l_7,
	plif_memwbporto_l_7,
	plif_memwbrtnaddr_l_7,
	plif_memwbdmemload_l_6,
	plif_memwbporto_l_6,
	plif_memwbrtnaddr_l_6,
	plif_memwbdmemload_l_5,
	plif_memwbporto_l_5,
	plif_memwbrtnaddr_l_5,
	plif_memwbdmemload_l_2,
	plif_memwbporto_l_2,
	plif_memwbrtnaddr_l_2,
	plif_memwbdmemload_l_1,
	plif_memwbporto_l_1,
	plif_memwbrtnaddr_l_1,
	plif_memwbdmemload_l_0,
	plif_memwbporto_l_0,
	plif_memwbrtnaddr_l_0,
	plif_memwbdmemload_l_4,
	plif_memwbporto_l_4,
	plif_memwbrtnaddr_l_4,
	plif_memwbdmemload_l_3,
	plif_memwbporto_l_3,
	plif_memwbrtnaddr_l_3,
	plif_memwbbtype_l,
	plif_memwbzero_l,
	plif_memwbjaddr_l_1,
	plif_memwbextimm_l_1,
	plif_memwbextimm_l_0,
	plif_memwbjaddr_l_0,
	plif_memwbjaddr_l_3,
	plif_memwbextimm_l_3,
	plif_memwbextimm_l_2,
	plif_memwbjaddr_l_2,
	plif_memwbjaddr_l_5,
	plif_memwbextimm_l_5,
	plif_memwbextimm_l_4,
	plif_memwbjaddr_l_4,
	plif_memwbjaddr_l_7,
	plif_memwbextimm_l_7,
	plif_memwbextimm_l_6,
	plif_memwbjaddr_l_6,
	plif_memwbjaddr_l_9,
	plif_memwbextimm_l_9,
	plif_memwbextimm_l_8,
	plif_memwbjaddr_l_8,
	plif_memwbjaddr_l_11,
	plif_memwbextimm_l_11,
	plif_memwbextimm_l_10,
	plif_memwbjaddr_l_10,
	plif_memwbjaddr_l_13,
	plif_memwbextimm_l_13,
	plif_memwbextimm_l_12,
	plif_memwbjaddr_l_12,
	plif_memwbjaddr_l_15,
	plif_memwbextimm_l_15,
	plif_memwbextimm_l_14,
	plif_memwbjaddr_l_14,
	plif_memwbjaddr_l_17,
	plif_memwbextimm_l_17,
	plif_memwbextimm_l_16,
	plif_memwbjaddr_l_16,
	plif_memwbjaddr_l_19,
	plif_memwbextimm_l_19,
	plif_memwbextimm_l_18,
	plif_memwbjaddr_l_18,
	plif_memwbjaddr_l_21,
	plif_memwbextimm_l_21,
	plif_memwbextimm_l_20,
	plif_memwbjaddr_l_20,
	plif_memwbjaddr_l_23,
	plif_memwbextimm_l_23,
	plif_memwbextimm_l_22,
	plif_memwbjaddr_l_22,
	plif_memwbjaddr_l_25,
	plif_memwbextimm_l_25,
	plif_memwbextimm_l_24,
	plif_memwbjaddr_l_24,
	plif_memwbextimm_l_27,
	plif_memwbextimm_l_26,
	plif_memwbextimm_l_29,
	plif_memwbextimm_l_28,
	plif_exmemregsrc_l_0,
	plif_exmemregsrc_l_1,
	plif_exmemrtnaddr_l_31,
	plif_exmemrtnaddr_l_30,
	plif_exmemrtnaddr_l_29,
	plif_exmemrtnaddr_l_28,
	plif_exmemrtnaddr_l_27,
	plif_exmemrtnaddr_l_26,
	plif_exmemrtnaddr_l_25,
	plif_exmemrtnaddr_l_24,
	plif_exmemrtnaddr_l_23,
	plif_exmemrtnaddr_l_22,
	plif_exmemrtnaddr_l_21,
	plif_exmemrtnaddr_l_20,
	plif_exmemrtnaddr_l_19,
	plif_exmemrtnaddr_l_18,
	plif_exmemrtnaddr_l_17,
	plif_exmemrtnaddr_l_16,
	plif_exmemrtnaddr_l_15,
	plif_exmemrtnaddr_l_14,
	plif_exmemrtnaddr_l_13,
	plif_exmemrtnaddr_l_12,
	plif_exmemrtnaddr_l_11,
	plif_exmemrtnaddr_l_10,
	plif_exmemrtnaddr_l_9,
	plif_exmemrtnaddr_l_8,
	plif_exmemrtnaddr_l_7,
	plif_exmemrtnaddr_l_6,
	plif_exmemrtnaddr_l_5,
	plif_exmemrtnaddr_l_2,
	plif_exmemrtnaddr_l_1,
	plif_exmemrtnaddr_l_0,
	plif_exmemrtnaddr_l_4,
	plif_exmemrtnaddr_l_3,
	plif_exmembtype_l,
	plif_exmemzero_l,
	plif_exmemjaddr_l_1,
	plif_exmemextimm_l_1,
	plif_exmemextimm_l_0,
	plif_exmemjaddr_l_0,
	plif_exmemjaddr_l_3,
	plif_exmemextimm_l_3,
	plif_exmemextimm_l_2,
	plif_exmemjaddr_l_2,
	plif_exmemjaddr_l_5,
	plif_exmemextimm_l_5,
	plif_exmemextimm_l_4,
	plif_exmemjaddr_l_4,
	plif_exmemjaddr_l_7,
	plif_exmemextimm_l_7,
	plif_exmemextimm_l_6,
	plif_exmemjaddr_l_6,
	plif_exmemjaddr_l_9,
	plif_exmemextimm_l_9,
	plif_exmemextimm_l_8,
	plif_exmemjaddr_l_8,
	plif_exmemjaddr_l_11,
	plif_exmemextimm_l_11,
	plif_exmemextimm_l_10,
	plif_exmemjaddr_l_10,
	plif_exmemjaddr_l_13,
	plif_exmemextimm_l_13,
	plif_exmemextimm_l_12,
	plif_exmemjaddr_l_12,
	plif_exmemjaddr_l_15,
	plif_exmemextimm_l_15,
	plif_exmemextimm_l_14,
	plif_exmemjaddr_l_14,
	plif_exmemjaddr_l_17,
	plif_exmemextimm_l_17,
	plif_exmemextimm_l_16,
	plif_exmemjaddr_l_16,
	plif_exmemjaddr_l_19,
	plif_exmemextimm_l_19,
	plif_exmemextimm_l_18,
	plif_exmemjaddr_l_18,
	plif_exmemjaddr_l_21,
	plif_exmemextimm_l_21,
	plif_exmemextimm_l_20,
	plif_exmemjaddr_l_20,
	plif_exmemjaddr_l_23,
	plif_exmemextimm_l_23,
	plif_exmemextimm_l_22,
	plif_exmemjaddr_l_22,
	plif_exmemjaddr_l_25,
	plif_exmemextimm_l_25,
	plif_exmemextimm_l_24,
	plif_exmemjaddr_l_24,
	plif_exmemextimm_l_27,
	plif_exmemextimm_l_26,
	plif_exmemextimm_l_29,
	plif_exmemextimm_l_28,
	CPUCLK,
	nRST,
	devpor,
	devclrn,
	devoe);
input 	plif_exmemporto_l_1;
input 	plif_exmemporto_l_0;
input 	plif_exmemporto_l_3;
input 	plif_exmemporto_l_2;
input 	plif_exmemporto_l_5;
input 	plif_exmemporto_l_4;
input 	plif_exmemporto_l_7;
input 	plif_exmemporto_l_6;
input 	plif_exmemporto_l_9;
input 	plif_exmemporto_l_8;
input 	plif_exmemporto_l_11;
input 	plif_exmemporto_l_10;
input 	plif_exmemporto_l_13;
input 	plif_exmemporto_l_12;
input 	plif_exmemporto_l_15;
input 	plif_exmemporto_l_14;
input 	plif_exmemporto_l_17;
input 	plif_exmemporto_l_16;
input 	plif_exmemporto_l_19;
input 	plif_exmemporto_l_18;
input 	plif_exmemporto_l_21;
input 	plif_exmemporto_l_20;
input 	plif_exmemporto_l_23;
input 	plif_exmemporto_l_22;
input 	plif_exmemporto_l_25;
input 	plif_exmemporto_l_24;
input 	plif_exmemporto_l_27;
input 	plif_exmemporto_l_26;
input 	plif_exmemporto_l_29;
input 	plif_exmemporto_l_28;
input 	plif_exmemporto_l_31;
input 	plif_exmemporto_l_30;
input 	ramiframload_0;
input 	ramiframload_1;
input 	ramiframload_2;
input 	ramiframload_3;
input 	ramiframload_4;
input 	ramiframload_5;
input 	ramiframload_6;
input 	ramiframload_7;
input 	ramiframload_8;
input 	ramiframload_9;
input 	ramiframload_10;
input 	ramiframload_11;
input 	ramiframload_12;
input 	ramiframload_13;
input 	ramiframload_14;
input 	ramiframload_15;
input 	ramiframload_16;
input 	ramiframload_17;
input 	ramiframload_18;
input 	ramiframload_19;
input 	ramiframload_20;
input 	ramiframload_21;
input 	ramiframload_22;
input 	ramiframload_23;
input 	ramiframload_24;
input 	ramiframload_25;
input 	ramiframload_26;
input 	ramiframload_27;
input 	ramiframload_28;
input 	ramiframload_29;
input 	ramiframload_30;
input 	ramiframload_31;
output 	plif_memwbpcsrc_l_1;
output 	plif_memwbpcsrc_l_0;
input 	plif_exmempcsrc_l_1;
input 	plif_exmempcsrc_l_0;
input 	plif_exmemregen_l;
input 	plif_exmemwsel_l_0;
input 	plif_exmemwsel_l_1;
input 	plif_exmemwsel_l_4;
input 	plif_exmemwsel_l_3;
input 	plif_exmemwsel_l_2;
output 	plif_memwbdmemload_l_31;
output 	plif_memwbporto_l_31;
output 	plif_memwbregsrc_l_0;
output 	plif_memwbregsrc_l_1;
output 	plif_memwbrtnaddr_l_31;
output 	plif_memwbwsel_l_4;
output 	plif_memwbwsel_l_3;
output 	plif_memwbwsel_l_0;
output 	plif_memwbwsel_l_2;
output 	plif_memwbwsel_l_1;
output 	plif_memwbregen_l;
output 	plif_memwbdmemload_l_30;
output 	plif_memwbporto_l_30;
output 	plif_memwbrtnaddr_l_30;
output 	plif_memwbdmemload_l_29;
output 	plif_memwbporto_l_29;
output 	plif_memwbrtnaddr_l_29;
output 	plif_memwbdmemload_l_28;
output 	plif_memwbporto_l_28;
output 	plif_memwbrtnaddr_l_28;
output 	plif_memwbdmemload_l_27;
output 	plif_memwbporto_l_27;
output 	plif_memwbrtnaddr_l_27;
output 	plif_memwbdmemload_l_26;
output 	plif_memwbporto_l_26;
output 	plif_memwbrtnaddr_l_26;
output 	plif_memwbdmemload_l_25;
output 	plif_memwbporto_l_25;
output 	plif_memwbrtnaddr_l_25;
output 	plif_memwbdmemload_l_24;
output 	plif_memwbporto_l_24;
output 	plif_memwbrtnaddr_l_24;
output 	plif_memwbdmemload_l_23;
output 	plif_memwbporto_l_23;
output 	plif_memwbrtnaddr_l_23;
output 	plif_memwbdmemload_l_22;
output 	plif_memwbporto_l_22;
output 	plif_memwbrtnaddr_l_22;
output 	plif_memwbdmemload_l_21;
output 	plif_memwbporto_l_21;
output 	plif_memwbrtnaddr_l_21;
output 	plif_memwbdmemload_l_20;
output 	plif_memwbporto_l_20;
output 	plif_memwbrtnaddr_l_20;
output 	plif_memwbdmemload_l_19;
output 	plif_memwbporto_l_19;
output 	plif_memwbrtnaddr_l_19;
output 	plif_memwbdmemload_l_18;
output 	plif_memwbporto_l_18;
output 	plif_memwbrtnaddr_l_18;
output 	plif_memwbdmemload_l_17;
output 	plif_memwbporto_l_17;
output 	plif_memwbrtnaddr_l_17;
output 	plif_memwbdmemload_l_16;
output 	plif_memwbporto_l_16;
output 	plif_memwbrtnaddr_l_16;
output 	plif_memwbdmemload_l_15;
output 	plif_memwbporto_l_15;
output 	plif_memwbrtnaddr_l_15;
output 	plif_memwbdmemload_l_14;
output 	plif_memwbporto_l_14;
output 	plif_memwbrtnaddr_l_14;
output 	plif_memwbdmemload_l_13;
output 	plif_memwbporto_l_13;
output 	plif_memwbrtnaddr_l_13;
output 	plif_memwbdmemload_l_12;
output 	plif_memwbporto_l_12;
output 	plif_memwbrtnaddr_l_12;
output 	plif_memwbdmemload_l_11;
output 	plif_memwbporto_l_11;
output 	plif_memwbrtnaddr_l_11;
output 	plif_memwbdmemload_l_10;
output 	plif_memwbporto_l_10;
output 	plif_memwbrtnaddr_l_10;
output 	plif_memwbdmemload_l_9;
output 	plif_memwbporto_l_9;
output 	plif_memwbrtnaddr_l_9;
output 	plif_memwbdmemload_l_8;
output 	plif_memwbporto_l_8;
output 	plif_memwbrtnaddr_l_8;
output 	plif_memwbdmemload_l_7;
output 	plif_memwbporto_l_7;
output 	plif_memwbrtnaddr_l_7;
output 	plif_memwbdmemload_l_6;
output 	plif_memwbporto_l_6;
output 	plif_memwbrtnaddr_l_6;
output 	plif_memwbdmemload_l_5;
output 	plif_memwbporto_l_5;
output 	plif_memwbrtnaddr_l_5;
output 	plif_memwbdmemload_l_2;
output 	plif_memwbporto_l_2;
output 	plif_memwbrtnaddr_l_2;
output 	plif_memwbdmemload_l_1;
output 	plif_memwbporto_l_1;
output 	plif_memwbrtnaddr_l_1;
output 	plif_memwbdmemload_l_0;
output 	plif_memwbporto_l_0;
output 	plif_memwbrtnaddr_l_0;
output 	plif_memwbdmemload_l_4;
output 	plif_memwbporto_l_4;
output 	plif_memwbrtnaddr_l_4;
output 	plif_memwbdmemload_l_3;
output 	plif_memwbporto_l_3;
output 	plif_memwbrtnaddr_l_3;
output 	plif_memwbbtype_l;
output 	plif_memwbzero_l;
output 	plif_memwbjaddr_l_1;
output 	plif_memwbextimm_l_1;
output 	plif_memwbextimm_l_0;
output 	plif_memwbjaddr_l_0;
output 	plif_memwbjaddr_l_3;
output 	plif_memwbextimm_l_3;
output 	plif_memwbextimm_l_2;
output 	plif_memwbjaddr_l_2;
output 	plif_memwbjaddr_l_5;
output 	plif_memwbextimm_l_5;
output 	plif_memwbextimm_l_4;
output 	plif_memwbjaddr_l_4;
output 	plif_memwbjaddr_l_7;
output 	plif_memwbextimm_l_7;
output 	plif_memwbextimm_l_6;
output 	plif_memwbjaddr_l_6;
output 	plif_memwbjaddr_l_9;
output 	plif_memwbextimm_l_9;
output 	plif_memwbextimm_l_8;
output 	plif_memwbjaddr_l_8;
output 	plif_memwbjaddr_l_11;
output 	plif_memwbextimm_l_11;
output 	plif_memwbextimm_l_10;
output 	plif_memwbjaddr_l_10;
output 	plif_memwbjaddr_l_13;
output 	plif_memwbextimm_l_13;
output 	plif_memwbextimm_l_12;
output 	plif_memwbjaddr_l_12;
output 	plif_memwbjaddr_l_15;
output 	plif_memwbextimm_l_15;
output 	plif_memwbextimm_l_14;
output 	plif_memwbjaddr_l_14;
output 	plif_memwbjaddr_l_17;
output 	plif_memwbextimm_l_17;
output 	plif_memwbextimm_l_16;
output 	plif_memwbjaddr_l_16;
output 	plif_memwbjaddr_l_19;
output 	plif_memwbextimm_l_19;
output 	plif_memwbextimm_l_18;
output 	plif_memwbjaddr_l_18;
output 	plif_memwbjaddr_l_21;
output 	plif_memwbextimm_l_21;
output 	plif_memwbextimm_l_20;
output 	plif_memwbjaddr_l_20;
output 	plif_memwbjaddr_l_23;
output 	plif_memwbextimm_l_23;
output 	plif_memwbextimm_l_22;
output 	plif_memwbjaddr_l_22;
output 	plif_memwbjaddr_l_25;
output 	plif_memwbextimm_l_25;
output 	plif_memwbextimm_l_24;
output 	plif_memwbjaddr_l_24;
output 	plif_memwbextimm_l_27;
output 	plif_memwbextimm_l_26;
output 	plif_memwbextimm_l_29;
output 	plif_memwbextimm_l_28;
input 	plif_exmemregsrc_l_0;
input 	plif_exmemregsrc_l_1;
input 	plif_exmemrtnaddr_l_31;
input 	plif_exmemrtnaddr_l_30;
input 	plif_exmemrtnaddr_l_29;
input 	plif_exmemrtnaddr_l_28;
input 	plif_exmemrtnaddr_l_27;
input 	plif_exmemrtnaddr_l_26;
input 	plif_exmemrtnaddr_l_25;
input 	plif_exmemrtnaddr_l_24;
input 	plif_exmemrtnaddr_l_23;
input 	plif_exmemrtnaddr_l_22;
input 	plif_exmemrtnaddr_l_21;
input 	plif_exmemrtnaddr_l_20;
input 	plif_exmemrtnaddr_l_19;
input 	plif_exmemrtnaddr_l_18;
input 	plif_exmemrtnaddr_l_17;
input 	plif_exmemrtnaddr_l_16;
input 	plif_exmemrtnaddr_l_15;
input 	plif_exmemrtnaddr_l_14;
input 	plif_exmemrtnaddr_l_13;
input 	plif_exmemrtnaddr_l_12;
input 	plif_exmemrtnaddr_l_11;
input 	plif_exmemrtnaddr_l_10;
input 	plif_exmemrtnaddr_l_9;
input 	plif_exmemrtnaddr_l_8;
input 	plif_exmemrtnaddr_l_7;
input 	plif_exmemrtnaddr_l_6;
input 	plif_exmemrtnaddr_l_5;
input 	plif_exmemrtnaddr_l_2;
input 	plif_exmemrtnaddr_l_1;
input 	plif_exmemrtnaddr_l_0;
input 	plif_exmemrtnaddr_l_4;
input 	plif_exmemrtnaddr_l_3;
input 	plif_exmembtype_l;
input 	plif_exmemzero_l;
input 	plif_exmemjaddr_l_1;
input 	plif_exmemextimm_l_1;
input 	plif_exmemextimm_l_0;
input 	plif_exmemjaddr_l_0;
input 	plif_exmemjaddr_l_3;
input 	plif_exmemextimm_l_3;
input 	plif_exmemextimm_l_2;
input 	plif_exmemjaddr_l_2;
input 	plif_exmemjaddr_l_5;
input 	plif_exmemextimm_l_5;
input 	plif_exmemextimm_l_4;
input 	plif_exmemjaddr_l_4;
input 	plif_exmemjaddr_l_7;
input 	plif_exmemextimm_l_7;
input 	plif_exmemextimm_l_6;
input 	plif_exmemjaddr_l_6;
input 	plif_exmemjaddr_l_9;
input 	plif_exmemextimm_l_9;
input 	plif_exmemextimm_l_8;
input 	plif_exmemjaddr_l_8;
input 	plif_exmemjaddr_l_11;
input 	plif_exmemextimm_l_11;
input 	plif_exmemextimm_l_10;
input 	plif_exmemjaddr_l_10;
input 	plif_exmemjaddr_l_13;
input 	plif_exmemextimm_l_13;
input 	plif_exmemextimm_l_12;
input 	plif_exmemjaddr_l_12;
input 	plif_exmemjaddr_l_15;
input 	plif_exmemextimm_l_15;
input 	plif_exmemextimm_l_14;
input 	plif_exmemjaddr_l_14;
input 	plif_exmemjaddr_l_17;
input 	plif_exmemextimm_l_17;
input 	plif_exmemextimm_l_16;
input 	plif_exmemjaddr_l_16;
input 	plif_exmemjaddr_l_19;
input 	plif_exmemextimm_l_19;
input 	plif_exmemextimm_l_18;
input 	plif_exmemjaddr_l_18;
input 	plif_exmemjaddr_l_21;
input 	plif_exmemextimm_l_21;
input 	plif_exmemextimm_l_20;
input 	plif_exmemjaddr_l_20;
input 	plif_exmemjaddr_l_23;
input 	plif_exmemextimm_l_23;
input 	plif_exmemextimm_l_22;
input 	plif_exmemjaddr_l_22;
input 	plif_exmemjaddr_l_25;
input 	plif_exmemextimm_l_25;
input 	plif_exmemextimm_l_24;
input 	plif_exmemjaddr_l_24;
input 	plif_exmemextimm_l_27;
input 	plif_exmemextimm_l_26;
input 	plif_exmemextimm_l_29;
input 	plif_exmemextimm_l_28;
input 	CPUCLK;
input 	nRST;

// Design Ports Information

input 	devpor;
input 	devclrn;
input 	devoe;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
assign unknown = 1'bx;

wire \plif_memwb.regsrc_l[0]~feeder_combout ;
wire \plif_memwb.regsrc_l[1]~feeder_combout ;
wire \plif_memwb.porto_l[29]~feeder_combout ;
wire \plif_memwb.porto_l[28]~feeder_combout ;
wire \plif_memwb.rtnaddr_l[28]~feeder_combout ;
wire \plif_memwb.porto_l[27]~feeder_combout ;
wire \plif_memwb.porto_l[24]~feeder_combout ;
wire \plif_memwb.porto_l[23]~feeder_combout ;
wire \plif_memwb.rtnaddr_l[23]~feeder_combout ;
wire \plif_memwb.rtnaddr_l[22]~feeder_combout ;
wire \plif_memwb.porto_l[21]~feeder_combout ;
wire \plif_memwb.porto_l[19]~feeder_combout ;
wire \plif_memwb.rtnaddr_l[16]~feeder_combout ;
wire \plif_memwb.porto_l[10]~feeder_combout ;
wire \plif_memwb.porto_l[9]~feeder_combout ;
wire \plif_memwb.rtnaddr_l[9]~feeder_combout ;
wire \plif_memwb.porto_l[8]~feeder_combout ;
wire \plif_memwb.rtnaddr_l[2]~feeder_combout ;
wire \plif_memwb.porto_l[1]~feeder_combout ;
wire \plif_memwb.rtnaddr_l[1]~feeder_combout ;
wire \plif_memwb.porto_l[0]~feeder_combout ;
wire \plif_memwb.rtnaddr_l[0]~feeder_combout ;
wire \plif_memwb.porto_l[4]~feeder_combout ;
wire \plif_memwb.rtnaddr_l[4]~feeder_combout ;
wire \plif_memwb.porto_l[3]~feeder_combout ;
wire \plif_memwb.rtnaddr_l[3]~feeder_combout ;
wire \plif_memwb.btype_l~feeder_combout ;
wire \plif_memwb.jaddr_l[1]~feeder_combout ;
wire \plif_memwb.extimm_l[0]~feeder_combout ;
wire \plif_memwb.jaddr_l[5]~feeder_combout ;
wire \plif_memwb.extimm_l[7]~feeder_combout ;
wire \plif_memwb.jaddr_l[9]~feeder_combout ;
wire \plif_memwb.extimm_l[8]~feeder_combout ;
wire \plif_memwb.jaddr_l[11]~feeder_combout ;
wire \plif_memwb.extimm_l[11]~feeder_combout ;
wire \plif_memwb.extimm_l[12]~feeder_combout ;
wire \plif_memwb.jaddr_l[15]~feeder_combout ;
wire \plif_memwb.extimm_l[15]~feeder_combout ;
wire \plif_memwb.extimm_l[14]~feeder_combout ;
wire \plif_memwb.jaddr_l[17]~feeder_combout ;
wire \plif_memwb.extimm_l[17]~feeder_combout ;
wire \plif_memwb.jaddr_l[19]~feeder_combout ;
wire \plif_memwb.extimm_l[18]~feeder_combout ;
wire \plif_memwb.jaddr_l[21]~feeder_combout ;
wire \plif_memwb.extimm_l[23]~feeder_combout ;
wire \plif_memwb.jaddr_l[25]~feeder_combout ;
wire \plif_memwb.extimm_l[24]~feeder_combout ;
wire \plif_memwb.extimm_l[28]~feeder_combout ;


// Location: FF_X55_Y32_N25
dffeas \plif_memwb.pcsrc_l[1] (
	.clk(CPUCLK),
	.d(gnd),
	.asdata(plif_exmempcsrc_l_1),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(plif_memwbpcsrc_l_1),
	.prn(vcc));
// synopsys translate_off
defparam \plif_memwb.pcsrc_l[1] .is_wysiwyg = "true";
defparam \plif_memwb.pcsrc_l[1] .power_up = "low";
// synopsys translate_on

// Location: FF_X55_Y32_N7
dffeas \plif_memwb.pcsrc_l[0] (
	.clk(CPUCLK),
	.d(gnd),
	.asdata(plif_exmempcsrc_l_0),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(plif_memwbpcsrc_l_0),
	.prn(vcc));
// synopsys translate_off
defparam \plif_memwb.pcsrc_l[0] .is_wysiwyg = "true";
defparam \plif_memwb.pcsrc_l[0] .power_up = "low";
// synopsys translate_on

// Location: FF_X55_Y41_N1
dffeas \plif_memwb.dmemload_l[31] (
	.clk(CPUCLK),
	.d(gnd),
	.asdata(ramiframload_31),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(plif_memwbdmemload_l_31),
	.prn(vcc));
// synopsys translate_off
defparam \plif_memwb.dmemload_l[31] .is_wysiwyg = "true";
defparam \plif_memwb.dmemload_l[31] .power_up = "low";
// synopsys translate_on

// Location: FF_X55_Y41_N3
dffeas \plif_memwb.porto_l[31] (
	.clk(CPUCLK),
	.d(gnd),
	.asdata(plif_exmemporto_l_31),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(plif_memwbporto_l_31),
	.prn(vcc));
// synopsys translate_off
defparam \plif_memwb.porto_l[31] .is_wysiwyg = "true";
defparam \plif_memwb.porto_l[31] .power_up = "low";
// synopsys translate_on

// Location: FF_X56_Y35_N5
dffeas \plif_memwb.regsrc_l[0] (
	.clk(CPUCLK),
	.d(\plif_memwb.regsrc_l[0]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(plif_memwbregsrc_l_0),
	.prn(vcc));
// synopsys translate_off
defparam \plif_memwb.regsrc_l[0] .is_wysiwyg = "true";
defparam \plif_memwb.regsrc_l[0] .power_up = "low";
// synopsys translate_on

// Location: FF_X56_Y35_N31
dffeas \plif_memwb.regsrc_l[1] (
	.clk(CPUCLK),
	.d(\plif_memwb.regsrc_l[1]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(plif_memwbregsrc_l_1),
	.prn(vcc));
// synopsys translate_off
defparam \plif_memwb.regsrc_l[1] .is_wysiwyg = "true";
defparam \plif_memwb.regsrc_l[1] .power_up = "low";
// synopsys translate_on

// Location: FF_X55_Y41_N9
dffeas \plif_memwb.rtnaddr_l[31] (
	.clk(CPUCLK),
	.d(gnd),
	.asdata(plif_exmemrtnaddr_l_31),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(plif_memwbrtnaddr_l_31),
	.prn(vcc));
// synopsys translate_off
defparam \plif_memwb.rtnaddr_l[31] .is_wysiwyg = "true";
defparam \plif_memwb.rtnaddr_l[31] .power_up = "low";
// synopsys translate_on

// Location: FF_X57_Y37_N29
dffeas \plif_memwb.wsel_l[4] (
	.clk(CPUCLK),
	.d(gnd),
	.asdata(plif_exmemwsel_l_4),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(plif_memwbwsel_l_4),
	.prn(vcc));
// synopsys translate_off
defparam \plif_memwb.wsel_l[4] .is_wysiwyg = "true";
defparam \plif_memwb.wsel_l[4] .power_up = "low";
// synopsys translate_on

// Location: FF_X57_Y37_N5
dffeas \plif_memwb.wsel_l[3] (
	.clk(CPUCLK),
	.d(gnd),
	.asdata(plif_exmemwsel_l_3),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(plif_memwbwsel_l_3),
	.prn(vcc));
// synopsys translate_off
defparam \plif_memwb.wsel_l[3] .is_wysiwyg = "true";
defparam \plif_memwb.wsel_l[3] .power_up = "low";
// synopsys translate_on

// Location: FF_X57_Y37_N9
dffeas \plif_memwb.wsel_l[0] (
	.clk(CPUCLK),
	.d(gnd),
	.asdata(plif_exmemwsel_l_0),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(plif_memwbwsel_l_0),
	.prn(vcc));
// synopsys translate_off
defparam \plif_memwb.wsel_l[0] .is_wysiwyg = "true";
defparam \plif_memwb.wsel_l[0] .power_up = "low";
// synopsys translate_on

// Location: FF_X58_Y37_N31
dffeas \plif_memwb.wsel_l[2] (
	.clk(CPUCLK),
	.d(gnd),
	.asdata(plif_exmemwsel_l_2),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(plif_memwbwsel_l_2),
	.prn(vcc));
// synopsys translate_off
defparam \plif_memwb.wsel_l[2] .is_wysiwyg = "true";
defparam \plif_memwb.wsel_l[2] .power_up = "low";
// synopsys translate_on

// Location: FF_X58_Y37_N13
dffeas \plif_memwb.wsel_l[1] (
	.clk(CPUCLK),
	.d(gnd),
	.asdata(plif_exmemwsel_l_1),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(plif_memwbwsel_l_1),
	.prn(vcc));
// synopsys translate_off
defparam \plif_memwb.wsel_l[1] .is_wysiwyg = "true";
defparam \plif_memwb.wsel_l[1] .power_up = "low";
// synopsys translate_on

// Location: FF_X57_Y37_N25
dffeas \plif_memwb.regen_l (
	.clk(CPUCLK),
	.d(gnd),
	.asdata(plif_exmemregen_l),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(plif_memwbregen_l),
	.prn(vcc));
// synopsys translate_off
defparam \plif_memwb.regen_l .is_wysiwyg = "true";
defparam \plif_memwb.regen_l .power_up = "low";
// synopsys translate_on

// Location: FF_X55_Y42_N11
dffeas \plif_memwb.dmemload_l[30] (
	.clk(CPUCLK),
	.d(gnd),
	.asdata(ramiframload_30),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(plif_memwbdmemload_l_30),
	.prn(vcc));
// synopsys translate_off
defparam \plif_memwb.dmemload_l[30] .is_wysiwyg = "true";
defparam \plif_memwb.dmemload_l[30] .power_up = "low";
// synopsys translate_on

// Location: FF_X55_Y42_N3
dffeas \plif_memwb.porto_l[30] (
	.clk(CPUCLK),
	.d(gnd),
	.asdata(plif_exmemporto_l_30),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(plif_memwbporto_l_30),
	.prn(vcc));
// synopsys translate_off
defparam \plif_memwb.porto_l[30] .is_wysiwyg = "true";
defparam \plif_memwb.porto_l[30] .power_up = "low";
// synopsys translate_on

// Location: FF_X55_Y42_N17
dffeas \plif_memwb.rtnaddr_l[30] (
	.clk(CPUCLK),
	.d(gnd),
	.asdata(plif_exmemrtnaddr_l_30),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(plif_memwbrtnaddr_l_30),
	.prn(vcc));
// synopsys translate_off
defparam \plif_memwb.rtnaddr_l[30] .is_wysiwyg = "true";
defparam \plif_memwb.rtnaddr_l[30] .power_up = "low";
// synopsys translate_on

// Location: FF_X56_Y35_N29
dffeas \plif_memwb.dmemload_l[29] (
	.clk(CPUCLK),
	.d(gnd),
	.asdata(ramiframload_29),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(plif_memwbdmemload_l_29),
	.prn(vcc));
// synopsys translate_off
defparam \plif_memwb.dmemload_l[29] .is_wysiwyg = "true";
defparam \plif_memwb.dmemload_l[29] .power_up = "low";
// synopsys translate_on

// Location: FF_X55_Y35_N29
dffeas \plif_memwb.porto_l[29] (
	.clk(CPUCLK),
	.d(\plif_memwb.porto_l[29]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(plif_memwbporto_l_29),
	.prn(vcc));
// synopsys translate_off
defparam \plif_memwb.porto_l[29] .is_wysiwyg = "true";
defparam \plif_memwb.porto_l[29] .power_up = "low";
// synopsys translate_on

// Location: FF_X56_Y35_N15
dffeas \plif_memwb.rtnaddr_l[29] (
	.clk(CPUCLK),
	.d(gnd),
	.asdata(plif_exmemrtnaddr_l_29),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(plif_memwbrtnaddr_l_29),
	.prn(vcc));
// synopsys translate_off
defparam \plif_memwb.rtnaddr_l[29] .is_wysiwyg = "true";
defparam \plif_memwb.rtnaddr_l[29] .power_up = "low";
// synopsys translate_on

// Location: FF_X57_Y35_N21
dffeas \plif_memwb.dmemload_l[28] (
	.clk(CPUCLK),
	.d(gnd),
	.asdata(ramiframload_28),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(plif_memwbdmemload_l_28),
	.prn(vcc));
// synopsys translate_off
defparam \plif_memwb.dmemload_l[28] .is_wysiwyg = "true";
defparam \plif_memwb.dmemload_l[28] .power_up = "low";
// synopsys translate_on

// Location: FF_X57_Y35_N19
dffeas \plif_memwb.porto_l[28] (
	.clk(CPUCLK),
	.d(\plif_memwb.porto_l[28]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(plif_memwbporto_l_28),
	.prn(vcc));
// synopsys translate_off
defparam \plif_memwb.porto_l[28] .is_wysiwyg = "true";
defparam \plif_memwb.porto_l[28] .power_up = "low";
// synopsys translate_on

// Location: FF_X57_Y35_N17
dffeas \plif_memwb.rtnaddr_l[28] (
	.clk(CPUCLK),
	.d(\plif_memwb.rtnaddr_l[28]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(plif_memwbrtnaddr_l_28),
	.prn(vcc));
// synopsys translate_off
defparam \plif_memwb.rtnaddr_l[28] .is_wysiwyg = "true";
defparam \plif_memwb.rtnaddr_l[28] .power_up = "low";
// synopsys translate_on

// Location: FF_X56_Y36_N21
dffeas \plif_memwb.dmemload_l[27] (
	.clk(CPUCLK),
	.d(gnd),
	.asdata(ramiframload_27),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(plif_memwbdmemload_l_27),
	.prn(vcc));
// synopsys translate_off
defparam \plif_memwb.dmemload_l[27] .is_wysiwyg = "true";
defparam \plif_memwb.dmemload_l[27] .power_up = "low";
// synopsys translate_on

// Location: FF_X56_Y36_N31
dffeas \plif_memwb.porto_l[27] (
	.clk(CPUCLK),
	.d(\plif_memwb.porto_l[27]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(plif_memwbporto_l_27),
	.prn(vcc));
// synopsys translate_off
defparam \plif_memwb.porto_l[27] .is_wysiwyg = "true";
defparam \plif_memwb.porto_l[27] .power_up = "low";
// synopsys translate_on

// Location: FF_X57_Y36_N1
dffeas \plif_memwb.rtnaddr_l[27] (
	.clk(CPUCLK),
	.d(gnd),
	.asdata(plif_exmemrtnaddr_l_27),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(plif_memwbrtnaddr_l_27),
	.prn(vcc));
// synopsys translate_off
defparam \plif_memwb.rtnaddr_l[27] .is_wysiwyg = "true";
defparam \plif_memwb.rtnaddr_l[27] .power_up = "low";
// synopsys translate_on

// Location: FF_X56_Y36_N5
dffeas \plif_memwb.dmemload_l[26] (
	.clk(CPUCLK),
	.d(gnd),
	.asdata(ramiframload_26),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(plif_memwbdmemload_l_26),
	.prn(vcc));
// synopsys translate_off
defparam \plif_memwb.dmemload_l[26] .is_wysiwyg = "true";
defparam \plif_memwb.dmemload_l[26] .power_up = "low";
// synopsys translate_on

// Location: FF_X56_Y36_N7
dffeas \plif_memwb.porto_l[26] (
	.clk(CPUCLK),
	.d(gnd),
	.asdata(plif_exmemporto_l_26),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(plif_memwbporto_l_26),
	.prn(vcc));
// synopsys translate_off
defparam \plif_memwb.porto_l[26] .is_wysiwyg = "true";
defparam \plif_memwb.porto_l[26] .power_up = "low";
// synopsys translate_on

// Location: FF_X56_Y36_N9
dffeas \plif_memwb.rtnaddr_l[26] (
	.clk(CPUCLK),
	.d(gnd),
	.asdata(plif_exmemrtnaddr_l_26),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(plif_memwbrtnaddr_l_26),
	.prn(vcc));
// synopsys translate_off
defparam \plif_memwb.rtnaddr_l[26] .is_wysiwyg = "true";
defparam \plif_memwb.rtnaddr_l[26] .power_up = "low";
// synopsys translate_on

// Location: FF_X56_Y36_N15
dffeas \plif_memwb.dmemload_l[25] (
	.clk(CPUCLK),
	.d(gnd),
	.asdata(ramiframload_25),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(plif_memwbdmemload_l_25),
	.prn(vcc));
// synopsys translate_off
defparam \plif_memwb.dmemload_l[25] .is_wysiwyg = "true";
defparam \plif_memwb.dmemload_l[25] .power_up = "low";
// synopsys translate_on

// Location: FF_X56_Y36_N13
dffeas \plif_memwb.porto_l[25] (
	.clk(CPUCLK),
	.d(gnd),
	.asdata(plif_exmemporto_l_25),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(plif_memwbporto_l_25),
	.prn(vcc));
// synopsys translate_off
defparam \plif_memwb.porto_l[25] .is_wysiwyg = "true";
defparam \plif_memwb.porto_l[25] .power_up = "low";
// synopsys translate_on

// Location: FF_X57_Y36_N31
dffeas \plif_memwb.rtnaddr_l[25] (
	.clk(CPUCLK),
	.d(gnd),
	.asdata(plif_exmemrtnaddr_l_25),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(plif_memwbrtnaddr_l_25),
	.prn(vcc));
// synopsys translate_off
defparam \plif_memwb.rtnaddr_l[25] .is_wysiwyg = "true";
defparam \plif_memwb.rtnaddr_l[25] .power_up = "low";
// synopsys translate_on

// Location: FF_X53_Y35_N15
dffeas \plif_memwb.dmemload_l[24] (
	.clk(CPUCLK),
	.d(gnd),
	.asdata(ramiframload_24),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(plif_memwbdmemload_l_24),
	.prn(vcc));
// synopsys translate_off
defparam \plif_memwb.dmemload_l[24] .is_wysiwyg = "true";
defparam \plif_memwb.dmemload_l[24] .power_up = "low";
// synopsys translate_on

// Location: FF_X53_Y35_N29
dffeas \plif_memwb.porto_l[24] (
	.clk(CPUCLK),
	.d(\plif_memwb.porto_l[24]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(plif_memwbporto_l_24),
	.prn(vcc));
// synopsys translate_off
defparam \plif_memwb.porto_l[24] .is_wysiwyg = "true";
defparam \plif_memwb.porto_l[24] .power_up = "low";
// synopsys translate_on

// Location: FF_X53_Y35_N3
dffeas \plif_memwb.rtnaddr_l[24] (
	.clk(CPUCLK),
	.d(gnd),
	.asdata(plif_exmemrtnaddr_l_24),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(plif_memwbrtnaddr_l_24),
	.prn(vcc));
// synopsys translate_off
defparam \plif_memwb.rtnaddr_l[24] .is_wysiwyg = "true";
defparam \plif_memwb.rtnaddr_l[24] .power_up = "low";
// synopsys translate_on

// Location: FF_X56_Y35_N11
dffeas \plif_memwb.dmemload_l[23] (
	.clk(CPUCLK),
	.d(gnd),
	.asdata(ramiframload_23),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(plif_memwbdmemload_l_23),
	.prn(vcc));
// synopsys translate_off
defparam \plif_memwb.dmemload_l[23] .is_wysiwyg = "true";
defparam \plif_memwb.dmemload_l[23] .power_up = "low";
// synopsys translate_on

// Location: FF_X55_Y35_N23
dffeas \plif_memwb.porto_l[23] (
	.clk(CPUCLK),
	.d(\plif_memwb.porto_l[23]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(plif_memwbporto_l_23),
	.prn(vcc));
// synopsys translate_off
defparam \plif_memwb.porto_l[23] .is_wysiwyg = "true";
defparam \plif_memwb.porto_l[23] .power_up = "low";
// synopsys translate_on

// Location: FF_X52_Y39_N9
dffeas \plif_memwb.rtnaddr_l[23] (
	.clk(CPUCLK),
	.d(\plif_memwb.rtnaddr_l[23]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(plif_memwbrtnaddr_l_23),
	.prn(vcc));
// synopsys translate_off
defparam \plif_memwb.rtnaddr_l[23] .is_wysiwyg = "true";
defparam \plif_memwb.rtnaddr_l[23] .power_up = "low";
// synopsys translate_on

// Location: FF_X58_Y39_N5
dffeas \plif_memwb.dmemload_l[22] (
	.clk(CPUCLK),
	.d(gnd),
	.asdata(ramiframload_22),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(plif_memwbdmemload_l_22),
	.prn(vcc));
// synopsys translate_off
defparam \plif_memwb.dmemload_l[22] .is_wysiwyg = "true";
defparam \plif_memwb.dmemload_l[22] .power_up = "low";
// synopsys translate_on

// Location: FF_X58_Y39_N3
dffeas \plif_memwb.porto_l[22] (
	.clk(CPUCLK),
	.d(gnd),
	.asdata(plif_exmemporto_l_22),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(plif_memwbporto_l_22),
	.prn(vcc));
// synopsys translate_off
defparam \plif_memwb.porto_l[22] .is_wysiwyg = "true";
defparam \plif_memwb.porto_l[22] .power_up = "low";
// synopsys translate_on

// Location: FF_X58_Y39_N9
dffeas \plif_memwb.rtnaddr_l[22] (
	.clk(CPUCLK),
	.d(\plif_memwb.rtnaddr_l[22]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(plif_memwbrtnaddr_l_22),
	.prn(vcc));
// synopsys translate_off
defparam \plif_memwb.rtnaddr_l[22] .is_wysiwyg = "true";
defparam \plif_memwb.rtnaddr_l[22] .power_up = "low";
// synopsys translate_on

// Location: FF_X56_Y35_N21
dffeas \plif_memwb.dmemload_l[21] (
	.clk(CPUCLK),
	.d(gnd),
	.asdata(ramiframload_21),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(plif_memwbdmemload_l_21),
	.prn(vcc));
// synopsys translate_off
defparam \plif_memwb.dmemload_l[21] .is_wysiwyg = "true";
defparam \plif_memwb.dmemload_l[21] .power_up = "low";
// synopsys translate_on

// Location: FF_X56_Y35_N23
dffeas \plif_memwb.porto_l[21] (
	.clk(CPUCLK),
	.d(\plif_memwb.porto_l[21]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(plif_memwbporto_l_21),
	.prn(vcc));
// synopsys translate_off
defparam \plif_memwb.porto_l[21] .is_wysiwyg = "true";
defparam \plif_memwb.porto_l[21] .power_up = "low";
// synopsys translate_on

// Location: FF_X56_Y35_N1
dffeas \plif_memwb.rtnaddr_l[21] (
	.clk(CPUCLK),
	.d(gnd),
	.asdata(plif_exmemrtnaddr_l_21),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(plif_memwbrtnaddr_l_21),
	.prn(vcc));
// synopsys translate_off
defparam \plif_memwb.rtnaddr_l[21] .is_wysiwyg = "true";
defparam \plif_memwb.rtnaddr_l[21] .power_up = "low";
// synopsys translate_on

// Location: FF_X54_Y39_N9
dffeas \plif_memwb.dmemload_l[20] (
	.clk(CPUCLK),
	.d(gnd),
	.asdata(ramiframload_20),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(plif_memwbdmemload_l_20),
	.prn(vcc));
// synopsys translate_off
defparam \plif_memwb.dmemload_l[20] .is_wysiwyg = "true";
defparam \plif_memwb.dmemload_l[20] .power_up = "low";
// synopsys translate_on

// Location: FF_X54_Y39_N13
dffeas \plif_memwb.porto_l[20] (
	.clk(CPUCLK),
	.d(gnd),
	.asdata(plif_exmemporto_l_20),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(plif_memwbporto_l_20),
	.prn(vcc));
// synopsys translate_off
defparam \plif_memwb.porto_l[20] .is_wysiwyg = "true";
defparam \plif_memwb.porto_l[20] .power_up = "low";
// synopsys translate_on

// Location: FF_X54_Y39_N17
dffeas \plif_memwb.rtnaddr_l[20] (
	.clk(CPUCLK),
	.d(gnd),
	.asdata(plif_exmemrtnaddr_l_20),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(plif_memwbrtnaddr_l_20),
	.prn(vcc));
// synopsys translate_off
defparam \plif_memwb.rtnaddr_l[20] .is_wysiwyg = "true";
defparam \plif_memwb.rtnaddr_l[20] .power_up = "low";
// synopsys translate_on

// Location: FF_X56_Y34_N29
dffeas \plif_memwb.dmemload_l[19] (
	.clk(CPUCLK),
	.d(gnd),
	.asdata(ramiframload_19),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(plif_memwbdmemload_l_19),
	.prn(vcc));
// synopsys translate_off
defparam \plif_memwb.dmemload_l[19] .is_wysiwyg = "true";
defparam \plif_memwb.dmemload_l[19] .power_up = "low";
// synopsys translate_on

// Location: FF_X56_Y34_N15
dffeas \plif_memwb.porto_l[19] (
	.clk(CPUCLK),
	.d(\plif_memwb.porto_l[19]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(plif_memwbporto_l_19),
	.prn(vcc));
// synopsys translate_off
defparam \plif_memwb.porto_l[19] .is_wysiwyg = "true";
defparam \plif_memwb.porto_l[19] .power_up = "low";
// synopsys translate_on

// Location: FF_X56_Y34_N25
dffeas \plif_memwb.rtnaddr_l[19] (
	.clk(CPUCLK),
	.d(gnd),
	.asdata(plif_exmemrtnaddr_l_19),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(plif_memwbrtnaddr_l_19),
	.prn(vcc));
// synopsys translate_off
defparam \plif_memwb.rtnaddr_l[19] .is_wysiwyg = "true";
defparam \plif_memwb.rtnaddr_l[19] .power_up = "low";
// synopsys translate_on

// Location: FF_X55_Y37_N13
dffeas \plif_memwb.dmemload_l[18] (
	.clk(CPUCLK),
	.d(gnd),
	.asdata(ramiframload_18),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(plif_memwbdmemload_l_18),
	.prn(vcc));
// synopsys translate_off
defparam \plif_memwb.dmemload_l[18] .is_wysiwyg = "true";
defparam \plif_memwb.dmemload_l[18] .power_up = "low";
// synopsys translate_on

// Location: FF_X55_Y37_N7
dffeas \plif_memwb.porto_l[18] (
	.clk(CPUCLK),
	.d(gnd),
	.asdata(plif_exmemporto_l_18),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(plif_memwbporto_l_18),
	.prn(vcc));
// synopsys translate_off
defparam \plif_memwb.porto_l[18] .is_wysiwyg = "true";
defparam \plif_memwb.porto_l[18] .power_up = "low";
// synopsys translate_on

// Location: FF_X55_Y37_N15
dffeas \plif_memwb.rtnaddr_l[18] (
	.clk(CPUCLK),
	.d(gnd),
	.asdata(plif_exmemrtnaddr_l_18),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(plif_memwbrtnaddr_l_18),
	.prn(vcc));
// synopsys translate_off
defparam \plif_memwb.rtnaddr_l[18] .is_wysiwyg = "true";
defparam \plif_memwb.rtnaddr_l[18] .power_up = "low";
// synopsys translate_on

// Location: FF_X56_Y35_N7
dffeas \plif_memwb.dmemload_l[17] (
	.clk(CPUCLK),
	.d(gnd),
	.asdata(ramiframload_17),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(plif_memwbdmemload_l_17),
	.prn(vcc));
// synopsys translate_off
defparam \plif_memwb.dmemload_l[17] .is_wysiwyg = "true";
defparam \plif_memwb.dmemload_l[17] .power_up = "low";
// synopsys translate_on

// Location: FF_X56_Y35_N9
dffeas \plif_memwb.porto_l[17] (
	.clk(CPUCLK),
	.d(gnd),
	.asdata(plif_exmemporto_l_17),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(plif_memwbporto_l_17),
	.prn(vcc));
// synopsys translate_off
defparam \plif_memwb.porto_l[17] .is_wysiwyg = "true";
defparam \plif_memwb.porto_l[17] .power_up = "low";
// synopsys translate_on

// Location: FF_X56_Y35_N25
dffeas \plif_memwb.rtnaddr_l[17] (
	.clk(CPUCLK),
	.d(gnd),
	.asdata(plif_exmemrtnaddr_l_17),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(plif_memwbrtnaddr_l_17),
	.prn(vcc));
// synopsys translate_off
defparam \plif_memwb.rtnaddr_l[17] .is_wysiwyg = "true";
defparam \plif_memwb.rtnaddr_l[17] .power_up = "low";
// synopsys translate_on

// Location: FF_X55_Y35_N1
dffeas \plif_memwb.dmemload_l[16] (
	.clk(CPUCLK),
	.d(gnd),
	.asdata(ramiframload_16),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(plif_memwbdmemload_l_16),
	.prn(vcc));
// synopsys translate_off
defparam \plif_memwb.dmemload_l[16] .is_wysiwyg = "true";
defparam \plif_memwb.dmemload_l[16] .power_up = "low";
// synopsys translate_on

// Location: FF_X55_Y35_N15
dffeas \plif_memwb.porto_l[16] (
	.clk(CPUCLK),
	.d(gnd),
	.asdata(plif_exmemporto_l_16),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(plif_memwbporto_l_16),
	.prn(vcc));
// synopsys translate_off
defparam \plif_memwb.porto_l[16] .is_wysiwyg = "true";
defparam \plif_memwb.porto_l[16] .power_up = "low";
// synopsys translate_on

// Location: FF_X55_Y35_N9
dffeas \plif_memwb.rtnaddr_l[16] (
	.clk(CPUCLK),
	.d(\plif_memwb.rtnaddr_l[16]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(plif_memwbrtnaddr_l_16),
	.prn(vcc));
// synopsys translate_off
defparam \plif_memwb.rtnaddr_l[16] .is_wysiwyg = "true";
defparam \plif_memwb.rtnaddr_l[16] .power_up = "low";
// synopsys translate_on

// Location: FF_X57_Y38_N25
dffeas \plif_memwb.dmemload_l[15] (
	.clk(CPUCLK),
	.d(gnd),
	.asdata(ramiframload_15),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(plif_memwbdmemload_l_15),
	.prn(vcc));
// synopsys translate_off
defparam \plif_memwb.dmemload_l[15] .is_wysiwyg = "true";
defparam \plif_memwb.dmemload_l[15] .power_up = "low";
// synopsys translate_on

// Location: FF_X56_Y36_N11
dffeas \plif_memwb.porto_l[15] (
	.clk(CPUCLK),
	.d(gnd),
	.asdata(plif_exmemporto_l_15),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(plif_memwbporto_l_15),
	.prn(vcc));
// synopsys translate_off
defparam \plif_memwb.porto_l[15] .is_wysiwyg = "true";
defparam \plif_memwb.porto_l[15] .power_up = "low";
// synopsys translate_on

// Location: FF_X57_Y38_N3
dffeas \plif_memwb.rtnaddr_l[15] (
	.clk(CPUCLK),
	.d(gnd),
	.asdata(plif_exmemrtnaddr_l_15),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(plif_memwbrtnaddr_l_15),
	.prn(vcc));
// synopsys translate_off
defparam \plif_memwb.rtnaddr_l[15] .is_wysiwyg = "true";
defparam \plif_memwb.rtnaddr_l[15] .power_up = "low";
// synopsys translate_on

// Location: FF_X58_Y35_N3
dffeas \plif_memwb.dmemload_l[14] (
	.clk(CPUCLK),
	.d(gnd),
	.asdata(ramiframload_14),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(plif_memwbdmemload_l_14),
	.prn(vcc));
// synopsys translate_off
defparam \plif_memwb.dmemload_l[14] .is_wysiwyg = "true";
defparam \plif_memwb.dmemload_l[14] .power_up = "low";
// synopsys translate_on

// Location: FF_X58_Y35_N29
dffeas \plif_memwb.porto_l[14] (
	.clk(CPUCLK),
	.d(gnd),
	.asdata(plif_exmemporto_l_14),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(plif_memwbporto_l_14),
	.prn(vcc));
// synopsys translate_off
defparam \plif_memwb.porto_l[14] .is_wysiwyg = "true";
defparam \plif_memwb.porto_l[14] .power_up = "low";
// synopsys translate_on

// Location: FF_X58_Y35_N31
dffeas \plif_memwb.rtnaddr_l[14] (
	.clk(CPUCLK),
	.d(gnd),
	.asdata(plif_exmemrtnaddr_l_14),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(plif_memwbrtnaddr_l_14),
	.prn(vcc));
// synopsys translate_off
defparam \plif_memwb.rtnaddr_l[14] .is_wysiwyg = "true";
defparam \plif_memwb.rtnaddr_l[14] .power_up = "low";
// synopsys translate_on

// Location: FF_X57_Y38_N1
dffeas \plif_memwb.dmemload_l[13] (
	.clk(CPUCLK),
	.d(gnd),
	.asdata(ramiframload_13),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(plif_memwbdmemload_l_13),
	.prn(vcc));
// synopsys translate_off
defparam \plif_memwb.dmemload_l[13] .is_wysiwyg = "true";
defparam \plif_memwb.dmemload_l[13] .power_up = "low";
// synopsys translate_on

// Location: FF_X57_Y38_N7
dffeas \plif_memwb.porto_l[13] (
	.clk(CPUCLK),
	.d(gnd),
	.asdata(plif_exmemporto_l_13),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(plif_memwbporto_l_13),
	.prn(vcc));
// synopsys translate_off
defparam \plif_memwb.porto_l[13] .is_wysiwyg = "true";
defparam \plif_memwb.porto_l[13] .power_up = "low";
// synopsys translate_on

// Location: FF_X57_Y38_N9
dffeas \plif_memwb.rtnaddr_l[13] (
	.clk(CPUCLK),
	.d(gnd),
	.asdata(plif_exmemrtnaddr_l_13),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(plif_memwbrtnaddr_l_13),
	.prn(vcc));
// synopsys translate_off
defparam \plif_memwb.rtnaddr_l[13] .is_wysiwyg = "true";
defparam \plif_memwb.rtnaddr_l[13] .power_up = "low";
// synopsys translate_on

// Location: FF_X57_Y34_N27
dffeas \plif_memwb.dmemload_l[12] (
	.clk(CPUCLK),
	.d(gnd),
	.asdata(ramiframload_12),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(plif_memwbdmemload_l_12),
	.prn(vcc));
// synopsys translate_off
defparam \plif_memwb.dmemload_l[12] .is_wysiwyg = "true";
defparam \plif_memwb.dmemload_l[12] .power_up = "low";
// synopsys translate_on

// Location: FF_X57_Y34_N13
dffeas \plif_memwb.porto_l[12] (
	.clk(CPUCLK),
	.d(gnd),
	.asdata(plif_exmemporto_l_12),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(plif_memwbporto_l_12),
	.prn(vcc));
// synopsys translate_off
defparam \plif_memwb.porto_l[12] .is_wysiwyg = "true";
defparam \plif_memwb.porto_l[12] .power_up = "low";
// synopsys translate_on

// Location: FF_X57_Y34_N3
dffeas \plif_memwb.rtnaddr_l[12] (
	.clk(CPUCLK),
	.d(gnd),
	.asdata(plif_exmemrtnaddr_l_12),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(plif_memwbrtnaddr_l_12),
	.prn(vcc));
// synopsys translate_off
defparam \plif_memwb.rtnaddr_l[12] .is_wysiwyg = "true";
defparam \plif_memwb.rtnaddr_l[12] .power_up = "low";
// synopsys translate_on

// Location: FF_X58_Y38_N9
dffeas \plif_memwb.dmemload_l[11] (
	.clk(CPUCLK),
	.d(gnd),
	.asdata(ramiframload_11),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(plif_memwbdmemload_l_11),
	.prn(vcc));
// synopsys translate_off
defparam \plif_memwb.dmemload_l[11] .is_wysiwyg = "true";
defparam \plif_memwb.dmemload_l[11] .power_up = "low";
// synopsys translate_on

// Location: FF_X58_Y38_N23
dffeas \plif_memwb.porto_l[11] (
	.clk(CPUCLK),
	.d(gnd),
	.asdata(plif_exmemporto_l_11),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(plif_memwbporto_l_11),
	.prn(vcc));
// synopsys translate_off
defparam \plif_memwb.porto_l[11] .is_wysiwyg = "true";
defparam \plif_memwb.porto_l[11] .power_up = "low";
// synopsys translate_on

// Location: FF_X58_Y38_N5
dffeas \plif_memwb.rtnaddr_l[11] (
	.clk(CPUCLK),
	.d(gnd),
	.asdata(plif_exmemrtnaddr_l_11),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(plif_memwbrtnaddr_l_11),
	.prn(vcc));
// synopsys translate_off
defparam \plif_memwb.rtnaddr_l[11] .is_wysiwyg = "true";
defparam \plif_memwb.rtnaddr_l[11] .power_up = "low";
// synopsys translate_on

// Location: FF_X56_Y34_N31
dffeas \plif_memwb.dmemload_l[10] (
	.clk(CPUCLK),
	.d(gnd),
	.asdata(ramiframload_10),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(plif_memwbdmemload_l_10),
	.prn(vcc));
// synopsys translate_off
defparam \plif_memwb.dmemload_l[10] .is_wysiwyg = "true";
defparam \plif_memwb.dmemload_l[10] .power_up = "low";
// synopsys translate_on

// Location: FF_X56_Y34_N9
dffeas \plif_memwb.porto_l[10] (
	.clk(CPUCLK),
	.d(\plif_memwb.porto_l[10]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(plif_memwbporto_l_10),
	.prn(vcc));
// synopsys translate_off
defparam \plif_memwb.porto_l[10] .is_wysiwyg = "true";
defparam \plif_memwb.porto_l[10] .power_up = "low";
// synopsys translate_on

// Location: FF_X56_Y34_N19
dffeas \plif_memwb.rtnaddr_l[10] (
	.clk(CPUCLK),
	.d(gnd),
	.asdata(plif_exmemrtnaddr_l_10),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(plif_memwbrtnaddr_l_10),
	.prn(vcc));
// synopsys translate_off
defparam \plif_memwb.rtnaddr_l[10] .is_wysiwyg = "true";
defparam \plif_memwb.rtnaddr_l[10] .power_up = "low";
// synopsys translate_on

// Location: FF_X58_Y35_N11
dffeas \plif_memwb.dmemload_l[9] (
	.clk(CPUCLK),
	.d(gnd),
	.asdata(ramiframload_9),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(plif_memwbdmemload_l_9),
	.prn(vcc));
// synopsys translate_off
defparam \plif_memwb.dmemload_l[9] .is_wysiwyg = "true";
defparam \plif_memwb.dmemload_l[9] .power_up = "low";
// synopsys translate_on

// Location: FF_X58_Y35_N13
dffeas \plif_memwb.porto_l[9] (
	.clk(CPUCLK),
	.d(\plif_memwb.porto_l[9]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(plif_memwbporto_l_9),
	.prn(vcc));
// synopsys translate_off
defparam \plif_memwb.porto_l[9] .is_wysiwyg = "true";
defparam \plif_memwb.porto_l[9] .power_up = "low";
// synopsys translate_on

// Location: FF_X58_Y35_N27
dffeas \plif_memwb.rtnaddr_l[9] (
	.clk(CPUCLK),
	.d(\plif_memwb.rtnaddr_l[9]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(plif_memwbrtnaddr_l_9),
	.prn(vcc));
// synopsys translate_off
defparam \plif_memwb.rtnaddr_l[9] .is_wysiwyg = "true";
defparam \plif_memwb.rtnaddr_l[9] .power_up = "low";
// synopsys translate_on

// Location: FF_X55_Y33_N3
dffeas \plif_memwb.dmemload_l[8] (
	.clk(CPUCLK),
	.d(gnd),
	.asdata(ramiframload_8),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(plif_memwbdmemload_l_8),
	.prn(vcc));
// synopsys translate_off
defparam \plif_memwb.dmemload_l[8] .is_wysiwyg = "true";
defparam \plif_memwb.dmemload_l[8] .power_up = "low";
// synopsys translate_on

// Location: FF_X55_Y33_N9
dffeas \plif_memwb.porto_l[8] (
	.clk(CPUCLK),
	.d(\plif_memwb.porto_l[8]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(plif_memwbporto_l_8),
	.prn(vcc));
// synopsys translate_off
defparam \plif_memwb.porto_l[8] .is_wysiwyg = "true";
defparam \plif_memwb.porto_l[8] .power_up = "low";
// synopsys translate_on

// Location: FF_X55_Y33_N23
dffeas \plif_memwb.rtnaddr_l[8] (
	.clk(CPUCLK),
	.d(gnd),
	.asdata(plif_exmemrtnaddr_l_8),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(plif_memwbrtnaddr_l_8),
	.prn(vcc));
// synopsys translate_off
defparam \plif_memwb.rtnaddr_l[8] .is_wysiwyg = "true";
defparam \plif_memwb.rtnaddr_l[8] .power_up = "low";
// synopsys translate_on

// Location: FF_X56_Y38_N1
dffeas \plif_memwb.dmemload_l[7] (
	.clk(CPUCLK),
	.d(gnd),
	.asdata(ramiframload_7),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(plif_memwbdmemload_l_7),
	.prn(vcc));
// synopsys translate_off
defparam \plif_memwb.dmemload_l[7] .is_wysiwyg = "true";
defparam \plif_memwb.dmemload_l[7] .power_up = "low";
// synopsys translate_on

// Location: FF_X56_Y38_N31
dffeas \plif_memwb.porto_l[7] (
	.clk(CPUCLK),
	.d(gnd),
	.asdata(plif_exmemporto_l_7),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(plif_memwbporto_l_7),
	.prn(vcc));
// synopsys translate_off
defparam \plif_memwb.porto_l[7] .is_wysiwyg = "true";
defparam \plif_memwb.porto_l[7] .power_up = "low";
// synopsys translate_on

// Location: FF_X56_Y38_N17
dffeas \plif_memwb.rtnaddr_l[7] (
	.clk(CPUCLK),
	.d(gnd),
	.asdata(plif_exmemrtnaddr_l_7),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(plif_memwbrtnaddr_l_7),
	.prn(vcc));
// synopsys translate_off
defparam \plif_memwb.rtnaddr_l[7] .is_wysiwyg = "true";
defparam \plif_memwb.rtnaddr_l[7] .power_up = "low";
// synopsys translate_on

// Location: FF_X56_Y39_N17
dffeas \plif_memwb.dmemload_l[6] (
	.clk(CPUCLK),
	.d(gnd),
	.asdata(ramiframload_6),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(plif_memwbdmemload_l_6),
	.prn(vcc));
// synopsys translate_off
defparam \plif_memwb.dmemload_l[6] .is_wysiwyg = "true";
defparam \plif_memwb.dmemload_l[6] .power_up = "low";
// synopsys translate_on

// Location: FF_X56_Y39_N5
dffeas \plif_memwb.porto_l[6] (
	.clk(CPUCLK),
	.d(gnd),
	.asdata(plif_exmemporto_l_6),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(plif_memwbporto_l_6),
	.prn(vcc));
// synopsys translate_off
defparam \plif_memwb.porto_l[6] .is_wysiwyg = "true";
defparam \plif_memwb.porto_l[6] .power_up = "low";
// synopsys translate_on

// Location: FF_X56_Y39_N31
dffeas \plif_memwb.rtnaddr_l[6] (
	.clk(CPUCLK),
	.d(gnd),
	.asdata(plif_exmemrtnaddr_l_6),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(plif_memwbrtnaddr_l_6),
	.prn(vcc));
// synopsys translate_off
defparam \plif_memwb.rtnaddr_l[6] .is_wysiwyg = "true";
defparam \plif_memwb.rtnaddr_l[6] .power_up = "low";
// synopsys translate_on

// Location: FF_X56_Y38_N9
dffeas \plif_memwb.dmemload_l[5] (
	.clk(CPUCLK),
	.d(gnd),
	.asdata(ramiframload_5),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(plif_memwbdmemload_l_5),
	.prn(vcc));
// synopsys translate_off
defparam \plif_memwb.dmemload_l[5] .is_wysiwyg = "true";
defparam \plif_memwb.dmemload_l[5] .power_up = "low";
// synopsys translate_on

// Location: FF_X56_Y38_N15
dffeas \plif_memwb.porto_l[5] (
	.clk(CPUCLK),
	.d(gnd),
	.asdata(plif_exmemporto_l_5),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(plif_memwbporto_l_5),
	.prn(vcc));
// synopsys translate_off
defparam \plif_memwb.porto_l[5] .is_wysiwyg = "true";
defparam \plif_memwb.porto_l[5] .power_up = "low";
// synopsys translate_on

// Location: FF_X56_Y38_N29
dffeas \plif_memwb.rtnaddr_l[5] (
	.clk(CPUCLK),
	.d(gnd),
	.asdata(plif_exmemrtnaddr_l_5),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(plif_memwbrtnaddr_l_5),
	.prn(vcc));
// synopsys translate_off
defparam \plif_memwb.rtnaddr_l[5] .is_wysiwyg = "true";
defparam \plif_memwb.rtnaddr_l[5] .power_up = "low";
// synopsys translate_on

// Location: FF_X58_Y35_N7
dffeas \plif_memwb.dmemload_l[2] (
	.clk(CPUCLK),
	.d(gnd),
	.asdata(ramiframload_2),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(plif_memwbdmemload_l_2),
	.prn(vcc));
// synopsys translate_off
defparam \plif_memwb.dmemload_l[2] .is_wysiwyg = "true";
defparam \plif_memwb.dmemload_l[2] .power_up = "low";
// synopsys translate_on

// Location: FF_X58_Y35_N21
dffeas \plif_memwb.porto_l[2] (
	.clk(CPUCLK),
	.d(gnd),
	.asdata(plif_exmemporto_l_2),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(plif_memwbporto_l_2),
	.prn(vcc));
// synopsys translate_off
defparam \plif_memwb.porto_l[2] .is_wysiwyg = "true";
defparam \plif_memwb.porto_l[2] .power_up = "low";
// synopsys translate_on

// Location: FF_X56_Y39_N15
dffeas \plif_memwb.rtnaddr_l[2] (
	.clk(CPUCLK),
	.d(\plif_memwb.rtnaddr_l[2]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(plif_memwbrtnaddr_l_2),
	.prn(vcc));
// synopsys translate_off
defparam \plif_memwb.rtnaddr_l[2] .is_wysiwyg = "true";
defparam \plif_memwb.rtnaddr_l[2] .power_up = "low";
// synopsys translate_on

// Location: FF_X57_Y34_N1
dffeas \plif_memwb.dmemload_l[1] (
	.clk(CPUCLK),
	.d(gnd),
	.asdata(ramiframload_1),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(plif_memwbdmemload_l_1),
	.prn(vcc));
// synopsys translate_off
defparam \plif_memwb.dmemload_l[1] .is_wysiwyg = "true";
defparam \plif_memwb.dmemload_l[1] .power_up = "low";
// synopsys translate_on

// Location: FF_X57_Y34_N23
dffeas \plif_memwb.porto_l[1] (
	.clk(CPUCLK),
	.d(\plif_memwb.porto_l[1]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(plif_memwbporto_l_1),
	.prn(vcc));
// synopsys translate_off
defparam \plif_memwb.porto_l[1] .is_wysiwyg = "true";
defparam \plif_memwb.porto_l[1] .power_up = "low";
// synopsys translate_on

// Location: FF_X57_Y34_N5
dffeas \plif_memwb.rtnaddr_l[1] (
	.clk(CPUCLK),
	.d(\plif_memwb.rtnaddr_l[1]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(plif_memwbrtnaddr_l_1),
	.prn(vcc));
// synopsys translate_off
defparam \plif_memwb.rtnaddr_l[1] .is_wysiwyg = "true";
defparam \plif_memwb.rtnaddr_l[1] .power_up = "low";
// synopsys translate_on

// Location: FF_X56_Y33_N17
dffeas \plif_memwb.dmemload_l[0] (
	.clk(CPUCLK),
	.d(gnd),
	.asdata(ramiframload_0),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(plif_memwbdmemload_l_0),
	.prn(vcc));
// synopsys translate_off
defparam \plif_memwb.dmemload_l[0] .is_wysiwyg = "true";
defparam \plif_memwb.dmemload_l[0] .power_up = "low";
// synopsys translate_on

// Location: FF_X56_Y33_N27
dffeas \plif_memwb.porto_l[0] (
	.clk(CPUCLK),
	.d(\plif_memwb.porto_l[0]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(plif_memwbporto_l_0),
	.prn(vcc));
// synopsys translate_off
defparam \plif_memwb.porto_l[0] .is_wysiwyg = "true";
defparam \plif_memwb.porto_l[0] .power_up = "low";
// synopsys translate_on

// Location: FF_X56_Y33_N1
dffeas \plif_memwb.rtnaddr_l[0] (
	.clk(CPUCLK),
	.d(\plif_memwb.rtnaddr_l[0]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(plif_memwbrtnaddr_l_0),
	.prn(vcc));
// synopsys translate_off
defparam \plif_memwb.rtnaddr_l[0] .is_wysiwyg = "true";
defparam \plif_memwb.rtnaddr_l[0] .power_up = "low";
// synopsys translate_on

// Location: FF_X56_Y33_N21
dffeas \plif_memwb.dmemload_l[4] (
	.clk(CPUCLK),
	.d(gnd),
	.asdata(ramiframload_4),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(plif_memwbdmemload_l_4),
	.prn(vcc));
// synopsys translate_off
defparam \plif_memwb.dmemload_l[4] .is_wysiwyg = "true";
defparam \plif_memwb.dmemload_l[4] .power_up = "low";
// synopsys translate_on

// Location: FF_X56_Y33_N19
dffeas \plif_memwb.porto_l[4] (
	.clk(CPUCLK),
	.d(\plif_memwb.porto_l[4]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(plif_memwbporto_l_4),
	.prn(vcc));
// synopsys translate_off
defparam \plif_memwb.porto_l[4] .is_wysiwyg = "true";
defparam \plif_memwb.porto_l[4] .power_up = "low";
// synopsys translate_on

// Location: FF_X56_Y33_N25
dffeas \plif_memwb.rtnaddr_l[4] (
	.clk(CPUCLK),
	.d(\plif_memwb.rtnaddr_l[4]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(plif_memwbrtnaddr_l_4),
	.prn(vcc));
// synopsys translate_off
defparam \plif_memwb.rtnaddr_l[4] .is_wysiwyg = "true";
defparam \plif_memwb.rtnaddr_l[4] .power_up = "low";
// synopsys translate_on

// Location: FF_X57_Y35_N25
dffeas \plif_memwb.dmemload_l[3] (
	.clk(CPUCLK),
	.d(gnd),
	.asdata(ramiframload_3),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(plif_memwbdmemload_l_3),
	.prn(vcc));
// synopsys translate_off
defparam \plif_memwb.dmemload_l[3] .is_wysiwyg = "true";
defparam \plif_memwb.dmemload_l[3] .power_up = "low";
// synopsys translate_on

// Location: FF_X57_Y35_N11
dffeas \plif_memwb.porto_l[3] (
	.clk(CPUCLK),
	.d(\plif_memwb.porto_l[3]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(plif_memwbporto_l_3),
	.prn(vcc));
// synopsys translate_off
defparam \plif_memwb.porto_l[3] .is_wysiwyg = "true";
defparam \plif_memwb.porto_l[3] .power_up = "low";
// synopsys translate_on

// Location: FF_X57_Y35_N13
dffeas \plif_memwb.rtnaddr_l[3] (
	.clk(CPUCLK),
	.d(\plif_memwb.rtnaddr_l[3]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(plif_memwbrtnaddr_l_3),
	.prn(vcc));
// synopsys translate_off
defparam \plif_memwb.rtnaddr_l[3] .is_wysiwyg = "true";
defparam \plif_memwb.rtnaddr_l[3] .power_up = "low";
// synopsys translate_on

// Location: FF_X55_Y32_N13
dffeas \plif_memwb.btype_l (
	.clk(CPUCLK),
	.d(\plif_memwb.btype_l~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(plif_memwbbtype_l),
	.prn(vcc));
// synopsys translate_off
defparam \plif_memwb.btype_l .is_wysiwyg = "true";
defparam \plif_memwb.btype_l .power_up = "low";
// synopsys translate_on

// Location: FF_X55_Y32_N17
dffeas \plif_memwb.zero_l (
	.clk(CPUCLK),
	.d(gnd),
	.asdata(plif_exmemzero_l),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(plif_memwbzero_l),
	.prn(vcc));
// synopsys translate_off
defparam \plif_memwb.zero_l .is_wysiwyg = "true";
defparam \plif_memwb.zero_l .power_up = "low";
// synopsys translate_on

// Location: FF_X54_Y29_N17
dffeas \plif_memwb.jaddr_l[1] (
	.clk(CPUCLK),
	.d(\plif_memwb.jaddr_l[1]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(plif_memwbjaddr_l_1),
	.prn(vcc));
// synopsys translate_off
defparam \plif_memwb.jaddr_l[1] .is_wysiwyg = "true";
defparam \plif_memwb.jaddr_l[1] .power_up = "low";
// synopsys translate_on

// Location: FF_X56_Y32_N5
dffeas \plif_memwb.extimm_l[1] (
	.clk(CPUCLK),
	.d(gnd),
	.asdata(plif_exmemextimm_l_1),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(plif_memwbextimm_l_1),
	.prn(vcc));
// synopsys translate_off
defparam \plif_memwb.extimm_l[1] .is_wysiwyg = "true";
defparam \plif_memwb.extimm_l[1] .power_up = "low";
// synopsys translate_on

// Location: FF_X56_Y29_N23
dffeas \plif_memwb.extimm_l[0] (
	.clk(CPUCLK),
	.d(\plif_memwb.extimm_l[0]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(plif_memwbextimm_l_0),
	.prn(vcc));
// synopsys translate_off
defparam \plif_memwb.extimm_l[0] .is_wysiwyg = "true";
defparam \plif_memwb.extimm_l[0] .power_up = "low";
// synopsys translate_on

// Location: FF_X52_Y33_N1
dffeas \plif_memwb.jaddr_l[0] (
	.clk(CPUCLK),
	.d(gnd),
	.asdata(plif_exmemjaddr_l_0),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(plif_memwbjaddr_l_0),
	.prn(vcc));
// synopsys translate_off
defparam \plif_memwb.jaddr_l[0] .is_wysiwyg = "true";
defparam \plif_memwb.jaddr_l[0] .power_up = "low";
// synopsys translate_on

// Location: FF_X59_Y39_N17
dffeas \plif_memwb.jaddr_l[3] (
	.clk(CPUCLK),
	.d(gnd),
	.asdata(plif_exmemjaddr_l_3),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(plif_memwbjaddr_l_3),
	.prn(vcc));
// synopsys translate_off
defparam \plif_memwb.jaddr_l[3] .is_wysiwyg = "true";
defparam \plif_memwb.jaddr_l[3] .power_up = "low";
// synopsys translate_on

// Location: FF_X56_Y32_N25
dffeas \plif_memwb.extimm_l[3] (
	.clk(CPUCLK),
	.d(gnd),
	.asdata(plif_exmemextimm_l_3),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(plif_memwbextimm_l_3),
	.prn(vcc));
// synopsys translate_off
defparam \plif_memwb.extimm_l[3] .is_wysiwyg = "true";
defparam \plif_memwb.extimm_l[3] .power_up = "low";
// synopsys translate_on

// Location: FF_X56_Y32_N7
dffeas \plif_memwb.extimm_l[2] (
	.clk(CPUCLK),
	.d(gnd),
	.asdata(plif_exmemextimm_l_2),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(plif_memwbextimm_l_2),
	.prn(vcc));
// synopsys translate_off
defparam \plif_memwb.extimm_l[2] .is_wysiwyg = "true";
defparam \plif_memwb.extimm_l[2] .power_up = "low";
// synopsys translate_on

// Location: FF_X50_Y33_N25
dffeas \plif_memwb.jaddr_l[2] (
	.clk(CPUCLK),
	.d(gnd),
	.asdata(plif_exmemjaddr_l_2),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(plif_memwbjaddr_l_2),
	.prn(vcc));
// synopsys translate_off
defparam \plif_memwb.jaddr_l[2] .is_wysiwyg = "true";
defparam \plif_memwb.jaddr_l[2] .power_up = "low";
// synopsys translate_on

// Location: FF_X57_Y29_N1
dffeas \plif_memwb.jaddr_l[5] (
	.clk(CPUCLK),
	.d(\plif_memwb.jaddr_l[5]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(plif_memwbjaddr_l_5),
	.prn(vcc));
// synopsys translate_off
defparam \plif_memwb.jaddr_l[5] .is_wysiwyg = "true";
defparam \plif_memwb.jaddr_l[5] .power_up = "low";
// synopsys translate_on

// Location: FF_X56_Y32_N9
dffeas \plif_memwb.extimm_l[5] (
	.clk(CPUCLK),
	.d(gnd),
	.asdata(plif_exmemextimm_l_5),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(plif_memwbextimm_l_5),
	.prn(vcc));
// synopsys translate_off
defparam \plif_memwb.extimm_l[5] .is_wysiwyg = "true";
defparam \plif_memwb.extimm_l[5] .power_up = "low";
// synopsys translate_on

// Location: FF_X56_Y32_N27
dffeas \plif_memwb.extimm_l[4] (
	.clk(CPUCLK),
	.d(gnd),
	.asdata(plif_exmemextimm_l_4),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(plif_memwbextimm_l_4),
	.prn(vcc));
// synopsys translate_off
defparam \plif_memwb.extimm_l[4] .is_wysiwyg = "true";
defparam \plif_memwb.extimm_l[4] .power_up = "low";
// synopsys translate_on

// Location: FF_X50_Y33_N11
dffeas \plif_memwb.jaddr_l[4] (
	.clk(CPUCLK),
	.d(gnd),
	.asdata(plif_exmemjaddr_l_4),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(plif_memwbjaddr_l_4),
	.prn(vcc));
// synopsys translate_off
defparam \plif_memwb.jaddr_l[4] .is_wysiwyg = "true";
defparam \plif_memwb.jaddr_l[4] .power_up = "low";
// synopsys translate_on

// Location: FF_X53_Y33_N31
dffeas \plif_memwb.jaddr_l[7] (
	.clk(CPUCLK),
	.d(gnd),
	.asdata(plif_exmemjaddr_l_7),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(plif_memwbjaddr_l_7),
	.prn(vcc));
// synopsys translate_off
defparam \plif_memwb.jaddr_l[7] .is_wysiwyg = "true";
defparam \plif_memwb.jaddr_l[7] .power_up = "low";
// synopsys translate_on

// Location: FF_X57_Y29_N11
dffeas \plif_memwb.extimm_l[7] (
	.clk(CPUCLK),
	.d(\plif_memwb.extimm_l[7]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(plif_memwbextimm_l_7),
	.prn(vcc));
// synopsys translate_off
defparam \plif_memwb.extimm_l[7] .is_wysiwyg = "true";
defparam \plif_memwb.extimm_l[7] .power_up = "low";
// synopsys translate_on

// Location: FF_X56_Y32_N21
dffeas \plif_memwb.extimm_l[6] (
	.clk(CPUCLK),
	.d(gnd),
	.asdata(plif_exmemextimm_l_6),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(plif_memwbextimm_l_6),
	.prn(vcc));
// synopsys translate_off
defparam \plif_memwb.extimm_l[6] .is_wysiwyg = "true";
defparam \plif_memwb.extimm_l[6] .power_up = "low";
// synopsys translate_on

// Location: FF_X55_Y33_N5
dffeas \plif_memwb.jaddr_l[6] (
	.clk(CPUCLK),
	.d(gnd),
	.asdata(plif_exmemjaddr_l_6),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(plif_memwbjaddr_l_6),
	.prn(vcc));
// synopsys translate_off
defparam \plif_memwb.jaddr_l[6] .is_wysiwyg = "true";
defparam \plif_memwb.jaddr_l[6] .power_up = "low";
// synopsys translate_on

// Location: FF_X58_Y32_N13
dffeas \plif_memwb.jaddr_l[9] (
	.clk(CPUCLK),
	.d(\plif_memwb.jaddr_l[9]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(plif_memwbjaddr_l_9),
	.prn(vcc));
// synopsys translate_off
defparam \plif_memwb.jaddr_l[9] .is_wysiwyg = "true";
defparam \plif_memwb.jaddr_l[9] .power_up = "low";
// synopsys translate_on

// Location: FF_X58_Y32_N15
dffeas \plif_memwb.extimm_l[9] (
	.clk(CPUCLK),
	.d(gnd),
	.asdata(plif_exmemextimm_l_9),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(plif_memwbextimm_l_9),
	.prn(vcc));
// synopsys translate_off
defparam \plif_memwb.extimm_l[9] .is_wysiwyg = "true";
defparam \plif_memwb.extimm_l[9] .power_up = "low";
// synopsys translate_on

// Location: FF_X58_Y32_N9
dffeas \plif_memwb.extimm_l[8] (
	.clk(CPUCLK),
	.d(\plif_memwb.extimm_l[8]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(plif_memwbextimm_l_8),
	.prn(vcc));
// synopsys translate_off
defparam \plif_memwb.extimm_l[8] .is_wysiwyg = "true";
defparam \plif_memwb.extimm_l[8] .power_up = "low";
// synopsys translate_on

// Location: FF_X56_Y34_N5
dffeas \plif_memwb.jaddr_l[8] (
	.clk(CPUCLK),
	.d(gnd),
	.asdata(plif_exmemjaddr_l_8),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(plif_memwbjaddr_l_8),
	.prn(vcc));
// synopsys translate_off
defparam \plif_memwb.jaddr_l[8] .is_wysiwyg = "true";
defparam \plif_memwb.jaddr_l[8] .power_up = "low";
// synopsys translate_on

// Location: FF_X58_Y32_N7
dffeas \plif_memwb.jaddr_l[11] (
	.clk(CPUCLK),
	.d(\plif_memwb.jaddr_l[11]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(plif_memwbjaddr_l_11),
	.prn(vcc));
// synopsys translate_off
defparam \plif_memwb.jaddr_l[11] .is_wysiwyg = "true";
defparam \plif_memwb.jaddr_l[11] .power_up = "low";
// synopsys translate_on

// Location: FF_X58_Y32_N17
dffeas \plif_memwb.extimm_l[11] (
	.clk(CPUCLK),
	.d(\plif_memwb.extimm_l[11]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(plif_memwbextimm_l_11),
	.prn(vcc));
// synopsys translate_off
defparam \plif_memwb.extimm_l[11] .is_wysiwyg = "true";
defparam \plif_memwb.extimm_l[11] .power_up = "low";
// synopsys translate_on

// Location: FF_X58_Y32_N27
dffeas \plif_memwb.extimm_l[10] (
	.clk(CPUCLK),
	.d(gnd),
	.asdata(plif_exmemextimm_l_10),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(plif_memwbextimm_l_10),
	.prn(vcc));
// synopsys translate_off
defparam \plif_memwb.extimm_l[10] .is_wysiwyg = "true";
defparam \plif_memwb.extimm_l[10] .power_up = "low";
// synopsys translate_on

// Location: FF_X50_Y33_N15
dffeas \plif_memwb.jaddr_l[10] (
	.clk(CPUCLK),
	.d(gnd),
	.asdata(plif_exmemjaddr_l_10),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(plif_memwbjaddr_l_10),
	.prn(vcc));
// synopsys translate_off
defparam \plif_memwb.jaddr_l[10] .is_wysiwyg = "true";
defparam \plif_memwb.jaddr_l[10] .power_up = "low";
// synopsys translate_on

// Location: FF_X58_Y32_N29
dffeas \plif_memwb.jaddr_l[13] (
	.clk(CPUCLK),
	.d(gnd),
	.asdata(plif_exmemjaddr_l_13),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(plif_memwbjaddr_l_13),
	.prn(vcc));
// synopsys translate_off
defparam \plif_memwb.jaddr_l[13] .is_wysiwyg = "true";
defparam \plif_memwb.jaddr_l[13] .power_up = "low";
// synopsys translate_on

// Location: FF_X56_Y32_N3
dffeas \plif_memwb.extimm_l[13] (
	.clk(CPUCLK),
	.d(gnd),
	.asdata(plif_exmemextimm_l_13),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(plif_memwbextimm_l_13),
	.prn(vcc));
// synopsys translate_off
defparam \plif_memwb.extimm_l[13] .is_wysiwyg = "true";
defparam \plif_memwb.extimm_l[13] .power_up = "low";
// synopsys translate_on

// Location: FF_X60_Y31_N13
dffeas \plif_memwb.extimm_l[12] (
	.clk(CPUCLK),
	.d(\plif_memwb.extimm_l[12]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(plif_memwbextimm_l_12),
	.prn(vcc));
// synopsys translate_off
defparam \plif_memwb.extimm_l[12] .is_wysiwyg = "true";
defparam \plif_memwb.extimm_l[12] .power_up = "low";
// synopsys translate_on

// Location: FF_X50_Y33_N3
dffeas \plif_memwb.jaddr_l[12] (
	.clk(CPUCLK),
	.d(gnd),
	.asdata(plif_exmemjaddr_l_12),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(plif_memwbjaddr_l_12),
	.prn(vcc));
// synopsys translate_off
defparam \plif_memwb.jaddr_l[12] .is_wysiwyg = "true";
defparam \plif_memwb.jaddr_l[12] .power_up = "low";
// synopsys translate_on

// Location: FF_X60_Y31_N27
dffeas \plif_memwb.jaddr_l[15] (
	.clk(CPUCLK),
	.d(\plif_memwb.jaddr_l[15]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(plif_memwbjaddr_l_15),
	.prn(vcc));
// synopsys translate_off
defparam \plif_memwb.jaddr_l[15] .is_wysiwyg = "true";
defparam \plif_memwb.jaddr_l[15] .power_up = "low";
// synopsys translate_on

// Location: FF_X60_Y31_N21
dffeas \plif_memwb.extimm_l[15] (
	.clk(CPUCLK),
	.d(\plif_memwb.extimm_l[15]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(plif_memwbextimm_l_15),
	.prn(vcc));
// synopsys translate_off
defparam \plif_memwb.extimm_l[15] .is_wysiwyg = "true";
defparam \plif_memwb.extimm_l[15] .power_up = "low";
// synopsys translate_on

// Location: FF_X60_Y31_N7
dffeas \plif_memwb.extimm_l[14] (
	.clk(CPUCLK),
	.d(\plif_memwb.extimm_l[14]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(plif_memwbextimm_l_14),
	.prn(vcc));
// synopsys translate_off
defparam \plif_memwb.extimm_l[14] .is_wysiwyg = "true";
defparam \plif_memwb.extimm_l[14] .power_up = "low";
// synopsys translate_on

// Location: FF_X50_Y33_N1
dffeas \plif_memwb.jaddr_l[14] (
	.clk(CPUCLK),
	.d(gnd),
	.asdata(plif_exmemjaddr_l_14),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(plif_memwbjaddr_l_14),
	.prn(vcc));
// synopsys translate_off
defparam \plif_memwb.jaddr_l[14] .is_wysiwyg = "true";
defparam \plif_memwb.jaddr_l[14] .power_up = "low";
// synopsys translate_on

// Location: FF_X53_Y32_N1
dffeas \plif_memwb.jaddr_l[17] (
	.clk(CPUCLK),
	.d(\plif_memwb.jaddr_l[17]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(plif_memwbjaddr_l_17),
	.prn(vcc));
// synopsys translate_off
defparam \plif_memwb.jaddr_l[17] .is_wysiwyg = "true";
defparam \plif_memwb.jaddr_l[17] .power_up = "low";
// synopsys translate_on

// Location: FF_X55_Y31_N29
dffeas \plif_memwb.extimm_l[17] (
	.clk(CPUCLK),
	.d(\plif_memwb.extimm_l[17]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(plif_memwbextimm_l_17),
	.prn(vcc));
// synopsys translate_off
defparam \plif_memwb.extimm_l[17] .is_wysiwyg = "true";
defparam \plif_memwb.extimm_l[17] .power_up = "low";
// synopsys translate_on

// Location: FF_X56_Y31_N25
dffeas \plif_memwb.extimm_l[16] (
	.clk(CPUCLK),
	.d(gnd),
	.asdata(plif_exmemextimm_l_16),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(plif_memwbextimm_l_16),
	.prn(vcc));
// synopsys translate_off
defparam \plif_memwb.extimm_l[16] .is_wysiwyg = "true";
defparam \plif_memwb.extimm_l[16] .power_up = "low";
// synopsys translate_on

// Location: FF_X53_Y33_N3
dffeas \plif_memwb.jaddr_l[16] (
	.clk(CPUCLK),
	.d(gnd),
	.asdata(plif_exmemjaddr_l_16),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(plif_memwbjaddr_l_16),
	.prn(vcc));
// synopsys translate_off
defparam \plif_memwb.jaddr_l[16] .is_wysiwyg = "true";
defparam \plif_memwb.jaddr_l[16] .power_up = "low";
// synopsys translate_on

// Location: FF_X53_Y33_N9
dffeas \plif_memwb.jaddr_l[19] (
	.clk(CPUCLK),
	.d(\plif_memwb.jaddr_l[19]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(plif_memwbjaddr_l_19),
	.prn(vcc));
// synopsys translate_off
defparam \plif_memwb.jaddr_l[19] .is_wysiwyg = "true";
defparam \plif_memwb.jaddr_l[19] .power_up = "low";
// synopsys translate_on

// Location: FF_X56_Y31_N29
dffeas \plif_memwb.extimm_l[19] (
	.clk(CPUCLK),
	.d(gnd),
	.asdata(plif_exmemextimm_l_19),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(plif_memwbextimm_l_19),
	.prn(vcc));
// synopsys translate_off
defparam \plif_memwb.extimm_l[19] .is_wysiwyg = "true";
defparam \plif_memwb.extimm_l[19] .power_up = "low";
// synopsys translate_on

// Location: FF_X55_Y31_N15
dffeas \plif_memwb.extimm_l[18] (
	.clk(CPUCLK),
	.d(\plif_memwb.extimm_l[18]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(plif_memwbextimm_l_18),
	.prn(vcc));
// synopsys translate_off
defparam \plif_memwb.extimm_l[18] .is_wysiwyg = "true";
defparam \plif_memwb.extimm_l[18] .power_up = "low";
// synopsys translate_on

// Location: FF_X53_Y33_N15
dffeas \plif_memwb.jaddr_l[18] (
	.clk(CPUCLK),
	.d(gnd),
	.asdata(plif_exmemjaddr_l_18),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(plif_memwbjaddr_l_18),
	.prn(vcc));
// synopsys translate_off
defparam \plif_memwb.jaddr_l[18] .is_wysiwyg = "true";
defparam \plif_memwb.jaddr_l[18] .power_up = "low";
// synopsys translate_on

// Location: FF_X55_Y31_N1
dffeas \plif_memwb.jaddr_l[21] (
	.clk(CPUCLK),
	.d(\plif_memwb.jaddr_l[21]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(plif_memwbjaddr_l_21),
	.prn(vcc));
// synopsys translate_off
defparam \plif_memwb.jaddr_l[21] .is_wysiwyg = "true";
defparam \plif_memwb.jaddr_l[21] .power_up = "low";
// synopsys translate_on

// Location: FF_X55_Y31_N31
dffeas \plif_memwb.extimm_l[21] (
	.clk(CPUCLK),
	.d(gnd),
	.asdata(plif_exmemextimm_l_21),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(plif_memwbextimm_l_21),
	.prn(vcc));
// synopsys translate_off
defparam \plif_memwb.extimm_l[21] .is_wysiwyg = "true";
defparam \plif_memwb.extimm_l[21] .power_up = "low";
// synopsys translate_on

// Location: FF_X56_Y31_N5
dffeas \plif_memwb.extimm_l[20] (
	.clk(CPUCLK),
	.d(gnd),
	.asdata(plif_exmemextimm_l_20),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(plif_memwbextimm_l_20),
	.prn(vcc));
// synopsys translate_off
defparam \plif_memwb.extimm_l[20] .is_wysiwyg = "true";
defparam \plif_memwb.extimm_l[20] .power_up = "low";
// synopsys translate_on

// Location: FF_X53_Y33_N5
dffeas \plif_memwb.jaddr_l[20] (
	.clk(CPUCLK),
	.d(gnd),
	.asdata(plif_exmemjaddr_l_20),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(plif_memwbjaddr_l_20),
	.prn(vcc));
// synopsys translate_off
defparam \plif_memwb.jaddr_l[20] .is_wysiwyg = "true";
defparam \plif_memwb.jaddr_l[20] .power_up = "low";
// synopsys translate_on

// Location: FF_X58_Y35_N9
dffeas \plif_memwb.jaddr_l[23] (
	.clk(CPUCLK),
	.d(gnd),
	.asdata(plif_exmemjaddr_l_23),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(plif_memwbjaddr_l_23),
	.prn(vcc));
// synopsys translate_off
defparam \plif_memwb.jaddr_l[23] .is_wysiwyg = "true";
defparam \plif_memwb.jaddr_l[23] .power_up = "low";
// synopsys translate_on

// Location: FF_X55_Y31_N25
dffeas \plif_memwb.extimm_l[23] (
	.clk(CPUCLK),
	.d(\plif_memwb.extimm_l[23]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(plif_memwbextimm_l_23),
	.prn(vcc));
// synopsys translate_off
defparam \plif_memwb.extimm_l[23] .is_wysiwyg = "true";
defparam \plif_memwb.extimm_l[23] .power_up = "low";
// synopsys translate_on

// Location: FF_X56_Y31_N13
dffeas \plif_memwb.extimm_l[22] (
	.clk(CPUCLK),
	.d(gnd),
	.asdata(plif_exmemextimm_l_22),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(plif_memwbextimm_l_22),
	.prn(vcc));
// synopsys translate_off
defparam \plif_memwb.extimm_l[22] .is_wysiwyg = "true";
defparam \plif_memwb.extimm_l[22] .power_up = "low";
// synopsys translate_on

// Location: FF_X53_Y33_N19
dffeas \plif_memwb.jaddr_l[22] (
	.clk(CPUCLK),
	.d(gnd),
	.asdata(plif_exmemjaddr_l_22),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(plif_memwbjaddr_l_22),
	.prn(vcc));
// synopsys translate_off
defparam \plif_memwb.jaddr_l[22] .is_wysiwyg = "true";
defparam \plif_memwb.jaddr_l[22] .power_up = "low";
// synopsys translate_on

// Location: FF_X55_Y31_N7
dffeas \plif_memwb.jaddr_l[25] (
	.clk(CPUCLK),
	.d(\plif_memwb.jaddr_l[25]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(plif_memwbjaddr_l_25),
	.prn(vcc));
// synopsys translate_off
defparam \plif_memwb.jaddr_l[25] .is_wysiwyg = "true";
defparam \plif_memwb.jaddr_l[25] .power_up = "low";
// synopsys translate_on

// Location: FF_X56_Y31_N9
dffeas \plif_memwb.extimm_l[25] (
	.clk(CPUCLK),
	.d(gnd),
	.asdata(plif_exmemextimm_l_25),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(plif_memwbextimm_l_25),
	.prn(vcc));
// synopsys translate_off
defparam \plif_memwb.extimm_l[25] .is_wysiwyg = "true";
defparam \plif_memwb.extimm_l[25] .power_up = "low";
// synopsys translate_on

// Location: FF_X56_Y28_N5
dffeas \plif_memwb.extimm_l[24] (
	.clk(CPUCLK),
	.d(\plif_memwb.extimm_l[24]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(plif_memwbextimm_l_24),
	.prn(vcc));
// synopsys translate_off
defparam \plif_memwb.extimm_l[24] .is_wysiwyg = "true";
defparam \plif_memwb.extimm_l[24] .power_up = "low";
// synopsys translate_on

// Location: FF_X55_Y33_N15
dffeas \plif_memwb.jaddr_l[24] (
	.clk(CPUCLK),
	.d(gnd),
	.asdata(plif_exmemjaddr_l_24),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(plif_memwbjaddr_l_24),
	.prn(vcc));
// synopsys translate_off
defparam \plif_memwb.jaddr_l[24] .is_wysiwyg = "true";
defparam \plif_memwb.jaddr_l[24] .power_up = "low";
// synopsys translate_on

// Location: FF_X56_Y31_N23
dffeas \plif_memwb.extimm_l[27] (
	.clk(CPUCLK),
	.d(gnd),
	.asdata(plif_exmemextimm_l_27),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(plif_memwbextimm_l_27),
	.prn(vcc));
// synopsys translate_off
defparam \plif_memwb.extimm_l[27] .is_wysiwyg = "true";
defparam \plif_memwb.extimm_l[27] .power_up = "low";
// synopsys translate_on

// Location: FF_X56_Y31_N21
dffeas \plif_memwb.extimm_l[26] (
	.clk(CPUCLK),
	.d(gnd),
	.asdata(plif_exmemextimm_l_26),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(plif_memwbextimm_l_26),
	.prn(vcc));
// synopsys translate_off
defparam \plif_memwb.extimm_l[26] .is_wysiwyg = "true";
defparam \plif_memwb.extimm_l[26] .power_up = "low";
// synopsys translate_on

// Location: FF_X56_Y31_N1
dffeas \plif_memwb.extimm_l[29] (
	.clk(CPUCLK),
	.d(gnd),
	.asdata(plif_exmemextimm_l_29),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(plif_memwbextimm_l_29),
	.prn(vcc));
// synopsys translate_off
defparam \plif_memwb.extimm_l[29] .is_wysiwyg = "true";
defparam \plif_memwb.extimm_l[29] .power_up = "low";
// synopsys translate_on

// Location: FF_X55_Y31_N9
dffeas \plif_memwb.extimm_l[28] (
	.clk(CPUCLK),
	.d(\plif_memwb.extimm_l[28]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(plif_memwbextimm_l_28),
	.prn(vcc));
// synopsys translate_off
defparam \plif_memwb.extimm_l[28] .is_wysiwyg = "true";
defparam \plif_memwb.extimm_l[28] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X56_Y35_N4
cycloneive_lcell_comb \plif_memwb.regsrc_l[0]~feeder (
// Equation(s):
// \plif_memwb.regsrc_l[0]~feeder_combout  = plif_exmemregsrc_l_0

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(plif_exmemregsrc_l_0),
	.cin(gnd),
	.combout(\plif_memwb.regsrc_l[0]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \plif_memwb.regsrc_l[0]~feeder .lut_mask = 16'hFF00;
defparam \plif_memwb.regsrc_l[0]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y35_N30
cycloneive_lcell_comb \plif_memwb.regsrc_l[1]~feeder (
// Equation(s):
// \plif_memwb.regsrc_l[1]~feeder_combout  = plif_exmemregsrc_l_1

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(plif_exmemregsrc_l_1),
	.cin(gnd),
	.combout(\plif_memwb.regsrc_l[1]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \plif_memwb.regsrc_l[1]~feeder .lut_mask = 16'hFF00;
defparam \plif_memwb.regsrc_l[1]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y35_N28
cycloneive_lcell_comb \plif_memwb.porto_l[29]~feeder (
// Equation(s):
// \plif_memwb.porto_l[29]~feeder_combout  = plif_exmemporto_l_29

	.dataa(gnd),
	.datab(gnd),
	.datac(plif_exmemporto_l_29),
	.datad(gnd),
	.cin(gnd),
	.combout(\plif_memwb.porto_l[29]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \plif_memwb.porto_l[29]~feeder .lut_mask = 16'hF0F0;
defparam \plif_memwb.porto_l[29]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y35_N18
cycloneive_lcell_comb \plif_memwb.porto_l[28]~feeder (
// Equation(s):
// \plif_memwb.porto_l[28]~feeder_combout  = plif_exmemporto_l_28

	.dataa(gnd),
	.datab(gnd),
	.datac(plif_exmemporto_l_28),
	.datad(gnd),
	.cin(gnd),
	.combout(\plif_memwb.porto_l[28]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \plif_memwb.porto_l[28]~feeder .lut_mask = 16'hF0F0;
defparam \plif_memwb.porto_l[28]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y35_N16
cycloneive_lcell_comb \plif_memwb.rtnaddr_l[28]~feeder (
// Equation(s):
// \plif_memwb.rtnaddr_l[28]~feeder_combout  = plif_exmemrtnaddr_l_28

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(plif_exmemrtnaddr_l_28),
	.cin(gnd),
	.combout(\plif_memwb.rtnaddr_l[28]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \plif_memwb.rtnaddr_l[28]~feeder .lut_mask = 16'hFF00;
defparam \plif_memwb.rtnaddr_l[28]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y36_N30
cycloneive_lcell_comb \plif_memwb.porto_l[27]~feeder (
// Equation(s):
// \plif_memwb.porto_l[27]~feeder_combout  = plif_exmemporto_l_27

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(plif_exmemporto_l_27),
	.cin(gnd),
	.combout(\plif_memwb.porto_l[27]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \plif_memwb.porto_l[27]~feeder .lut_mask = 16'hFF00;
defparam \plif_memwb.porto_l[27]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y35_N28
cycloneive_lcell_comb \plif_memwb.porto_l[24]~feeder (
// Equation(s):
// \plif_memwb.porto_l[24]~feeder_combout  = plif_exmemporto_l_24

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(plif_exmemporto_l_24),
	.cin(gnd),
	.combout(\plif_memwb.porto_l[24]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \plif_memwb.porto_l[24]~feeder .lut_mask = 16'hFF00;
defparam \plif_memwb.porto_l[24]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y35_N22
cycloneive_lcell_comb \plif_memwb.porto_l[23]~feeder (
// Equation(s):
// \plif_memwb.porto_l[23]~feeder_combout  = plif_exmemporto_l_23

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(plif_exmemporto_l_23),
	.cin(gnd),
	.combout(\plif_memwb.porto_l[23]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \plif_memwb.porto_l[23]~feeder .lut_mask = 16'hFF00;
defparam \plif_memwb.porto_l[23]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X52_Y39_N8
cycloneive_lcell_comb \plif_memwb.rtnaddr_l[23]~feeder (
// Equation(s):
// \plif_memwb.rtnaddr_l[23]~feeder_combout  = plif_exmemrtnaddr_l_23

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(plif_exmemrtnaddr_l_23),
	.cin(gnd),
	.combout(\plif_memwb.rtnaddr_l[23]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \plif_memwb.rtnaddr_l[23]~feeder .lut_mask = 16'hFF00;
defparam \plif_memwb.rtnaddr_l[23]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y39_N8
cycloneive_lcell_comb \plif_memwb.rtnaddr_l[22]~feeder (
// Equation(s):
// \plif_memwb.rtnaddr_l[22]~feeder_combout  = plif_exmemrtnaddr_l_22

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(plif_exmemrtnaddr_l_22),
	.cin(gnd),
	.combout(\plif_memwb.rtnaddr_l[22]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \plif_memwb.rtnaddr_l[22]~feeder .lut_mask = 16'hFF00;
defparam \plif_memwb.rtnaddr_l[22]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y35_N22
cycloneive_lcell_comb \plif_memwb.porto_l[21]~feeder (
// Equation(s):
// \plif_memwb.porto_l[21]~feeder_combout  = plif_exmemporto_l_21

	.dataa(gnd),
	.datab(gnd),
	.datac(plif_exmemporto_l_21),
	.datad(gnd),
	.cin(gnd),
	.combout(\plif_memwb.porto_l[21]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \plif_memwb.porto_l[21]~feeder .lut_mask = 16'hF0F0;
defparam \plif_memwb.porto_l[21]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y34_N14
cycloneive_lcell_comb \plif_memwb.porto_l[19]~feeder (
// Equation(s):
// \plif_memwb.porto_l[19]~feeder_combout  = plif_exmemporto_l_19

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(plif_exmemporto_l_19),
	.cin(gnd),
	.combout(\plif_memwb.porto_l[19]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \plif_memwb.porto_l[19]~feeder .lut_mask = 16'hFF00;
defparam \plif_memwb.porto_l[19]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y35_N8
cycloneive_lcell_comb \plif_memwb.rtnaddr_l[16]~feeder (
// Equation(s):
// \plif_memwb.rtnaddr_l[16]~feeder_combout  = plif_exmemrtnaddr_l_16

	.dataa(gnd),
	.datab(gnd),
	.datac(plif_exmemrtnaddr_l_16),
	.datad(gnd),
	.cin(gnd),
	.combout(\plif_memwb.rtnaddr_l[16]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \plif_memwb.rtnaddr_l[16]~feeder .lut_mask = 16'hF0F0;
defparam \plif_memwb.rtnaddr_l[16]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y34_N8
cycloneive_lcell_comb \plif_memwb.porto_l[10]~feeder (
// Equation(s):
// \plif_memwb.porto_l[10]~feeder_combout  = plif_exmemporto_l_10

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(plif_exmemporto_l_10),
	.cin(gnd),
	.combout(\plif_memwb.porto_l[10]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \plif_memwb.porto_l[10]~feeder .lut_mask = 16'hFF00;
defparam \plif_memwb.porto_l[10]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y35_N12
cycloneive_lcell_comb \plif_memwb.porto_l[9]~feeder (
// Equation(s):
// \plif_memwb.porto_l[9]~feeder_combout  = plif_exmemporto_l_9

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(plif_exmemporto_l_9),
	.cin(gnd),
	.combout(\plif_memwb.porto_l[9]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \plif_memwb.porto_l[9]~feeder .lut_mask = 16'hFF00;
defparam \plif_memwb.porto_l[9]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y35_N26
cycloneive_lcell_comb \plif_memwb.rtnaddr_l[9]~feeder (
// Equation(s):
// \plif_memwb.rtnaddr_l[9]~feeder_combout  = plif_exmemrtnaddr_l_9

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(plif_exmemrtnaddr_l_9),
	.cin(gnd),
	.combout(\plif_memwb.rtnaddr_l[9]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \plif_memwb.rtnaddr_l[9]~feeder .lut_mask = 16'hFF00;
defparam \plif_memwb.rtnaddr_l[9]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y33_N8
cycloneive_lcell_comb \plif_memwb.porto_l[8]~feeder (
// Equation(s):
// \plif_memwb.porto_l[8]~feeder_combout  = plif_exmemporto_l_8

	.dataa(gnd),
	.datab(gnd),
	.datac(plif_exmemporto_l_8),
	.datad(gnd),
	.cin(gnd),
	.combout(\plif_memwb.porto_l[8]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \plif_memwb.porto_l[8]~feeder .lut_mask = 16'hF0F0;
defparam \plif_memwb.porto_l[8]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y39_N14
cycloneive_lcell_comb \plif_memwb.rtnaddr_l[2]~feeder (
// Equation(s):
// \plif_memwb.rtnaddr_l[2]~feeder_combout  = plif_exmemrtnaddr_l_2

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(plif_exmemrtnaddr_l_2),
	.cin(gnd),
	.combout(\plif_memwb.rtnaddr_l[2]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \plif_memwb.rtnaddr_l[2]~feeder .lut_mask = 16'hFF00;
defparam \plif_memwb.rtnaddr_l[2]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y34_N22
cycloneive_lcell_comb \plif_memwb.porto_l[1]~feeder (
// Equation(s):
// \plif_memwb.porto_l[1]~feeder_combout  = plif_exmemporto_l_1

	.dataa(gnd),
	.datab(gnd),
	.datac(plif_exmemporto_l_1),
	.datad(gnd),
	.cin(gnd),
	.combout(\plif_memwb.porto_l[1]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \plif_memwb.porto_l[1]~feeder .lut_mask = 16'hF0F0;
defparam \plif_memwb.porto_l[1]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y34_N4
cycloneive_lcell_comb \plif_memwb.rtnaddr_l[1]~feeder (
// Equation(s):
// \plif_memwb.rtnaddr_l[1]~feeder_combout  = plif_exmemrtnaddr_l_1

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(plif_exmemrtnaddr_l_1),
	.cin(gnd),
	.combout(\plif_memwb.rtnaddr_l[1]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \plif_memwb.rtnaddr_l[1]~feeder .lut_mask = 16'hFF00;
defparam \plif_memwb.rtnaddr_l[1]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y33_N26
cycloneive_lcell_comb \plif_memwb.porto_l[0]~feeder (
// Equation(s):
// \plif_memwb.porto_l[0]~feeder_combout  = plif_exmemporto_l_0

	.dataa(gnd),
	.datab(gnd),
	.datac(plif_exmemporto_l_0),
	.datad(gnd),
	.cin(gnd),
	.combout(\plif_memwb.porto_l[0]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \plif_memwb.porto_l[0]~feeder .lut_mask = 16'hF0F0;
defparam \plif_memwb.porto_l[0]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y33_N0
cycloneive_lcell_comb \plif_memwb.rtnaddr_l[0]~feeder (
// Equation(s):
// \plif_memwb.rtnaddr_l[0]~feeder_combout  = plif_exmemrtnaddr_l_0

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(plif_exmemrtnaddr_l_0),
	.cin(gnd),
	.combout(\plif_memwb.rtnaddr_l[0]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \plif_memwb.rtnaddr_l[0]~feeder .lut_mask = 16'hFF00;
defparam \plif_memwb.rtnaddr_l[0]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y33_N18
cycloneive_lcell_comb \plif_memwb.porto_l[4]~feeder (
// Equation(s):
// \plif_memwb.porto_l[4]~feeder_combout  = plif_exmemporto_l_4

	.dataa(gnd),
	.datab(gnd),
	.datac(plif_exmemporto_l_4),
	.datad(gnd),
	.cin(gnd),
	.combout(\plif_memwb.porto_l[4]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \plif_memwb.porto_l[4]~feeder .lut_mask = 16'hF0F0;
defparam \plif_memwb.porto_l[4]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y33_N24
cycloneive_lcell_comb \plif_memwb.rtnaddr_l[4]~feeder (
// Equation(s):
// \plif_memwb.rtnaddr_l[4]~feeder_combout  = plif_exmemrtnaddr_l_4

	.dataa(gnd),
	.datab(gnd),
	.datac(plif_exmemrtnaddr_l_4),
	.datad(gnd),
	.cin(gnd),
	.combout(\plif_memwb.rtnaddr_l[4]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \plif_memwb.rtnaddr_l[4]~feeder .lut_mask = 16'hF0F0;
defparam \plif_memwb.rtnaddr_l[4]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y35_N10
cycloneive_lcell_comb \plif_memwb.porto_l[3]~feeder (
// Equation(s):
// \plif_memwb.porto_l[3]~feeder_combout  = plif_exmemporto_l_3

	.dataa(gnd),
	.datab(gnd),
	.datac(plif_exmemporto_l_3),
	.datad(gnd),
	.cin(gnd),
	.combout(\plif_memwb.porto_l[3]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \plif_memwb.porto_l[3]~feeder .lut_mask = 16'hF0F0;
defparam \plif_memwb.porto_l[3]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y35_N12
cycloneive_lcell_comb \plif_memwb.rtnaddr_l[3]~feeder (
// Equation(s):
// \plif_memwb.rtnaddr_l[3]~feeder_combout  = plif_exmemrtnaddr_l_3

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(plif_exmemrtnaddr_l_3),
	.cin(gnd),
	.combout(\plif_memwb.rtnaddr_l[3]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \plif_memwb.rtnaddr_l[3]~feeder .lut_mask = 16'hFF00;
defparam \plif_memwb.rtnaddr_l[3]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y32_N12
cycloneive_lcell_comb \plif_memwb.btype_l~feeder (
// Equation(s):
// \plif_memwb.btype_l~feeder_combout  = plif_exmembtype_l

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(plif_exmembtype_l),
	.cin(gnd),
	.combout(\plif_memwb.btype_l~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \plif_memwb.btype_l~feeder .lut_mask = 16'hFF00;
defparam \plif_memwb.btype_l~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y29_N16
cycloneive_lcell_comb \plif_memwb.jaddr_l[1]~feeder (
// Equation(s):
// \plif_memwb.jaddr_l[1]~feeder_combout  = plif_exmemjaddr_l_1

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(plif_exmemjaddr_l_1),
	.cin(gnd),
	.combout(\plif_memwb.jaddr_l[1]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \plif_memwb.jaddr_l[1]~feeder .lut_mask = 16'hFF00;
defparam \plif_memwb.jaddr_l[1]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y29_N22
cycloneive_lcell_comb \plif_memwb.extimm_l[0]~feeder (
// Equation(s):
// \plif_memwb.extimm_l[0]~feeder_combout  = plif_exmemextimm_l_0

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(plif_exmemextimm_l_0),
	.cin(gnd),
	.combout(\plif_memwb.extimm_l[0]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \plif_memwb.extimm_l[0]~feeder .lut_mask = 16'hFF00;
defparam \plif_memwb.extimm_l[0]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y29_N0
cycloneive_lcell_comb \plif_memwb.jaddr_l[5]~feeder (
// Equation(s):
// \plif_memwb.jaddr_l[5]~feeder_combout  = plif_exmemjaddr_l_5

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(plif_exmemjaddr_l_5),
	.cin(gnd),
	.combout(\plif_memwb.jaddr_l[5]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \plif_memwb.jaddr_l[5]~feeder .lut_mask = 16'hFF00;
defparam \plif_memwb.jaddr_l[5]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y29_N10
cycloneive_lcell_comb \plif_memwb.extimm_l[7]~feeder (
// Equation(s):
// \plif_memwb.extimm_l[7]~feeder_combout  = plif_exmemextimm_l_7

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(plif_exmemextimm_l_7),
	.cin(gnd),
	.combout(\plif_memwb.extimm_l[7]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \plif_memwb.extimm_l[7]~feeder .lut_mask = 16'hFF00;
defparam \plif_memwb.extimm_l[7]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y32_N12
cycloneive_lcell_comb \plif_memwb.jaddr_l[9]~feeder (
// Equation(s):
// \plif_memwb.jaddr_l[9]~feeder_combout  = plif_exmemjaddr_l_9

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(plif_exmemjaddr_l_9),
	.cin(gnd),
	.combout(\plif_memwb.jaddr_l[9]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \plif_memwb.jaddr_l[9]~feeder .lut_mask = 16'hFF00;
defparam \plif_memwb.jaddr_l[9]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y32_N8
cycloneive_lcell_comb \plif_memwb.extimm_l[8]~feeder (
// Equation(s):
// \plif_memwb.extimm_l[8]~feeder_combout  = plif_exmemextimm_l_8

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(plif_exmemextimm_l_8),
	.cin(gnd),
	.combout(\plif_memwb.extimm_l[8]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \plif_memwb.extimm_l[8]~feeder .lut_mask = 16'hFF00;
defparam \plif_memwb.extimm_l[8]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y32_N6
cycloneive_lcell_comb \plif_memwb.jaddr_l[11]~feeder (
// Equation(s):
// \plif_memwb.jaddr_l[11]~feeder_combout  = plif_exmemjaddr_l_11

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(plif_exmemjaddr_l_11),
	.cin(gnd),
	.combout(\plif_memwb.jaddr_l[11]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \plif_memwb.jaddr_l[11]~feeder .lut_mask = 16'hFF00;
defparam \plif_memwb.jaddr_l[11]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y32_N16
cycloneive_lcell_comb \plif_memwb.extimm_l[11]~feeder (
// Equation(s):
// \plif_memwb.extimm_l[11]~feeder_combout  = plif_exmemextimm_l_11

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(plif_exmemextimm_l_11),
	.cin(gnd),
	.combout(\plif_memwb.extimm_l[11]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \plif_memwb.extimm_l[11]~feeder .lut_mask = 16'hFF00;
defparam \plif_memwb.extimm_l[11]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y31_N12
cycloneive_lcell_comb \plif_memwb.extimm_l[12]~feeder (
// Equation(s):
// \plif_memwb.extimm_l[12]~feeder_combout  = plif_exmemextimm_l_12

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(plif_exmemextimm_l_12),
	.cin(gnd),
	.combout(\plif_memwb.extimm_l[12]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \plif_memwb.extimm_l[12]~feeder .lut_mask = 16'hFF00;
defparam \plif_memwb.extimm_l[12]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y31_N26
cycloneive_lcell_comb \plif_memwb.jaddr_l[15]~feeder (
// Equation(s):
// \plif_memwb.jaddr_l[15]~feeder_combout  = plif_exmemjaddr_l_15

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(plif_exmemjaddr_l_15),
	.cin(gnd),
	.combout(\plif_memwb.jaddr_l[15]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \plif_memwb.jaddr_l[15]~feeder .lut_mask = 16'hFF00;
defparam \plif_memwb.jaddr_l[15]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y31_N20
cycloneive_lcell_comb \plif_memwb.extimm_l[15]~feeder (
// Equation(s):
// \plif_memwb.extimm_l[15]~feeder_combout  = plif_exmemextimm_l_15

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(plif_exmemextimm_l_15),
	.cin(gnd),
	.combout(\plif_memwb.extimm_l[15]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \plif_memwb.extimm_l[15]~feeder .lut_mask = 16'hFF00;
defparam \plif_memwb.extimm_l[15]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y31_N6
cycloneive_lcell_comb \plif_memwb.extimm_l[14]~feeder (
// Equation(s):
// \plif_memwb.extimm_l[14]~feeder_combout  = plif_exmemextimm_l_14

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(plif_exmemextimm_l_14),
	.cin(gnd),
	.combout(\plif_memwb.extimm_l[14]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \plif_memwb.extimm_l[14]~feeder .lut_mask = 16'hFF00;
defparam \plif_memwb.extimm_l[14]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y32_N0
cycloneive_lcell_comb \plif_memwb.jaddr_l[17]~feeder (
// Equation(s):
// \plif_memwb.jaddr_l[17]~feeder_combout  = plif_exmemjaddr_l_17

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(plif_exmemjaddr_l_17),
	.cin(gnd),
	.combout(\plif_memwb.jaddr_l[17]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \plif_memwb.jaddr_l[17]~feeder .lut_mask = 16'hFF00;
defparam \plif_memwb.jaddr_l[17]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y31_N28
cycloneive_lcell_comb \plif_memwb.extimm_l[17]~feeder (
// Equation(s):
// \plif_memwb.extimm_l[17]~feeder_combout  = plif_exmemextimm_l_17

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(plif_exmemextimm_l_17),
	.cin(gnd),
	.combout(\plif_memwb.extimm_l[17]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \plif_memwb.extimm_l[17]~feeder .lut_mask = 16'hFF00;
defparam \plif_memwb.extimm_l[17]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y33_N8
cycloneive_lcell_comb \plif_memwb.jaddr_l[19]~feeder (
// Equation(s):
// \plif_memwb.jaddr_l[19]~feeder_combout  = plif_exmemjaddr_l_19

	.dataa(gnd),
	.datab(gnd),
	.datac(plif_exmemjaddr_l_19),
	.datad(gnd),
	.cin(gnd),
	.combout(\plif_memwb.jaddr_l[19]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \plif_memwb.jaddr_l[19]~feeder .lut_mask = 16'hF0F0;
defparam \plif_memwb.jaddr_l[19]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y31_N14
cycloneive_lcell_comb \plif_memwb.extimm_l[18]~feeder (
// Equation(s):
// \plif_memwb.extimm_l[18]~feeder_combout  = plif_exmemextimm_l_18

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(plif_exmemextimm_l_18),
	.cin(gnd),
	.combout(\plif_memwb.extimm_l[18]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \plif_memwb.extimm_l[18]~feeder .lut_mask = 16'hFF00;
defparam \plif_memwb.extimm_l[18]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y31_N0
cycloneive_lcell_comb \plif_memwb.jaddr_l[21]~feeder (
// Equation(s):
// \plif_memwb.jaddr_l[21]~feeder_combout  = plif_exmemjaddr_l_21

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(plif_exmemjaddr_l_21),
	.cin(gnd),
	.combout(\plif_memwb.jaddr_l[21]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \plif_memwb.jaddr_l[21]~feeder .lut_mask = 16'hFF00;
defparam \plif_memwb.jaddr_l[21]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y31_N24
cycloneive_lcell_comb \plif_memwb.extimm_l[23]~feeder (
// Equation(s):
// \plif_memwb.extimm_l[23]~feeder_combout  = plif_exmemextimm_l_23

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(plif_exmemextimm_l_23),
	.cin(gnd),
	.combout(\plif_memwb.extimm_l[23]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \plif_memwb.extimm_l[23]~feeder .lut_mask = 16'hFF00;
defparam \plif_memwb.extimm_l[23]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y31_N6
cycloneive_lcell_comb \plif_memwb.jaddr_l[25]~feeder (
// Equation(s):
// \plif_memwb.jaddr_l[25]~feeder_combout  = plif_exmemjaddr_l_25

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(plif_exmemjaddr_l_25),
	.cin(gnd),
	.combout(\plif_memwb.jaddr_l[25]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \plif_memwb.jaddr_l[25]~feeder .lut_mask = 16'hFF00;
defparam \plif_memwb.jaddr_l[25]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y28_N4
cycloneive_lcell_comb \plif_memwb.extimm_l[24]~feeder (
// Equation(s):
// \plif_memwb.extimm_l[24]~feeder_combout  = plif_exmemextimm_l_24

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(plif_exmemextimm_l_24),
	.cin(gnd),
	.combout(\plif_memwb.extimm_l[24]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \plif_memwb.extimm_l[24]~feeder .lut_mask = 16'hFF00;
defparam \plif_memwb.extimm_l[24]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y31_N8
cycloneive_lcell_comb \plif_memwb.extimm_l[28]~feeder (
// Equation(s):
// \plif_memwb.extimm_l[28]~feeder_combout  = plif_exmemextimm_l_28

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(plif_exmemextimm_l_28),
	.cin(gnd),
	.combout(\plif_memwb.extimm_l[28]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \plif_memwb.extimm_l[28]~feeder .lut_mask = 16'hFF00;
defparam \plif_memwb.extimm_l[28]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

endmodule

module register_file (
	plif_memwbregsrc_l_1,
	wdat_31,
	plif_memwbrtnaddr_l_31,
	plif_memwbwsel_l_4,
	plif_memwbwsel_l_3,
	plif_memwbwsel_l_0,
	plif_memwbwsel_l_2,
	plif_memwbwsel_l_1,
	Decoder0,
	WideOr0,
	plif_memwbregen_l,
	wdat_30,
	plif_memwbrtnaddr_l_30,
	wdat_29,
	plif_memwbrtnaddr_l_29,
	wdat_28,
	plif_memwbrtnaddr_l_28,
	wdat_27,
	plif_memwbrtnaddr_l_27,
	wdat_26,
	plif_memwbrtnaddr_l_26,
	wdat_25,
	plif_memwbrtnaddr_l_25,
	wdat_24,
	plif_memwbrtnaddr_l_24,
	wdat_23,
	plif_memwbrtnaddr_l_23,
	wdat_22,
	plif_memwbrtnaddr_l_22,
	wdat_21,
	plif_memwbrtnaddr_l_21,
	wdat_20,
	plif_memwbrtnaddr_l_20,
	wdat_19,
	plif_memwbrtnaddr_l_19,
	wdat_18,
	plif_memwbrtnaddr_l_18,
	wdat_17,
	plif_memwbrtnaddr_l_17,
	wdat_16,
	plif_memwbrtnaddr_l_16,
	wdat_15,
	plif_memwbrtnaddr_l_15,
	wdat_14,
	plif_memwbrtnaddr_l_14,
	wdat_13,
	plif_memwbrtnaddr_l_13,
	wdat_12,
	plif_memwbrtnaddr_l_12,
	wdat_11,
	plif_memwbrtnaddr_l_11,
	wdat_10,
	plif_memwbrtnaddr_l_10,
	wdat_9,
	plif_memwbrtnaddr_l_9,
	wdat_8,
	plif_memwbrtnaddr_l_8,
	wdat_7,
	plif_memwbrtnaddr_l_7,
	wdat_6,
	plif_memwbrtnaddr_l_6,
	wdat_5,
	plif_memwbrtnaddr_l_5,
	wdat_2,
	plif_memwbrtnaddr_l_2,
	wdat_1,
	plif_memwbrtnaddr_l_1,
	wdat_0,
	plif_memwbrtnaddr_l_0,
	wdat_4,
	plif_memwbrtnaddr_l_4,
	wdat_3,
	plif_memwbrtnaddr_l_3,
	Selector4,
	plif_ifidinstr_l_22,
	Selector41,
	Selector5,
	Selector2,
	Selector3,
	Selector9,
	plif_ifidinstr_l_17,
	Selector91,
	Selector10,
	Selector7,
	Selector8,
	Mux32,
	Mux321,
	Mux33,
	Mux331,
	Mux34,
	Mux341,
	Mux35,
	Mux351,
	Mux36,
	Mux361,
	Mux37,
	Mux371,
	Mux38,
	Mux381,
	Mux39,
	Mux391,
	Mux40,
	Mux401,
	Mux41,
	Mux411,
	Mux42,
	Mux421,
	Mux43,
	Mux431,
	Mux44,
	Mux441,
	Mux45,
	Mux451,
	Mux46,
	Mux461,
	Mux47,
	Mux471,
	Mux48,
	Mux481,
	Mux49,
	Mux491,
	Mux50,
	Mux501,
	Mux51,
	Mux511,
	Mux52,
	Mux521,
	Mux53,
	Mux531,
	Mux54,
	Mux541,
	Mux55,
	Mux551,
	Mux56,
	Mux561,
	Mux57,
	Mux571,
	Mux58,
	Mux581,
	Mux29,
	Mux291,
	Mux30,
	Mux301,
	Mux63,
	Mux631,
	Mux62,
	Mux621,
	Mux27,
	Mux271,
	Mux28,
	Mux281,
	Mux61,
	Mux611,
	Mux23,
	Mux231,
	Mux24,
	Mux241,
	Mux25,
	Mux251,
	Mux26,
	Mux261,
	Mux60,
	Mux601,
	Mux15,
	Mux151,
	Mux16,
	Mux161,
	Mux17,
	Mux171,
	Mux18,
	Mux181,
	Mux19,
	Mux191,
	Mux20,
	Mux201,
	Mux21,
	Mux211,
	Mux22,
	Mux221,
	Mux59,
	Mux591,
	Mux0,
	Mux01,
	Mux2,
	Mux210,
	Mux1,
	Mux11,
	Mux3,
	Mux31,
	Mux4,
	Mux410,
	Mux5,
	Mux510,
	Mux6,
	Mux64,
	Mux7,
	Mux71,
	Mux8,
	Mux81,
	Mux9,
	Mux91,
	Mux10,
	Mux101,
	Mux111,
	Mux112,
	Mux12,
	Mux121,
	Mux13,
	Mux131,
	Mux14,
	Mux141,
	Mux311,
	Mux312,
	CLK,
	nRST,
	devpor,
	devclrn,
	devoe);
input 	plif_memwbregsrc_l_1;
input 	wdat_31;
input 	plif_memwbrtnaddr_l_31;
input 	plif_memwbwsel_l_4;
input 	plif_memwbwsel_l_3;
input 	plif_memwbwsel_l_0;
input 	plif_memwbwsel_l_2;
input 	plif_memwbwsel_l_1;
output 	Decoder0;
input 	WideOr0;
input 	plif_memwbregen_l;
input 	wdat_30;
input 	plif_memwbrtnaddr_l_30;
input 	wdat_29;
input 	plif_memwbrtnaddr_l_29;
input 	wdat_28;
input 	plif_memwbrtnaddr_l_28;
input 	wdat_27;
input 	plif_memwbrtnaddr_l_27;
input 	wdat_26;
input 	plif_memwbrtnaddr_l_26;
input 	wdat_25;
input 	plif_memwbrtnaddr_l_25;
input 	wdat_24;
input 	plif_memwbrtnaddr_l_24;
input 	wdat_23;
input 	plif_memwbrtnaddr_l_23;
input 	wdat_22;
input 	plif_memwbrtnaddr_l_22;
input 	wdat_21;
input 	plif_memwbrtnaddr_l_21;
input 	wdat_20;
input 	plif_memwbrtnaddr_l_20;
input 	wdat_19;
input 	plif_memwbrtnaddr_l_19;
input 	wdat_18;
input 	plif_memwbrtnaddr_l_18;
input 	wdat_17;
input 	plif_memwbrtnaddr_l_17;
input 	wdat_16;
input 	plif_memwbrtnaddr_l_16;
input 	wdat_15;
input 	plif_memwbrtnaddr_l_15;
input 	wdat_14;
input 	plif_memwbrtnaddr_l_14;
input 	wdat_13;
input 	plif_memwbrtnaddr_l_13;
input 	wdat_12;
input 	plif_memwbrtnaddr_l_12;
input 	wdat_11;
input 	plif_memwbrtnaddr_l_11;
input 	wdat_10;
input 	plif_memwbrtnaddr_l_10;
input 	wdat_9;
input 	plif_memwbrtnaddr_l_9;
input 	wdat_8;
input 	plif_memwbrtnaddr_l_8;
input 	wdat_7;
input 	plif_memwbrtnaddr_l_7;
input 	wdat_6;
input 	plif_memwbrtnaddr_l_6;
input 	wdat_5;
input 	plif_memwbrtnaddr_l_5;
input 	wdat_2;
input 	plif_memwbrtnaddr_l_2;
input 	wdat_1;
input 	plif_memwbrtnaddr_l_1;
input 	wdat_0;
input 	plif_memwbrtnaddr_l_0;
input 	wdat_4;
input 	plif_memwbrtnaddr_l_4;
input 	wdat_3;
input 	plif_memwbrtnaddr_l_3;
input 	Selector4;
input 	plif_ifidinstr_l_22;
input 	Selector41;
input 	Selector5;
input 	Selector2;
input 	Selector3;
input 	Selector9;
input 	plif_ifidinstr_l_17;
input 	Selector91;
input 	Selector10;
input 	Selector7;
input 	Selector8;
output 	Mux32;
output 	Mux321;
output 	Mux33;
output 	Mux331;
output 	Mux34;
output 	Mux341;
output 	Mux35;
output 	Mux351;
output 	Mux36;
output 	Mux361;
output 	Mux37;
output 	Mux371;
output 	Mux38;
output 	Mux381;
output 	Mux39;
output 	Mux391;
output 	Mux40;
output 	Mux401;
output 	Mux41;
output 	Mux411;
output 	Mux42;
output 	Mux421;
output 	Mux43;
output 	Mux431;
output 	Mux44;
output 	Mux441;
output 	Mux45;
output 	Mux451;
output 	Mux46;
output 	Mux461;
output 	Mux47;
output 	Mux471;
output 	Mux48;
output 	Mux481;
output 	Mux49;
output 	Mux491;
output 	Mux50;
output 	Mux501;
output 	Mux51;
output 	Mux511;
output 	Mux52;
output 	Mux521;
output 	Mux53;
output 	Mux531;
output 	Mux54;
output 	Mux541;
output 	Mux55;
output 	Mux551;
output 	Mux56;
output 	Mux561;
output 	Mux57;
output 	Mux571;
output 	Mux58;
output 	Mux581;
output 	Mux29;
output 	Mux291;
output 	Mux30;
output 	Mux301;
output 	Mux63;
output 	Mux631;
output 	Mux62;
output 	Mux621;
output 	Mux27;
output 	Mux271;
output 	Mux28;
output 	Mux281;
output 	Mux61;
output 	Mux611;
output 	Mux23;
output 	Mux231;
output 	Mux24;
output 	Mux241;
output 	Mux25;
output 	Mux251;
output 	Mux26;
output 	Mux261;
output 	Mux60;
output 	Mux601;
output 	Mux15;
output 	Mux151;
output 	Mux16;
output 	Mux161;
output 	Mux17;
output 	Mux171;
output 	Mux18;
output 	Mux181;
output 	Mux19;
output 	Mux191;
output 	Mux20;
output 	Mux201;
output 	Mux21;
output 	Mux211;
output 	Mux22;
output 	Mux221;
output 	Mux59;
output 	Mux591;
output 	Mux0;
output 	Mux01;
output 	Mux2;
output 	Mux210;
output 	Mux1;
output 	Mux11;
output 	Mux3;
output 	Mux31;
output 	Mux4;
output 	Mux410;
output 	Mux5;
output 	Mux510;
output 	Mux6;
output 	Mux64;
output 	Mux7;
output 	Mux71;
output 	Mux8;
output 	Mux81;
output 	Mux9;
output 	Mux91;
output 	Mux10;
output 	Mux101;
output 	Mux111;
output 	Mux112;
output 	Mux12;
output 	Mux121;
output 	Mux13;
output 	Mux131;
output 	Mux14;
output 	Mux141;
output 	Mux311;
output 	Mux312;
input 	CLK;
input 	nRST;

// Design Ports Information

input 	devpor;
input 	devclrn;
input 	devoe;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
assign unknown = 1'bx;

wire \register[28][30]~q ;
wire \register[3][29]~q ;
wire \Mux34~14_combout ;
wire \register[30][28]~q ;
wire \register[24][28]~q ;
wire \Mux35~4_combout ;
wire \register[3][28]~q ;
wire \register[1][28]~q ;
wire \Mux35~14_combout ;
wire \register[4][24]~q ;
wire \Mux39~12_combout ;
wire \register[1][23]~q ;
wire \Mux40~14_combout ;
wire \register[28][21]~q ;
wire \register[5][21]~q ;
wire \register[8][21]~q ;
wire \Mux42~12_combout ;
wire \register[26][20]~q ;
wire \Mux43~2_combout ;
wire \register[24][20]~q ;
wire \Mux43~4_combout ;
wire \register[4][19]~q ;
wire \register[13][19]~q ;
wire \register[8][18]~q ;
wire \Mux45~12_combout ;
wire \register[13][18]~q ;
wire \register[28][17]~q ;
wire \register[8][17]~q ;
wire \Mux46~12_combout ;
wire \register[18][16]~q ;
wire \Mux47~2_combout ;
wire \Mux48~12_combout ;
wire \register[22][13]~q ;
wire \register[22][12]~q ;
wire \register[10][10]~q ;
wire \register[26][8]~q ;
wire \Mux55~2_combout ;
wire \register[20][8]~q ;
wire \Mux56~12_combout ;
wire \register[18][6]~q ;
wire \Mux57~2_combout ;
wire \register[16][5]~q ;
wire \register[28][5]~q ;
wire \Mux58~12_combout ;
wire \register[3][2]~q ;
wire \register[1][2]~q ;
wire \Mux29~14_combout ;
wire \register[24][1]~q ;
wire \register[20][0]~q ;
wire \register[8][0]~q ;
wire \register[28][4]~q ;
wire \register[3][4]~q ;
wire \Mux61~14_combout ;
wire \Mux24~4_combout ;
wire \Mux25~2_combout ;
wire \Mux60~14_combout ;
wire \Mux15~4_combout ;
wire \Mux16~14_combout ;
wire \Mux17~14_combout ;
wire \Mux19~2_combout ;
wire \Mux21~12_combout ;
wire \Mux22~2_combout ;
wire \Mux59~14_combout ;
wire \Mux2~2_combout ;
wire \Mux2~12_combout ;
wire \Mux3~14_combout ;
wire \Mux6~14_combout ;
wire \Mux9~12_combout ;
wire \Mux9~14_combout ;
wire \Mux10~12_combout ;
wire \Mux12~12_combout ;
wire \Mux13~4_combout ;
wire \Mux13~12_combout ;
wire \Mux31~12_combout ;
wire \register[28][30]~feeder_combout ;
wire \register[30][28]~feeder_combout ;
wire \register[24][28]~feeder_combout ;
wire \register[28][21]~feeder_combout ;
wire \register[24][20]~feeder_combout ;
wire \register[13][19]~feeder_combout ;
wire \register[13][18]~feeder_combout ;
wire \register[28][17]~feeder_combout ;
wire \register[22][13]~feeder_combout ;
wire \register[20][8]~feeder_combout ;
wire \register[18][6]~feeder_combout ;
wire \register[28][5]~feeder_combout ;
wire \register[16][5]~feeder_combout ;
wire \register[24][1]~feeder_combout ;
wire \register[8][0]~feeder_combout ;
wire \register[20][0]~feeder_combout ;
wire \register[28][4]~feeder_combout ;
wire \register~64_combout ;
wire \Decoder0~32_combout ;
wire \Decoder0~37_combout ;
wire \register[23][31]~q ;
wire \Decoder0~40_combout ;
wire \register[31][31]~q ;
wire \register[27][31]~feeder_combout ;
wire \Decoder0~29_combout ;
wire \Decoder0~38_combout ;
wire \register[27][31]~q ;
wire \Decoder0~39_combout ;
wire \register[19][31]~q ;
wire \Mux32~7_combout ;
wire \Mux32~8_combout ;
wire \register[29][31]~feeder_combout ;
wire \Decoder0~27_combout ;
wire \Decoder0~28_combout ;
wire \register[29][31]~q ;
wire \Decoder0~21_combout ;
wire \Decoder0~22_combout ;
wire \register[21][31]~q ;
wire \register[25][31]~feeder_combout ;
wire \Decoder0~23_combout ;
wire \Decoder0~24_combout ;
wire \register[25][31]~q ;
wire \Mux32~0_combout ;
wire \Mux32~1_combout ;
wire \Decoder0~34_combout ;
wire \register[24][31]~q ;
wire \Decoder0~25_combout ;
wire \Decoder0~36_combout ;
wire \register[16][31]~q ;
wire \Mux32~4_combout ;
wire \register[28][31]~feeder_combout ;
wire \Decoder0~57_combout ;
wire \register[28][31]~q ;
wire \Mux32~5_combout ;
wire \register[26][31]~feeder_combout ;
wire \Decoder0~30_combout ;
wire \Decoder0~54_combout ;
wire \register[26][31]~q ;
wire \Decoder0~33_combout ;
wire \register[18][31]~q ;
wire \Decoder0~55_combout ;
wire \register[22][31]~q ;
wire \Mux32~2_combout ;
wire \register[30][31]~feeder_combout ;
wire \Decoder0~56_combout ;
wire \register[30][31]~q ;
wire \Mux32~3_combout ;
wire \Mux32~6_combout ;
wire \Decoder0~41_combout ;
wire \Decoder0~43_combout ;
wire \register[7][31]~q ;
wire \Decoder0~58_combout ;
wire \register[6][31]~q ;
wire \Decoder0~59_combout ;
wire \register[5][31]~q ;
wire \Mux32~10_combout ;
wire \Mux32~11_combout ;
wire \register[14][31]~feeder_combout ;
wire \Decoder0~61_combout ;
wire \register[14][31]~q ;
wire \Decoder0~51_combout ;
wire \Decoder0~62_combout ;
wire \register[13][31]~q ;
wire \Mux32~17_combout ;
wire \register[15][31]~feeder_combout ;
wire \Decoder0~53_combout ;
wire \register[15][31]~q ;
wire \Mux32~18_combout ;
wire \Decoder0~50_combout ;
wire \register[2][31]~q ;
wire \Decoder0~48_combout ;
wire \register[3][31]~q ;
wire \Decoder0~42_combout ;
wire \Decoder0~49_combout ;
wire \register[1][31]~q ;
wire \Mux32~14_combout ;
wire \Mux32~15_combout ;
wire \Decoder0~44_combout ;
wire \register[9][31]~q ;
wire \Decoder0~46_combout ;
wire \register[8][31]~q ;
wire \Decoder0~45_combout ;
wire \register[10][31]~q ;
wire \Mux32~12_combout ;
wire \Mux32~13_combout ;
wire \Mux32~16_combout ;
wire \register~65_combout ;
wire \Decoder0~35_combout ;
wire \register[20][30]~q ;
wire \register[16][30]~q ;
wire \Mux33~4_combout ;
wire \Mux33~5_combout ;
wire \register[18][30]~q ;
wire \Mux33~2_combout ;
wire \register[30][30]~feeder_combout ;
wire \register[30][30]~q ;
wire \Mux33~3_combout ;
wire \Mux33~6_combout ;
wire \register[27][30]~q ;
wire \register[31][30]~q ;
wire \register[23][30]~feeder_combout ;
wire \register[23][30]~q ;
wire \register[19][30]~feeder_combout ;
wire \register[19][30]~q ;
wire \Mux33~7_combout ;
wire \Mux33~8_combout ;
wire \register[25][30]~feeder_combout ;
wire \register[25][30]~q ;
wire \register[21][30]~q ;
wire \Mux33~0_combout ;
wire \register[29][30]~q ;
wire \Mux33~1_combout ;
wire \register[14][30]~q ;
wire \register[15][30]~q ;
wire \register[13][30]~q ;
wire \Decoder0~31_combout ;
wire \Decoder0~52_combout ;
wire \register[12][30]~q ;
wire \Mux33~17_combout ;
wire \Mux33~18_combout ;
wire \register[10][30]~q ;
wire \register[8][30]~q ;
wire \Mux33~10_combout ;
wire \Decoder0~47_combout ;
wire \register[11][30]~q ;
wire \register[9][30]~q ;
wire \Mux33~11_combout ;
wire \register[6][30]~q ;
wire \register[7][30]~q ;
wire \register[5][30]~q ;
wire \Mux33~12_combout ;
wire \Mux33~13_combout ;
wire \register[2][30]~q ;
wire \register[3][30]~q ;
wire \register[1][30]~q ;
wire \Mux33~14_combout ;
wire \Mux33~15_combout ;
wire \Mux33~16_combout ;
wire \register~66_combout ;
wire \register[31][29]~q ;
wire \register[23][29]~q ;
wire \register[19][29]~q ;
wire \register[27][29]~q ;
wire \Mux34~7_combout ;
wire \Mux34~8_combout ;
wire \register[29][29]~feeder_combout ;
wire \register[29][29]~q ;
wire \register[21][29]~q ;
wire \register[25][29]~q ;
wire \Decoder0~26_combout ;
wire \register[17][29]~q ;
wire \Mux34~0_combout ;
wire \Mux34~1_combout ;
wire \register[22][29]~q ;
wire \register[18][29]~q ;
wire \Mux34~2_combout ;
wire \register[26][29]~q ;
wire \Mux34~3_combout ;
wire \register[28][29]~q ;
wire \register[16][29]~q ;
wire \register[20][29]~feeder_combout ;
wire \register[20][29]~q ;
wire \Mux34~4_combout ;
wire \Mux34~5_combout ;
wire \Mux34~6_combout ;
wire \register[14][29]~q ;
wire \register[15][29]~feeder_combout ;
wire \register[15][29]~q ;
wire \register[12][29]~q ;
wire \register[13][29]~feeder_combout ;
wire \register[13][29]~q ;
wire \Mux34~17_combout ;
wire \Mux34~18_combout ;
wire \register[7][29]~q ;
wire \register[6][29]~q ;
wire \Decoder0~60_combout ;
wire \register[4][29]~q ;
wire \register[5][29]~q ;
wire \Mux34~10_combout ;
wire \Mux34~11_combout ;
wire \register[2][29]~feeder_combout ;
wire \register[2][29]~q ;
wire \Mux34~15_combout ;
wire \register[9][29]~q ;
wire \register[11][29]~q ;
wire \register[10][29]~q ;
wire \Mux34~12_combout ;
wire \Mux34~13_combout ;
wire \Mux34~16_combout ;
wire \register~67_combout ;
wire \register[27][28]~feeder_combout ;
wire \register[27][28]~q ;
wire \register[31][28]~feeder_combout ;
wire \register[31][28]~q ;
wire \register[19][28]~q ;
wire \register[23][28]~q ;
wire \Mux35~7_combout ;
wire \Mux35~8_combout ;
wire \register[21][28]~feeder_combout ;
wire \register[21][28]~q ;
wire \Mux35~0_combout ;
wire \register[29][28]~feeder_combout ;
wire \register[29][28]~q ;
wire \register[25][28]~q ;
wire \Mux35~1_combout ;
wire \register[20][28]~q ;
wire \register[28][28]~feeder_combout ;
wire \register[28][28]~q ;
wire \Mux35~5_combout ;
wire \register[18][28]~q ;
wire \register[26][28]~q ;
wire \Mux35~2_combout ;
wire \register[22][28]~feeder_combout ;
wire \register[22][28]~q ;
wire \Mux35~3_combout ;
wire \Mux35~6_combout ;
wire \register[15][28]~feeder_combout ;
wire \register[15][28]~q ;
wire \register[14][28]~q ;
wire \register[12][28]~q ;
wire \Mux35~17_combout ;
wire \Mux35~18_combout ;
wire \register[2][28]~feeder_combout ;
wire \register[2][28]~q ;
wire \Mux35~15_combout ;
wire \register[7][28]~feeder_combout ;
wire \register[7][28]~q ;
wire \register[5][28]~q ;
wire \register[4][28]~q ;
wire \Mux35~12_combout ;
wire \Mux35~13_combout ;
wire \Mux35~16_combout ;
wire \register[11][28]~q ;
wire \register[9][28]~q ;
wire \register[8][28]~q ;
wire \register[10][28]~q ;
wire \Mux35~10_combout ;
wire \Mux35~11_combout ;
wire \register~68_combout ;
wire \register[23][27]~feeder_combout ;
wire \register[23][27]~q ;
wire \register[31][27]~q ;
wire \register[27][27]~q ;
wire \Mux36~7_combout ;
wire \Mux36~8_combout ;
wire \register[29][27]~feeder_combout ;
wire \register[29][27]~q ;
wire \register[17][27]~feeder_combout ;
wire \register[17][27]~q ;
wire \register[25][27]~q ;
wire \Mux36~0_combout ;
wire \register[21][27]~q ;
wire \Mux36~1_combout ;
wire \register[16][27]~q ;
wire \register[20][27]~q ;
wire \Mux36~4_combout ;
wire \register[24][27]~q ;
wire \register[28][27]~feeder_combout ;
wire \register[28][27]~q ;
wire \Mux36~5_combout ;
wire \register[30][27]~q ;
wire \register[22][27]~q ;
wire \register[18][27]~q ;
wire \Mux36~2_combout ;
wire \register[26][27]~q ;
wire \Mux36~3_combout ;
wire \Mux36~6_combout ;
wire \register[5][27]~q ;
wire \Mux36~10_combout ;
wire \register[6][27]~q ;
wire \register[7][27]~q ;
wire \Mux36~11_combout ;
wire \register[15][27]~feeder_combout ;
wire \register[15][27]~q ;
wire \register[14][27]~feeder_combout ;
wire \register[14][27]~q ;
wire \register[13][27]~q ;
wire \Mux36~17_combout ;
wire \Mux36~18_combout ;
wire \register[1][27]~q ;
wire \register[3][27]~q ;
wire \Mux36~14_combout ;
wire \Mux36~15_combout ;
wire \register[9][27]~q ;
wire \register[11][27]~q ;
wire \register[10][27]~q ;
wire \register[8][27]~q ;
wire \Mux36~12_combout ;
wire \Mux36~13_combout ;
wire \Mux36~16_combout ;
wire \register~69_combout ;
wire \register[17][26]~q ;
wire \register[21][26]~feeder_combout ;
wire \register[21][26]~q ;
wire \Mux37~0_combout ;
wire \register[29][26]~q ;
wire \register[25][26]~feeder_combout ;
wire \register[25][26]~q ;
wire \Mux37~1_combout ;
wire \register[19][26]~q ;
wire \register[23][26]~q ;
wire \Mux37~7_combout ;
wire \register[27][26]~feeder_combout ;
wire \register[27][26]~q ;
wire \register[31][26]~feeder_combout ;
wire \register[31][26]~q ;
wire \Mux37~8_combout ;
wire \register[30][26]~feeder_combout ;
wire \register[30][26]~q ;
wire \register[22][26]~q ;
wire \register[18][26]~q ;
wire \register[26][26]~q ;
wire \Mux37~2_combout ;
wire \Mux37~3_combout ;
wire \register[28][26]~feeder_combout ;
wire \register[28][26]~q ;
wire \register[20][26]~q ;
wire \register[24][26]~q ;
wire \Mux37~4_combout ;
wire \Mux37~5_combout ;
wire \Mux37~6_combout ;
wire \register[11][26]~feeder_combout ;
wire \register[11][26]~q ;
wire \register[9][26]~q ;
wire \register[10][26]~q ;
wire \register[8][26]~q ;
wire \Mux37~10_combout ;
wire \Mux37~11_combout ;
wire \register[1][26]~q ;
wire \register[3][26]~q ;
wire \Mux37~14_combout ;
wire \Mux37~15_combout ;
wire \register[5][26]~q ;
wire \register[4][26]~q ;
wire \Mux37~12_combout ;
wire \register[7][26]~q ;
wire \register[6][26]~q ;
wire \Mux37~13_combout ;
wire \Mux37~16_combout ;
wire \register[14][26]~feeder_combout ;
wire \register[14][26]~q ;
wire \register[15][26]~q ;
wire \register[13][26]~q ;
wire \register[12][26]~q ;
wire \Mux37~17_combout ;
wire \Mux37~18_combout ;
wire \register~70_combout ;
wire \register[29][25]~feeder_combout ;
wire \register[29][25]~q ;
wire \register[21][25]~q ;
wire \register[25][25]~q ;
wire \register[17][25]~q ;
wire \Mux38~0_combout ;
wire \Mux38~1_combout ;
wire \register[23][25]~feeder_combout ;
wire \register[23][25]~q ;
wire \register[31][25]~feeder_combout ;
wire \register[31][25]~q ;
wire \register[19][25]~q ;
wire \register[27][25]~q ;
wire \Mux38~7_combout ;
wire \Mux38~8_combout ;
wire \register[28][25]~q ;
wire \register[20][25]~q ;
wire \Mux38~4_combout ;
wire \Mux38~5_combout ;
wire \register[30][25]~feeder_combout ;
wire \register[30][25]~q ;
wire \register[26][25]~feeder_combout ;
wire \register[26][25]~q ;
wire \register[22][25]~q ;
wire \register[18][25]~q ;
wire \Mux38~2_combout ;
wire \Mux38~3_combout ;
wire \Mux38~6_combout ;
wire \register[12][25]~q ;
wire \Mux38~17_combout ;
wire \register[14][25]~q ;
wire \register[15][25]~q ;
wire \Mux38~18_combout ;
wire \register[5][25]~q ;
wire \Mux38~10_combout ;
wire \register[6][25]~q ;
wire \register[7][25]~q ;
wire \Mux38~11_combout ;
wire \register[2][25]~q ;
wire \register[3][25]~q ;
wire \register[1][25]~q ;
wire \Mux38~14_combout ;
wire \Mux38~15_combout ;
wire \register[9][25]~q ;
wire \register[11][25]~q ;
wire \register[8][25]~q ;
wire \register[10][25]~q ;
wire \Mux38~12_combout ;
wire \Mux38~13_combout ;
wire \Mux38~16_combout ;
wire \register~71_combout ;
wire \register[25][24]~feeder_combout ;
wire \register[25][24]~q ;
wire \register[29][24]~q ;
wire \register[17][24]~q ;
wire \Mux39~0_combout ;
wire \Mux39~1_combout ;
wire \register[16][24]~q ;
wire \register[24][24]~q ;
wire \Mux39~4_combout ;
wire \register[20][24]~q ;
wire \Mux39~5_combout ;
wire \register[22][24]~q ;
wire \register[30][24]~q ;
wire \register[26][24]~q ;
wire \Mux39~2_combout ;
wire \Mux39~3_combout ;
wire \Mux39~6_combout ;
wire \register[23][24]~q ;
wire \register[19][24]~q ;
wire \Mux39~7_combout ;
wire \register[27][24]~feeder_combout ;
wire \register[27][24]~q ;
wire \register[31][24]~feeder_combout ;
wire \register[31][24]~q ;
wire \Mux39~8_combout ;
wire \register[2][24]~feeder_combout ;
wire \register[2][24]~q ;
wire \register[1][24]~q ;
wire \register[3][24]~q ;
wire \Mux39~14_combout ;
wire \Mux39~15_combout ;
wire \register[7][24]~q ;
wire \register[6][24]~q ;
wire \Mux39~13_combout ;
wire \Mux39~16_combout ;
wire \register[15][24]~feeder_combout ;
wire \register[15][24]~q ;
wire \register[14][24]~feeder_combout ;
wire \register[14][24]~q ;
wire \register[12][24]~q ;
wire \register[13][24]~q ;
wire \Mux39~17_combout ;
wire \Mux39~18_combout ;
wire \register[11][24]~feeder_combout ;
wire \register[11][24]~q ;
wire \register[9][24]~feeder_combout ;
wire \register[9][24]~q ;
wire \register[8][24]~q ;
wire \register[10][24]~q ;
wire \Mux39~10_combout ;
wire \Mux39~11_combout ;
wire \register~72_combout ;
wire \register[31][23]~feeder_combout ;
wire \register[31][23]~q ;
wire \register[23][23]~q ;
wire \register[19][23]~q ;
wire \register[27][23]~feeder_combout ;
wire \register[27][23]~q ;
wire \Mux40~7_combout ;
wire \Mux40~8_combout ;
wire \register[29][23]~feeder_combout ;
wire \register[29][23]~q ;
wire \register[21][23]~q ;
wire \register[25][23]~q ;
wire \Mux40~0_combout ;
wire \Mux40~1_combout ;
wire \register[28][23]~feeder_combout ;
wire \register[28][23]~q ;
wire \register[24][23]~q ;
wire \register[20][23]~q ;
wire \Mux40~4_combout ;
wire \Mux40~5_combout ;
wire \register[22][23]~q ;
wire \Mux40~2_combout ;
wire \register[30][23]~q ;
wire \Mux40~3_combout ;
wire \Mux40~6_combout ;
wire \register[2][23]~q ;
wire \Mux40~15_combout ;
wire \register[9][23]~feeder_combout ;
wire \register[9][23]~q ;
wire \register[11][23]~q ;
wire \register[8][23]~q ;
wire \register[10][23]~q ;
wire \Mux40~12_combout ;
wire \Mux40~13_combout ;
wire \Mux40~16_combout ;
wire \register[15][23]~feeder_combout ;
wire \register[15][23]~q ;
wire \register[13][23]~q ;
wire \register[12][23]~q ;
wire \Mux40~17_combout ;
wire \register[14][23]~feeder_combout ;
wire \register[14][23]~q ;
wire \Mux40~18_combout ;
wire \register[5][23]~q ;
wire \register[4][23]~q ;
wire \Mux40~10_combout ;
wire \register[7][23]~q ;
wire \register[6][23]~q ;
wire \Mux40~11_combout ;
wire \register~73_combout ;
wire \register[29][22]~feeder_combout ;
wire \register[29][22]~q ;
wire \register[25][22]~feeder_combout ;
wire \register[25][22]~q ;
wire \register[17][22]~q ;
wire \register[21][22]~feeder_combout ;
wire \register[21][22]~q ;
wire \Mux41~0_combout ;
wire \Mux41~1_combout ;
wire \register[28][22]~feeder_combout ;
wire \register[28][22]~q ;
wire \register[16][22]~q ;
wire \register[24][22]~feeder_combout ;
wire \register[24][22]~q ;
wire \Mux41~4_combout ;
wire \register[20][22]~q ;
wire \Mux41~5_combout ;
wire \register[22][22]~q ;
wire \register[30][22]~q ;
wire \register[18][22]~q ;
wire \Mux41~2_combout ;
wire \Mux41~3_combout ;
wire \Mux41~6_combout ;
wire \register[27][22]~q ;
wire \register[31][22]~q ;
wire \register[19][22]~q ;
wire \Mux41~7_combout ;
wire \Mux41~8_combout ;
wire \register[15][22]~q ;
wire \register[13][22]~q ;
wire \register[12][22]~q ;
wire \Mux41~17_combout ;
wire \register[14][22]~q ;
wire \Mux41~18_combout ;
wire \register[2][22]~q ;
wire \register[1][22]~q ;
wire \register[3][22]~q ;
wire \Mux41~14_combout ;
wire \Mux41~15_combout ;
wire \register[7][22]~q ;
wire \register[5][22]~q ;
wire \register[4][22]~q ;
wire \Mux41~12_combout ;
wire \Mux41~13_combout ;
wire \Mux41~16_combout ;
wire \register[11][22]~q ;
wire \register[9][22]~q ;
wire \register[8][22]~q ;
wire \register[10][22]~q ;
wire \Mux41~10_combout ;
wire \Mux41~11_combout ;
wire \register~74_combout ;
wire \register[20][21]~q ;
wire \Mux42~4_combout ;
wire \register[24][21]~q ;
wire \Mux42~5_combout ;
wire \register[30][21]~feeder_combout ;
wire \register[30][21]~q ;
wire \register[26][21]~q ;
wire \register[18][21]~q ;
wire \register[22][21]~q ;
wire \Mux42~2_combout ;
wire \Mux42~3_combout ;
wire \Mux42~6_combout ;
wire \register[17][21]~q ;
wire \register[25][21]~feeder_combout ;
wire \register[25][21]~q ;
wire \Mux42~0_combout ;
wire \register[21][21]~q ;
wire \register[29][21]~q ;
wire \Mux42~1_combout ;
wire \register[23][21]~q ;
wire \register[31][21]~q ;
wire \register[19][21]~q ;
wire \register[27][21]~feeder_combout ;
wire \register[27][21]~q ;
wire \Mux42~7_combout ;
wire \Mux42~8_combout ;
wire \register[15][21]~feeder_combout ;
wire \register[15][21]~q ;
wire \register[14][21]~q ;
wire \register[13][21]~q ;
wire \register[12][21]~q ;
wire \Mux42~17_combout ;
wire \Mux42~18_combout ;
wire \register[7][21]~q ;
wire \register[6][21]~q ;
wire \register[4][21]~q ;
wire \Mux42~10_combout ;
wire \Mux42~11_combout ;
wire \register[11][21]~q ;
wire \register[9][21]~feeder_combout ;
wire \register[9][21]~q ;
wire \Mux42~13_combout ;
wire \register[2][21]~q ;
wire \register[3][21]~q ;
wire \register[1][21]~q ;
wire \Mux42~14_combout ;
wire \Mux42~15_combout ;
wire \Mux42~16_combout ;
wire \register~75_combout ;
wire \register[30][20]~feeder_combout ;
wire \register[30][20]~q ;
wire \register[22][20]~feeder_combout ;
wire \register[22][20]~q ;
wire \Mux43~3_combout ;
wire \register[28][20]~q ;
wire \register[20][20]~q ;
wire \Mux43~5_combout ;
wire \Mux43~6_combout ;
wire \register[31][20]~feeder_combout ;
wire \register[31][20]~q ;
wire \register[27][20]~q ;
wire \register[23][20]~feeder_combout ;
wire \register[23][20]~q ;
wire \register[19][20]~q ;
wire \Mux43~7_combout ;
wire \Mux43~8_combout ;
wire \register[29][20]~feeder_combout ;
wire \register[29][20]~q ;
wire \register[25][20]~q ;
wire \register[17][20]~q ;
wire \register[21][20]~feeder_combout ;
wire \register[21][20]~q ;
wire \Mux43~0_combout ;
wire \Mux43~1_combout ;
wire \register[6][20]~q ;
wire \register[7][20]~q ;
wire \register[5][20]~q ;
wire \Mux43~12_combout ;
wire \Mux43~13_combout ;
wire \register[3][20]~q ;
wire \register[1][20]~q ;
wire \Mux43~14_combout ;
wire \register[2][20]~q ;
wire \Mux43~15_combout ;
wire \Mux43~16_combout ;
wire \register[11][20]~q ;
wire \register[9][20]~q ;
wire \register[10][20]~q ;
wire \Mux43~10_combout ;
wire \Mux43~11_combout ;
wire \register[12][20]~q ;
wire \register[13][20]~q ;
wire \Mux43~17_combout ;
wire \register[14][20]~feeder_combout ;
wire \register[14][20]~q ;
wire \register[15][20]~q ;
wire \Mux43~18_combout ;
wire \register~76_combout ;
wire \register[31][19]~feeder_combout ;
wire \register[31][19]~q ;
wire \register[23][19]~q ;
wire \register[19][19]~q ;
wire \Mux44~7_combout ;
wire \Mux44~8_combout ;
wire \register[21][19]~q ;
wire \register[17][19]~q ;
wire \register[25][19]~feeder_combout ;
wire \register[25][19]~q ;
wire \Mux44~0_combout ;
wire \register[29][19]~feeder_combout ;
wire \register[29][19]~q ;
wire \Mux44~1_combout ;
wire \register[24][19]~q ;
wire \register[28][19]~q ;
wire \register[16][19]~feeder_combout ;
wire \register[16][19]~q ;
wire \register[20][19]~q ;
wire \Mux44~4_combout ;
wire \Mux44~5_combout ;
wire \register[30][19]~q ;
wire \register[26][19]~q ;
wire \register[22][19]~q ;
wire \Mux44~2_combout ;
wire \Mux44~3_combout ;
wire \Mux44~6_combout ;
wire \register[15][19]~q ;
wire \register[12][19]~q ;
wire \Mux44~17_combout ;
wire \register[14][19]~q ;
wire \Mux44~18_combout ;
wire \register[7][19]~q ;
wire \register[6][19]~q ;
wire \register[5][19]~q ;
wire \Mux44~10_combout ;
wire \Mux44~11_combout ;
wire \register[3][19]~q ;
wire \register[1][19]~q ;
wire \Mux44~14_combout ;
wire \Mux44~15_combout ;
wire \register[10][19]~q ;
wire \register[8][19]~q ;
wire \Mux44~12_combout ;
wire \register[11][19]~q ;
wire \register[9][19]~q ;
wire \Mux44~13_combout ;
wire \Mux44~16_combout ;
wire \register~77_combout ;
wire \register[22][18]~feeder_combout ;
wire \register[22][18]~q ;
wire \register[30][18]~q ;
wire \register[26][18]~q ;
wire \register[18][18]~q ;
wire \Mux45~2_combout ;
wire \Mux45~3_combout ;
wire \register[24][18]~feeder_combout ;
wire \register[24][18]~q ;
wire \register[16][18]~q ;
wire \Mux45~4_combout ;
wire \register[20][18]~q ;
wire \Mux45~5_combout ;
wire \Mux45~6_combout ;
wire \register[25][18]~feeder_combout ;
wire \register[25][18]~q ;
wire \register[29][18]~q ;
wire \register[17][18]~feeder_combout ;
wire \register[17][18]~q ;
wire \register[21][18]~feeder_combout ;
wire \register[21][18]~q ;
wire \Mux45~0_combout ;
wire \Mux45~1_combout ;
wire \register[27][18]~feeder_combout ;
wire \register[27][18]~q ;
wire \register[31][18]~q ;
wire \register[23][18]~q ;
wire \register[19][18]~q ;
wire \Mux45~7_combout ;
wire \Mux45~8_combout ;
wire \register[9][18]~feeder_combout ;
wire \register[9][18]~q ;
wire \register[10][18]~q ;
wire \Mux45~10_combout ;
wire \register[11][18]~q ;
wire \Mux45~11_combout ;
wire \register[12][18]~q ;
wire \Mux45~17_combout ;
wire \register[14][18]~q ;
wire \register[15][18]~q ;
wire \Mux45~18_combout ;
wire \register[7][18]~q ;
wire \register[6][18]~feeder_combout ;
wire \register[6][18]~q ;
wire \Mux45~13_combout ;
wire \register[2][18]~q ;
wire \register[3][18]~q ;
wire \Mux45~14_combout ;
wire \Mux45~15_combout ;
wire \Mux45~16_combout ;
wire \register~78_combout ;
wire \register[30][17]~q ;
wire \register[18][17]~q ;
wire \Mux46~2_combout ;
wire \Mux46~3_combout ;
wire \register[24][17]~q ;
wire \register[16][17]~feeder_combout ;
wire \register[16][17]~q ;
wire \register[20][17]~q ;
wire \Mux46~4_combout ;
wire \Mux46~5_combout ;
wire \Mux46~6_combout ;
wire \register[31][17]~feeder_combout ;
wire \register[31][17]~q ;
wire \register[23][17]~feeder_combout ;
wire \register[23][17]~q ;
wire \register[27][17]~q ;
wire \Mux46~7_combout ;
wire \Mux46~8_combout ;
wire \register[21][17]~q ;
wire \register[17][17]~q ;
wire \register[25][17]~feeder_combout ;
wire \register[25][17]~q ;
wire \Mux46~0_combout ;
wire \register[29][17]~feeder_combout ;
wire \register[29][17]~q ;
wire \Mux46~1_combout ;
wire \register[7][17]~q ;
wire \register[6][17]~q ;
wire \register[4][17]~q ;
wire \register[5][17]~q ;
wire \Mux46~10_combout ;
wire \Mux46~11_combout ;
wire \register[15][17]~q ;
wire \register[14][17]~q ;
wire \register[12][17]~q ;
wire \register[13][17]~q ;
wire \Mux46~17_combout ;
wire \Mux46~18_combout ;
wire \register[9][17]~q ;
wire \register[11][17]~q ;
wire \Mux46~13_combout ;
wire \register[1][17]~q ;
wire \register[3][17]~q ;
wire \Mux46~14_combout ;
wire \register[2][17]~feeder_combout ;
wire \register[2][17]~q ;
wire \Mux46~15_combout ;
wire \Mux46~16_combout ;
wire \register~79_combout ;
wire \register[27][16]~feeder_combout ;
wire \register[27][16]~q ;
wire \register[31][16]~feeder_combout ;
wire \register[31][16]~q ;
wire \register[23][16]~q ;
wire \Mux47~7_combout ;
wire \Mux47~8_combout ;
wire \register[22][16]~q ;
wire \register[30][16]~q ;
wire \Mux47~3_combout ;
wire \register[20][16]~q ;
wire \register[28][16]~q ;
wire \register[24][16]~q ;
wire \register[16][16]~feeder_combout ;
wire \register[16][16]~q ;
wire \Mux47~4_combout ;
wire \Mux47~5_combout ;
wire \Mux47~6_combout ;
wire \register[25][16]~q ;
wire \register[29][16]~feeder_combout ;
wire \register[29][16]~q ;
wire \register[17][16]~q ;
wire \Mux47~0_combout ;
wire \Mux47~1_combout ;
wire \register[10][16]~q ;
wire \register[8][16]~q ;
wire \Mux47~10_combout ;
wire \register[9][16]~q ;
wire \register[11][16]~q ;
wire \Mux47~11_combout ;
wire \register[15][16]~feeder_combout ;
wire \register[15][16]~q ;
wire \register[14][16]~q ;
wire \register[12][16]~q ;
wire \register[13][16]~q ;
wire \Mux47~17_combout ;
wire \Mux47~18_combout ;
wire \register[6][16]~q ;
wire \register[7][16]~q ;
wire \register[4][16]~q ;
wire \register[5][16]~q ;
wire \Mux47~12_combout ;
wire \Mux47~13_combout ;
wire \register[2][16]~q ;
wire \register[1][16]~q ;
wire \register[3][16]~q ;
wire \Mux47~14_combout ;
wire \Mux47~15_combout ;
wire \Mux47~16_combout ;
wire \register~80_combout ;
wire \register[28][15]~feeder_combout ;
wire \register[28][15]~q ;
wire \register[16][15]~q ;
wire \register[20][15]~feeder_combout ;
wire \register[20][15]~q ;
wire \Mux48~4_combout ;
wire \register[24][15]~feeder_combout ;
wire \register[24][15]~q ;
wire \Mux48~5_combout ;
wire \register[26][15]~q ;
wire \register[30][15]~feeder_combout ;
wire \register[30][15]~q ;
wire \register[18][15]~q ;
wire \register[22][15]~feeder_combout ;
wire \register[22][15]~q ;
wire \Mux48~2_combout ;
wire \Mux48~3_combout ;
wire \Mux48~6_combout ;
wire \register[23][15]~feeder_combout ;
wire \register[23][15]~q ;
wire \register[31][15]~feeder_combout ;
wire \register[31][15]~q ;
wire \register[27][15]~q ;
wire \register[19][15]~q ;
wire \Mux48~7_combout ;
wire \Mux48~8_combout ;
wire \register[29][15]~feeder_combout ;
wire \register[29][15]~q ;
wire \register[21][15]~q ;
wire \register[25][15]~feeder_combout ;
wire \register[25][15]~q ;
wire \register[17][15]~q ;
wire \Mux48~0_combout ;
wire \Mux48~1_combout ;
wire \register[7][15]~q ;
wire \register[6][15]~q ;
wire \register[5][15]~q ;
wire \register[4][15]~q ;
wire \Mux48~10_combout ;
wire \Mux48~11_combout ;
wire \register[14][15]~q ;
wire \register[12][15]~q ;
wire \register[13][15]~q ;
wire \Mux48~17_combout ;
wire \register[15][15]~q ;
wire \Mux48~18_combout ;
wire \register[3][15]~q ;
wire \register[1][15]~q ;
wire \Mux48~14_combout ;
wire \Mux48~15_combout ;
wire \register[11][15]~q ;
wire \register[9][15]~q ;
wire \Mux48~13_combout ;
wire \Mux48~16_combout ;
wire \register~81_combout ;
wire \register[27][14]~q ;
wire \register[31][14]~feeder_combout ;
wire \register[31][14]~q ;
wire \register[23][14]~q ;
wire \Mux49~7_combout ;
wire \Mux49~8_combout ;
wire \register[25][14]~q ;
wire \register[29][14]~q ;
wire \register[17][14]~q ;
wire \register[21][14]~feeder_combout ;
wire \register[21][14]~q ;
wire \Mux49~0_combout ;
wire \Mux49~1_combout ;
wire \register[30][14]~q ;
wire \register[26][14]~q ;
wire \register[18][14]~q ;
wire \Mux49~2_combout ;
wire \Mux49~3_combout ;
wire \register[20][14]~q ;
wire \register[28][14]~feeder_combout ;
wire \register[28][14]~q ;
wire \register[24][14]~q ;
wire \register[16][14]~feeder_combout ;
wire \register[16][14]~q ;
wire \Mux49~4_combout ;
wire \Mux49~5_combout ;
wire \Mux49~6_combout ;
wire \register[2][14]~q ;
wire \register[1][14]~q ;
wire \register[3][14]~q ;
wire \Mux49~14_combout ;
wire \Mux49~15_combout ;
wire \register[5][14]~q ;
wire \register[4][14]~q ;
wire \Mux49~12_combout ;
wire \register[7][14]~q ;
wire \register[6][14]~q ;
wire \Mux49~13_combout ;
wire \Mux49~16_combout ;
wire \register[9][14]~feeder_combout ;
wire \register[9][14]~q ;
wire \register[11][14]~q ;
wire \register[10][14]~q ;
wire \register[8][14]~q ;
wire \Mux49~10_combout ;
wire \Mux49~11_combout ;
wire \register[14][14]~q ;
wire \register[15][14]~q ;
wire \register[13][14]~q ;
wire \register[12][14]~q ;
wire \Mux49~17_combout ;
wire \Mux49~18_combout ;
wire \register~82_combout ;
wire \register[29][13]~feeder_combout ;
wire \register[29][13]~q ;
wire \register[21][13]~feeder_combout ;
wire \register[21][13]~q ;
wire \register[17][13]~q ;
wire \Mux50~0_combout ;
wire \Mux50~1_combout ;
wire \register[23][13]~feeder_combout ;
wire \register[23][13]~q ;
wire \register[31][13]~q ;
wire \register[27][13]~q ;
wire \register[19][13]~q ;
wire \Mux50~7_combout ;
wire \Mux50~8_combout ;
wire \register[24][13]~feeder_combout ;
wire \register[24][13]~q ;
wire \register[20][13]~q ;
wire \register[16][13]~q ;
wire \Mux50~4_combout ;
wire \Mux50~5_combout ;
wire \register[26][13]~q ;
wire \register[30][13]~q ;
wire \register[18][13]~q ;
wire \Mux50~2_combout ;
wire \Mux50~3_combout ;
wire \Mux50~6_combout ;
wire \register[12][13]~q ;
wire \Mux50~17_combout ;
wire \register[15][13]~q ;
wire \register[14][13]~q ;
wire \Mux50~18_combout ;
wire \register[7][13]~q ;
wire \register[5][13]~q ;
wire \Mux50~10_combout ;
wire \register[6][13]~q ;
wire \Mux50~11_combout ;
wire \register[2][13]~q ;
wire \register[1][13]~q ;
wire \Mux50~14_combout ;
wire \Mux50~15_combout ;
wire \register[9][13]~q ;
wire \register[10][13]~q ;
wire \Mux50~12_combout ;
wire \Mux50~13_combout ;
wire \Mux50~16_combout ;
wire \register~83_combout ;
wire \register[31][12]~feeder_combout ;
wire \register[31][12]~q ;
wire \register[19][12]~q ;
wire \register[23][12]~q ;
wire \Mux51~7_combout ;
wire \register[27][12]~feeder_combout ;
wire \register[27][12]~q ;
wire \Mux51~8_combout ;
wire \register[17][12]~q ;
wire \register[21][12]~feeder_combout ;
wire \register[21][12]~q ;
wire \Mux51~0_combout ;
wire \register[25][12]~q ;
wire \register[29][12]~feeder_combout ;
wire \register[29][12]~q ;
wire \Mux51~1_combout ;
wire \register[30][12]~feeder_combout ;
wire \register[30][12]~q ;
wire \register[26][12]~q ;
wire \register[18][12]~feeder_combout ;
wire \register[18][12]~q ;
wire \Mux51~2_combout ;
wire \Mux51~3_combout ;
wire \register[28][12]~feeder_combout ;
wire \register[28][12]~q ;
wire \register[20][12]~q ;
wire \register[16][12]~q ;
wire \register[24][12]~feeder_combout ;
wire \register[24][12]~q ;
wire \Mux51~4_combout ;
wire \Mux51~5_combout ;
wire \Mux51~6_combout ;
wire \register[9][12]~q ;
wire \register[11][12]~q ;
wire \register[10][12]~q ;
wire \register[8][12]~q ;
wire \Mux51~10_combout ;
wire \Mux51~11_combout ;
wire \register[14][12]~q ;
wire \register[15][12]~q ;
wire \register[12][12]~q ;
wire \register[13][12]~q ;
wire \Mux51~17_combout ;
wire \Mux51~18_combout ;
wire \register[6][12]~feeder_combout ;
wire \register[6][12]~q ;
wire \register[7][12]~q ;
wire \register[5][12]~q ;
wire \Mux51~12_combout ;
wire \Mux51~13_combout ;
wire \register[2][12]~q ;
wire \register[3][12]~q ;
wire \register[1][12]~q ;
wire \Mux51~14_combout ;
wire \Mux51~15_combout ;
wire \Mux51~16_combout ;
wire \register~84_combout ;
wire \register[21][11]~feeder_combout ;
wire \register[21][11]~q ;
wire \register[17][11]~q ;
wire \register[25][11]~feeder_combout ;
wire \register[25][11]~q ;
wire \Mux52~0_combout ;
wire \register[29][11]~q ;
wire \Mux52~1_combout ;
wire \register[23][11]~q ;
wire \register[31][11]~q ;
wire \register[19][11]~q ;
wire \register[27][11]~q ;
wire \Mux52~7_combout ;
wire \Mux52~8_combout ;
wire \register[26][11]~q ;
wire \register[30][11]~q ;
wire \register[18][11]~q ;
wire \Mux52~2_combout ;
wire \Mux52~3_combout ;
wire \register[28][11]~feeder_combout ;
wire \register[28][11]~q ;
wire \register[16][11]~feeder_combout ;
wire \register[16][11]~q ;
wire \register[20][11]~q ;
wire \Mux52~4_combout ;
wire \Mux52~5_combout ;
wire \Mux52~6_combout ;
wire \register[7][11]~q ;
wire \register[4][11]~q ;
wire \register[5][11]~q ;
wire \Mux52~10_combout ;
wire \register[6][11]~q ;
wire \Mux52~11_combout ;
wire \register[14][11]~feeder_combout ;
wire \register[14][11]~q ;
wire \register[13][11]~q ;
wire \register[12][11]~q ;
wire \Mux52~17_combout ;
wire \register[15][11]~q ;
wire \Mux52~18_combout ;
wire \register[2][11]~q ;
wire \register[1][11]~q ;
wire \register[3][11]~q ;
wire \Mux52~14_combout ;
wire \Mux52~15_combout ;
wire \register[9][11]~q ;
wire \register[10][11]~q ;
wire \register[8][11]~q ;
wire \Mux52~12_combout ;
wire \Mux52~13_combout ;
wire \Mux52~16_combout ;
wire \register~85_combout ;
wire \register[28][10]~feeder_combout ;
wire \register[28][10]~q ;
wire \register[24][10]~q ;
wire \register[16][10]~feeder_combout ;
wire \register[16][10]~q ;
wire \Mux53~4_combout ;
wire \Mux53~5_combout ;
wire \register[26][10]~feeder_combout ;
wire \register[26][10]~q ;
wire \register[18][10]~q ;
wire \Mux53~2_combout ;
wire \register[30][10]~q ;
wire \Mux53~3_combout ;
wire \Mux53~6_combout ;
wire \register[31][10]~feeder_combout ;
wire \register[31][10]~q ;
wire \register[23][10]~q ;
wire \register[19][10]~q ;
wire \Mux53~7_combout ;
wire \register[27][10]~q ;
wire \Mux53~8_combout ;
wire \register[29][10]~q ;
wire \register[25][10]~q ;
wire \register[21][10]~q ;
wire \Mux53~0_combout ;
wire \Mux53~1_combout ;
wire \register[11][10]~q ;
wire \register[9][10]~q ;
wire \register[8][10]~q ;
wire \Mux53~10_combout ;
wire \Mux53~11_combout ;
wire \register[15][10]~q ;
wire \register[14][10]~q ;
wire \register[12][10]~q ;
wire \register[13][10]~q ;
wire \Mux53~17_combout ;
wire \Mux53~18_combout ;
wire \register[1][10]~q ;
wire \register[3][10]~q ;
wire \Mux53~14_combout ;
wire \register[2][10]~q ;
wire \Mux53~15_combout ;
wire \register[4][10]~q ;
wire \register[5][10]~q ;
wire \Mux53~12_combout ;
wire \register[7][10]~feeder_combout ;
wire \register[7][10]~q ;
wire \Mux53~13_combout ;
wire \Mux53~16_combout ;
wire \register~86_combout ;
wire \register[28][9]~feeder_combout ;
wire \register[28][9]~q ;
wire \register[20][9]~q ;
wire \register[16][9]~q ;
wire \Mux54~4_combout ;
wire \Mux54~5_combout ;
wire \register[18][9]~q ;
wire \Mux54~2_combout ;
wire \register[26][9]~q ;
wire \Mux54~3_combout ;
wire \Mux54~6_combout ;
wire \register[23][9]~q ;
wire \register[31][9]~feeder_combout ;
wire \register[31][9]~q ;
wire \register[19][9]~q ;
wire \register[27][9]~feeder_combout ;
wire \register[27][9]~q ;
wire \Mux54~7_combout ;
wire \Mux54~8_combout ;
wire \register[29][9]~q ;
wire \register[25][9]~q ;
wire \Mux54~0_combout ;
wire \register[21][9]~feeder_combout ;
wire \register[21][9]~q ;
wire \Mux54~1_combout ;
wire \register[15][9]~q ;
wire \register[14][9]~feeder_combout ;
wire \register[14][9]~q ;
wire \register[12][9]~q ;
wire \register[13][9]~q ;
wire \Mux54~17_combout ;
wire \Mux54~18_combout ;
wire \register[6][9]~feeder_combout ;
wire \register[6][9]~q ;
wire \register[4][9]~q ;
wire \register[5][9]~q ;
wire \Mux54~10_combout ;
wire \register[7][9]~q ;
wire \Mux54~11_combout ;
wire \register[11][9]~feeder_combout ;
wire \register[11][9]~q ;
wire \register[9][9]~feeder_combout ;
wire \register[9][9]~q ;
wire \register[8][9]~q ;
wire \register[10][9]~q ;
wire \Mux54~12_combout ;
wire \Mux54~13_combout ;
wire \register[1][9]~q ;
wire \register[3][9]~q ;
wire \Mux54~14_combout ;
wire \register[2][9]~q ;
wire \Mux54~15_combout ;
wire \Mux54~16_combout ;
wire \register~87_combout ;
wire \register[29][8]~feeder_combout ;
wire \register[29][8]~q ;
wire \register[25][8]~q ;
wire \register[21][8]~q ;
wire \register[17][8]~q ;
wire \Mux55~0_combout ;
wire \Mux55~1_combout ;
wire \register[22][8]~feeder_combout ;
wire \register[22][8]~q ;
wire \register[30][8]~q ;
wire \Mux55~3_combout ;
wire \register[28][8]~q ;
wire \register[24][8]~feeder_combout ;
wire \register[24][8]~q ;
wire \register[16][8]~feeder_combout ;
wire \register[16][8]~q ;
wire \Mux55~4_combout ;
wire \Mux55~5_combout ;
wire \Mux55~6_combout ;
wire \register[27][8]~q ;
wire \register[31][8]~q ;
wire \register[19][8]~q ;
wire \register[23][8]~q ;
wire \Mux55~7_combout ;
wire \Mux55~8_combout ;
wire \register[13][8]~q ;
wire \Mux55~17_combout ;
wire \register[14][8]~feeder_combout ;
wire \register[14][8]~q ;
wire \register[15][8]~q ;
wire \Mux55~18_combout ;
wire \register[10][8]~q ;
wire \Mux55~10_combout ;
wire \register[11][8]~q ;
wire \register[9][8]~q ;
wire \Mux55~11_combout ;
wire \register[6][8]~q ;
wire \register[5][8]~q ;
wire \Mux55~12_combout ;
wire \Mux55~13_combout ;
wire \register[2][8]~q ;
wire \register[3][8]~q ;
wire \register[1][8]~q ;
wire \Mux55~14_combout ;
wire \Mux55~15_combout ;
wire \Mux55~16_combout ;
wire \register~88_combout ;
wire \register[23][7]~q ;
wire \register[31][7]~q ;
wire \register[19][7]~q ;
wire \register[27][7]~feeder_combout ;
wire \register[27][7]~q ;
wire \Mux56~7_combout ;
wire \Mux56~8_combout ;
wire \register[29][7]~feeder_combout ;
wire \register[29][7]~q ;
wire \register[21][7]~q ;
wire \register[25][7]~feeder_combout ;
wire \register[25][7]~q ;
wire \register[17][7]~q ;
wire \Mux56~0_combout ;
wire \Mux56~1_combout ;
wire \register[24][7]~feeder_combout ;
wire \register[24][7]~q ;
wire \register[28][7]~q ;
wire \register[16][7]~q ;
wire \Mux56~4_combout ;
wire \Mux56~5_combout ;
wire \register[26][7]~q ;
wire \register[30][7]~q ;
wire \register[18][7]~q ;
wire \register[22][7]~q ;
wire \Mux56~2_combout ;
wire \Mux56~3_combout ;
wire \Mux56~6_combout ;
wire \register[11][7]~q ;
wire \register[9][7]~q ;
wire \Mux56~13_combout ;
wire \register[2][7]~q ;
wire \register[3][7]~feeder_combout ;
wire \register[3][7]~q ;
wire \register[1][7]~feeder_combout ;
wire \register[1][7]~q ;
wire \Mux56~14_combout ;
wire \Mux56~15_combout ;
wire \Mux56~16_combout ;
wire \register[7][7]~q ;
wire \register[6][7]~q ;
wire \register[4][7]~q ;
wire \register[5][7]~q ;
wire \Mux56~10_combout ;
wire \Mux56~11_combout ;
wire \register[15][7]~feeder_combout ;
wire \register[15][7]~q ;
wire \register[14][7]~q ;
wire \register[13][7]~q ;
wire \register[12][7]~q ;
wire \Mux56~17_combout ;
wire \Mux56~18_combout ;
wire \register~89_combout ;
wire \register[23][6]~q ;
wire \register[19][6]~q ;
wire \Mux57~7_combout ;
wire \register[31][6]~feeder_combout ;
wire \register[31][6]~q ;
wire \register[27][6]~q ;
wire \Mux57~8_combout ;
wire \register[22][6]~q ;
wire \register[30][6]~q ;
wire \Mux57~3_combout ;
wire \register[20][6]~q ;
wire \register[28][6]~q ;
wire \register[24][6]~q ;
wire \Mux57~4_combout ;
wire \Mux57~5_combout ;
wire \Mux57~6_combout ;
wire \register[29][6]~feeder_combout ;
wire \register[29][6]~q ;
wire \register[21][6]~q ;
wire \Mux57~0_combout ;
wire \register[25][6]~feeder_combout ;
wire \register[25][6]~q ;
wire \Mux57~1_combout ;
wire \register[11][6]~q ;
wire \register[9][6]~feeder_combout ;
wire \register[9][6]~q ;
wire \register[8][6]~q ;
wire \register[10][6]~q ;
wire \Mux57~10_combout ;
wire \Mux57~11_combout ;
wire \register[2][6]~q ;
wire \register[1][6]~feeder_combout ;
wire \register[1][6]~q ;
wire \register[3][6]~feeder_combout ;
wire \register[3][6]~q ;
wire \Mux57~14_combout ;
wire \Mux57~15_combout ;
wire \register[7][6]~q ;
wire \register[4][6]~q ;
wire \Mux57~12_combout ;
wire \Mux57~13_combout ;
wire \Mux57~16_combout ;
wire \register[15][6]~q ;
wire \register[12][6]~q ;
wire \register[13][6]~q ;
wire \Mux57~17_combout ;
wire \register[14][6]~feeder_combout ;
wire \register[14][6]~q ;
wire \Mux57~18_combout ;
wire \register~90_combout ;
wire \register[23][5]~q ;
wire \register[31][5]~q ;
wire \register[19][5]~q ;
wire \register[27][5]~feeder_combout ;
wire \register[27][5]~q ;
wire \Mux58~7_combout ;
wire \Mux58~8_combout ;
wire \register[29][5]~feeder_combout ;
wire \register[29][5]~q ;
wire \register[21][5]~q ;
wire \register[17][5]~q ;
wire \register[25][5]~q ;
wire \Mux58~0_combout ;
wire \Mux58~1_combout ;
wire \register[26][5]~q ;
wire \register[30][5]~q ;
wire \register[18][5]~q ;
wire \register[22][5]~q ;
wire \Mux58~2_combout ;
wire \Mux58~3_combout ;
wire \register[20][5]~feeder_combout ;
wire \register[20][5]~q ;
wire \Mux58~4_combout ;
wire \register[24][5]~feeder_combout ;
wire \register[24][5]~q ;
wire \Mux58~5_combout ;
wire \Mux58~6_combout ;
wire \register[7][5]~q ;
wire \register[5][5]~q ;
wire \register[4][5]~q ;
wire \Mux58~10_combout ;
wire \register[6][5]~q ;
wire \Mux58~11_combout ;
wire \register[15][5]~q ;
wire \register[14][5]~feeder_combout ;
wire \register[14][5]~q ;
wire \register[12][5]~q ;
wire \register[13][5]~q ;
wire \Mux58~17_combout ;
wire \Mux58~18_combout ;
wire \register[2][5]~q ;
wire \register[1][5]~q ;
wire \register[3][5]~q ;
wire \Mux58~14_combout ;
wire \Mux58~15_combout ;
wire \register[9][5]~q ;
wire \register[11][5]~q ;
wire \Mux58~13_combout ;
wire \Mux58~16_combout ;
wire \register~91_combout ;
wire \register[23][2]~q ;
wire \register[31][2]~q ;
wire \register[19][2]~q ;
wire \register[27][2]~feeder_combout ;
wire \register[27][2]~q ;
wire \Mux29~7_combout ;
wire \Mux29~8_combout ;
wire \register[29][2]~q ;
wire \register[21][2]~q ;
wire \register[25][2]~q ;
wire \Mux29~0_combout ;
wire \Mux29~1_combout ;
wire \register[24][2]~feeder_combout ;
wire \register[24][2]~q ;
wire \register[28][2]~q ;
wire \register[20][2]~q ;
wire \register[16][2]~q ;
wire \Mux29~4_combout ;
wire \Mux29~5_combout ;
wire \register[30][2]~q ;
wire \register[22][2]~q ;
wire \register[18][2]~q ;
wire \Mux29~2_combout ;
wire \Mux29~3_combout ;
wire \Mux29~6_combout ;
wire \register[7][2]~q ;
wire \register[6][2]~q ;
wire \register[4][2]~q ;
wire \register[5][2]~q ;
wire \Mux29~10_combout ;
wire \Mux29~11_combout ;
wire \register[15][2]~q ;
wire \register[12][2]~q ;
wire \register[13][2]~q ;
wire \Mux29~17_combout ;
wire \register[14][2]~feeder_combout ;
wire \register[14][2]~q ;
wire \Mux29~18_combout ;
wire \register[2][2]~q ;
wire \Mux29~15_combout ;
wire \register[9][2]~q ;
wire \register[11][2]~q ;
wire \register[8][2]~q ;
wire \register[10][2]~q ;
wire \Mux29~12_combout ;
wire \Mux29~13_combout ;
wire \Mux29~16_combout ;
wire \register~92_combout ;
wire \register[29][1]~q ;
wire \register[21][1]~q ;
wire \register[17][1]~q ;
wire \Mux30~0_combout ;
wire \register[25][1]~feeder_combout ;
wire \register[25][1]~q ;
wire \Mux30~1_combout ;
wire \register[30][1]~feeder_combout ;
wire \register[30][1]~q ;
wire \register[22][1]~q ;
wire \register[18][1]~q ;
wire \Mux30~2_combout ;
wire \Mux30~3_combout ;
wire \register[28][1]~feeder_combout ;
wire \register[28][1]~q ;
wire \register[16][1]~feeder_combout ;
wire \register[16][1]~q ;
wire \Mux30~4_combout ;
wire \Mux30~5_combout ;
wire \Mux30~6_combout ;
wire \register[27][1]~feeder_combout ;
wire \register[27][1]~q ;
wire \register[31][1]~q ;
wire \register[19][1]~q ;
wire \register[23][1]~q ;
wire \Mux30~7_combout ;
wire \Mux30~8_combout ;
wire \register[3][1]~q ;
wire \register[1][1]~q ;
wire \Mux30~14_combout ;
wire \Mux30~15_combout ;
wire \register[6][1]~q ;
wire \register[7][1]~q ;
wire \register[5][1]~q ;
wire \register[4][1]~q ;
wire \Mux30~12_combout ;
wire \Mux30~13_combout ;
wire \Mux30~16_combout ;
wire \register[11][1]~q ;
wire \register[10][1]~q ;
wire \Mux30~10_combout ;
wire \register[9][1]~q ;
wire \Mux30~11_combout ;
wire \register[13][1]~q ;
wire \Mux30~17_combout ;
wire \register[14][1]~feeder_combout ;
wire \register[14][1]~q ;
wire \register[15][1]~q ;
wire \Mux30~18_combout ;
wire \register~93_combout ;
wire \register[29][0]~feeder_combout ;
wire \register[29][0]~q ;
wire \register[25][0]~feeder_combout ;
wire \register[25][0]~q ;
wire \register[17][0]~q ;
wire \register[21][0]~q ;
wire \Mux63~0_combout ;
wire \Mux63~1_combout ;
wire \register[27][0]~feeder_combout ;
wire \register[27][0]~q ;
wire \register[31][0]~feeder_combout ;
wire \register[31][0]~q ;
wire \register[19][0]~q ;
wire \register[23][0]~q ;
wire \Mux63~7_combout ;
wire \Mux63~8_combout ;
wire \register[30][0]~q ;
wire \register[18][0]~q ;
wire \register[26][0]~q ;
wire \Mux63~2_combout ;
wire \Mux63~3_combout ;
wire \register[28][0]~q ;
wire \register[24][0]~q ;
wire \register[16][0]~feeder_combout ;
wire \register[16][0]~q ;
wire \Mux63~4_combout ;
wire \Mux63~5_combout ;
wire \Mux63~6_combout ;
wire \register[11][0]~q ;
wire \register[9][0]~q ;
wire \register[10][0]~feeder_combout ;
wire \register[10][0]~q ;
wire \Mux63~10_combout ;
wire \Mux63~11_combout ;
wire \register[6][0]~q ;
wire \register[7][0]~q ;
wire \register[4][0]~q ;
wire \register[5][0]~q ;
wire \Mux63~12_combout ;
wire \Mux63~13_combout ;
wire \register[2][0]~feeder_combout ;
wire \register[2][0]~q ;
wire \register[3][0]~q ;
wire \Mux63~14_combout ;
wire \Mux63~15_combout ;
wire \Mux63~16_combout ;
wire \register[15][0]~q ;
wire \register[14][0]~q ;
wire \register[12][0]~q ;
wire \register[13][0]~q ;
wire \Mux63~17_combout ;
wire \Mux63~18_combout ;
wire \Mux62~2_combout ;
wire \register[26][1]~feeder_combout ;
wire \register[26][1]~q ;
wire \Mux62~3_combout ;
wire \register[20][1]~q ;
wire \Mux62~4_combout ;
wire \Mux62~5_combout ;
wire \Mux62~6_combout ;
wire \Mux62~0_combout ;
wire \Mux62~1_combout ;
wire \Mux62~7_combout ;
wire \Mux62~8_combout ;
wire \Mux62~10_combout ;
wire \Mux62~11_combout ;
wire \register[12][1]~q ;
wire \Mux62~17_combout ;
wire \Mux62~18_combout ;
wire \register[8][1]~q ;
wire \Mux62~12_combout ;
wire \Mux62~13_combout ;
wire \register[2][1]~q ;
wire \Mux62~14_combout ;
wire \Mux62~15_combout ;
wire \Mux62~16_combout ;
wire \register~94_combout ;
wire \register[21][4]~feeder_combout ;
wire \register[21][4]~q ;
wire \register[25][4]~q ;
wire \Mux27~0_combout ;
wire \register[29][4]~feeder_combout ;
wire \register[29][4]~q ;
wire \Mux27~1_combout ;
wire \register[23][4]~feeder_combout ;
wire \register[23][4]~q ;
wire \register[31][4]~q ;
wire \register[19][4]~q ;
wire \register[27][4]~q ;
wire \Mux27~7_combout ;
wire \Mux27~8_combout ;
wire \register[26][4]~q ;
wire \register[30][4]~q ;
wire \register[18][4]~q ;
wire \Mux27~2_combout ;
wire \Mux27~3_combout ;
wire \register[24][4]~q ;
wire \register[20][4]~q ;
wire \register[16][4]~q ;
wire \Mux27~4_combout ;
wire \Mux27~5_combout ;
wire \Mux27~6_combout ;
wire \register[7][4]~q ;
wire \register[6][4]~q ;
wire \register[5][4]~q ;
wire \register[4][4]~q ;
wire \Mux27~10_combout ;
wire \Mux27~11_combout ;
wire \register[14][4]~q ;
wire \register[15][4]~feeder_combout ;
wire \register[15][4]~q ;
wire \register[12][4]~q ;
wire \register[13][4]~q ;
wire \Mux27~17_combout ;
wire \Mux27~18_combout ;
wire \register[1][4]~q ;
wire \Mux27~14_combout ;
wire \Mux27~15_combout ;
wire \register[9][4]~q ;
wire \register[11][4]~q ;
wire \register[8][4]~q ;
wire \register[10][4]~q ;
wire \Mux27~12_combout ;
wire \Mux27~13_combout ;
wire \Mux27~16_combout ;
wire \register~95_combout ;
wire \register[20][3]~q ;
wire \register[16][3]~q ;
wire \register[24][3]~feeder_combout ;
wire \register[24][3]~q ;
wire \Mux28~4_combout ;
wire \Mux28~5_combout ;
wire \register[22][3]~q ;
wire \register[30][3]~q ;
wire \register[26][3]~feeder_combout ;
wire \register[26][3]~q ;
wire \register[18][3]~feeder_combout ;
wire \register[18][3]~q ;
wire \Mux28~2_combout ;
wire \Mux28~3_combout ;
wire \Mux28~6_combout ;
wire \register[31][3]~feeder_combout ;
wire \register[31][3]~q ;
wire \register[27][3]~feeder_combout ;
wire \register[27][3]~q ;
wire \register[23][3]~q ;
wire \register[19][3]~q ;
wire \Mux28~7_combout ;
wire \Mux28~8_combout ;
wire \register[29][3]~feeder_combout ;
wire \register[29][3]~q ;
wire \register[25][3]~feeder_combout ;
wire \register[25][3]~q ;
wire \register[21][3]~q ;
wire \register[17][3]~feeder_combout ;
wire \register[17][3]~q ;
wire \Mux28~0_combout ;
wire \Mux28~1_combout ;
wire \register[15][3]~q ;
wire \register[14][3]~q ;
wire \register[13][3]~q ;
wire \Mux28~17_combout ;
wire \Mux28~18_combout ;
wire \register[2][3]~q ;
wire \register[1][3]~q ;
wire \register[3][3]~q ;
wire \Mux28~14_combout ;
wire \Mux28~15_combout ;
wire \register[6][3]~q ;
wire \register[7][3]~q ;
wire \register[5][3]~q ;
wire \Mux28~12_combout ;
wire \Mux28~13_combout ;
wire \Mux28~16_combout ;
wire \register[9][3]~feeder_combout ;
wire \register[9][3]~q ;
wire \register[11][3]~q ;
wire \register[8][3]~q ;
wire \register[10][3]~q ;
wire \Mux28~10_combout ;
wire \Mux28~11_combout ;
wire \Mux61~7_combout ;
wire \Mux61~8_combout ;
wire \register[17][2]~q ;
wire \Mux61~0_combout ;
wire \Mux61~1_combout ;
wire \Mux61~4_combout ;
wire \Mux61~5_combout ;
wire \register[26][2]~q ;
wire \Mux61~2_combout ;
wire \Mux61~3_combout ;
wire \Mux61~6_combout ;
wire \Mux61~17_combout ;
wire \Mux61~18_combout ;
wire \Mux61~10_combout ;
wire \Mux61~11_combout ;
wire \Mux61~12_combout ;
wire \Mux61~13_combout ;
wire \Mux61~15_combout ;
wire \Mux61~16_combout ;
wire \Mux23~7_combout ;
wire \Mux23~8_combout ;
wire \Mux23~4_combout ;
wire \Mux23~5_combout ;
wire \register[18][8]~feeder_combout ;
wire \register[18][8]~q ;
wire \Mux23~2_combout ;
wire \Mux23~3_combout ;
wire \Mux23~6_combout ;
wire \Mux23~0_combout ;
wire \Mux23~1_combout ;
wire \register[12][8]~q ;
wire \Mux23~17_combout ;
wire \Mux23~18_combout ;
wire \register[7][8]~feeder_combout ;
wire \register[7][8]~q ;
wire \register[4][8]~q ;
wire \Mux23~10_combout ;
wire \Mux23~11_combout ;
wire \Mux23~14_combout ;
wire \Mux23~15_combout ;
wire \register[8][8]~q ;
wire \Mux23~12_combout ;
wire \Mux23~13_combout ;
wire \Mux23~16_combout ;
wire \Mux24~7_combout ;
wire \Mux24~8_combout ;
wire \Mux24~0_combout ;
wire \Mux24~1_combout ;
wire \Mux24~2_combout ;
wire \Mux24~3_combout ;
wire \register[20][7]~q ;
wire \Mux24~5_combout ;
wire \Mux24~6_combout ;
wire \Mux24~17_combout ;
wire \Mux24~18_combout ;
wire \register[10][7]~q ;
wire \register[8][7]~q ;
wire \Mux24~10_combout ;
wire \Mux24~11_combout ;
wire \Mux24~12_combout ;
wire \Mux24~13_combout ;
wire \Mux24~14_combout ;
wire \Mux24~15_combout ;
wire \Mux24~16_combout ;
wire \Mux25~7_combout ;
wire \Mux25~8_combout ;
wire \register[26][6]~q ;
wire \Mux25~3_combout ;
wire \register[16][6]~feeder_combout ;
wire \register[16][6]~q ;
wire \Mux25~4_combout ;
wire \Mux25~5_combout ;
wire \Mux25~6_combout ;
wire \register[17][6]~q ;
wire \Mux25~0_combout ;
wire \Mux25~1_combout ;
wire \Mux25~17_combout ;
wire \Mux25~18_combout ;
wire \register[5][6]~q ;
wire \Mux25~10_combout ;
wire \register[6][6]~q ;
wire \Mux25~11_combout ;
wire \Mux25~14_combout ;
wire \Mux25~15_combout ;
wire \Mux25~12_combout ;
wire \Mux25~13_combout ;
wire \Mux25~16_combout ;
wire \Mux26~7_combout ;
wire \Mux26~8_combout ;
wire \Mux26~2_combout ;
wire \Mux26~3_combout ;
wire \Mux26~4_combout ;
wire \Mux26~5_combout ;
wire \Mux26~6_combout ;
wire \Mux26~0_combout ;
wire \Mux26~1_combout ;
wire \Mux26~12_combout ;
wire \Mux26~13_combout ;
wire \Mux26~14_combout ;
wire \Mux26~15_combout ;
wire \Mux26~16_combout ;
wire \Mux26~17_combout ;
wire \Mux26~18_combout ;
wire \register[10][5]~q ;
wire \register[8][5]~q ;
wire \Mux26~10_combout ;
wire \Mux26~11_combout ;
wire \Mux60~7_combout ;
wire \Mux60~8_combout ;
wire \Mux60~0_combout ;
wire \Mux60~1_combout ;
wire \Mux60~4_combout ;
wire \register[28][3]~feeder_combout ;
wire \register[28][3]~q ;
wire \Mux60~5_combout ;
wire \Mux60~2_combout ;
wire \Mux60~3_combout ;
wire \Mux60~6_combout ;
wire \register[4][3]~q ;
wire \Mux60~10_combout ;
wire \Mux60~11_combout ;
wire \register[12][3]~q ;
wire \Mux60~17_combout ;
wire \Mux60~18_combout ;
wire \Mux60~15_combout ;
wire \Mux60~12_combout ;
wire \Mux60~13_combout ;
wire \Mux60~16_combout ;
wire \register[26][16]~q ;
wire \Mux15~2_combout ;
wire \Mux15~3_combout ;
wire \Mux15~5_combout ;
wire \Mux15~6_combout ;
wire \register[19][16]~q ;
wire \Mux15~7_combout ;
wire \Mux15~8_combout ;
wire \register[21][16]~q ;
wire \Mux15~0_combout ;
wire \Mux15~1_combout ;
wire \Mux15~10_combout ;
wire \Mux15~11_combout ;
wire \Mux15~17_combout ;
wire \Mux15~18_combout ;
wire \Mux15~14_combout ;
wire \Mux15~15_combout ;
wire \Mux15~12_combout ;
wire \Mux15~13_combout ;
wire \Mux15~16_combout ;
wire \Mux16~0_combout ;
wire \Mux16~1_combout ;
wire \Mux16~7_combout ;
wire \Mux16~8_combout ;
wire \Mux16~4_combout ;
wire \Mux16~5_combout ;
wire \Mux16~2_combout ;
wire \Mux16~3_combout ;
wire \Mux16~6_combout ;
wire \Mux16~17_combout ;
wire \Mux16~18_combout ;
wire \register[10][15]~q ;
wire \register[8][15]~q ;
wire \Mux16~10_combout ;
wire \Mux16~11_combout ;
wire \register[2][15]~q ;
wire \Mux16~15_combout ;
wire \Mux16~12_combout ;
wire \Mux16~13_combout ;
wire \Mux16~16_combout ;
wire \Mux17~4_combout ;
wire \Mux17~5_combout ;
wire \register[22][14]~q ;
wire \Mux17~2_combout ;
wire \Mux17~3_combout ;
wire \Mux17~6_combout ;
wire \register[19][14]~feeder_combout ;
wire \register[19][14]~q ;
wire \Mux17~7_combout ;
wire \Mux17~8_combout ;
wire \Mux17~0_combout ;
wire \Mux17~1_combout ;
wire \Mux17~17_combout ;
wire \Mux17~18_combout ;
wire \Mux17~15_combout ;
wire \Mux17~12_combout ;
wire \Mux17~13_combout ;
wire \Mux17~16_combout ;
wire \Mux17~10_combout ;
wire \Mux17~11_combout ;
wire \Mux18~7_combout ;
wire \Mux18~8_combout ;
wire \Mux18~2_combout ;
wire \Mux18~3_combout ;
wire \register[28][13]~q ;
wire \Mux18~4_combout ;
wire \Mux18~5_combout ;
wire \Mux18~6_combout ;
wire \register[25][13]~feeder_combout ;
wire \register[25][13]~q ;
wire \Mux18~0_combout ;
wire \Mux18~1_combout ;
wire \register[8][13]~q ;
wire \Mux18~10_combout ;
wire \register[11][13]~q ;
wire \Mux18~11_combout ;
wire \register[13][13]~q ;
wire \Mux18~17_combout ;
wire \Mux18~18_combout ;
wire \register[4][13]~q ;
wire \Mux18~12_combout ;
wire \Mux18~13_combout ;
wire \register[3][13]~q ;
wire \Mux18~14_combout ;
wire \Mux18~15_combout ;
wire \Mux18~16_combout ;
wire \Mux19~0_combout ;
wire \Mux19~1_combout ;
wire \Mux19~7_combout ;
wire \Mux19~8_combout ;
wire \Mux19~4_combout ;
wire \Mux19~5_combout ;
wire \Mux19~3_combout ;
wire \Mux19~6_combout ;
wire \Mux19~17_combout ;
wire \Mux19~18_combout ;
wire \register[4][12]~q ;
wire \Mux19~10_combout ;
wire \Mux19~11_combout ;
wire \Mux19~14_combout ;
wire \Mux19~15_combout ;
wire \Mux19~12_combout ;
wire \Mux19~13_combout ;
wire \Mux19~16_combout ;
wire \Mux20~7_combout ;
wire \Mux20~8_combout ;
wire \Mux20~0_combout ;
wire \Mux20~1_combout ;
wire \register[24][11]~q ;
wire \Mux20~4_combout ;
wire \Mux20~5_combout ;
wire \register[22][11]~feeder_combout ;
wire \register[22][11]~q ;
wire \Mux20~2_combout ;
wire \Mux20~3_combout ;
wire \Mux20~6_combout ;
wire \Mux20~17_combout ;
wire \Mux20~18_combout ;
wire \Mux20~14_combout ;
wire \Mux20~15_combout ;
wire \Mux20~12_combout ;
wire \Mux20~13_combout ;
wire \Mux20~16_combout ;
wire \Mux20~10_combout ;
wire \register[11][11]~q ;
wire \Mux20~11_combout ;
wire \register[17][10]~q ;
wire \Mux21~0_combout ;
wire \Mux21~1_combout ;
wire \register[22][10]~q ;
wire \Mux21~2_combout ;
wire \Mux21~3_combout ;
wire \register[20][10]~feeder_combout ;
wire \register[20][10]~q ;
wire \Mux21~4_combout ;
wire \Mux21~5_combout ;
wire \Mux21~6_combout ;
wire \Mux21~7_combout ;
wire \Mux21~8_combout ;
wire \register[6][10]~feeder_combout ;
wire \register[6][10]~q ;
wire \Mux21~10_combout ;
wire \Mux21~11_combout ;
wire \Mux21~17_combout ;
wire \Mux21~18_combout ;
wire \Mux21~13_combout ;
wire \Mux21~14_combout ;
wire \Mux21~15_combout ;
wire \Mux21~16_combout ;
wire \Mux22~7_combout ;
wire \Mux22~8_combout ;
wire \register[17][9]~q ;
wire \Mux22~0_combout ;
wire \Mux22~1_combout ;
wire \register[24][9]~feeder_combout ;
wire \register[24][9]~q ;
wire \Mux22~4_combout ;
wire \Mux22~5_combout ;
wire \register[22][9]~q ;
wire \register[30][9]~feeder_combout ;
wire \register[30][9]~q ;
wire \Mux22~3_combout ;
wire \Mux22~6_combout ;
wire \Mux22~17_combout ;
wire \Mux22~18_combout ;
wire \Mux22~10_combout ;
wire \Mux22~11_combout ;
wire \Mux22~14_combout ;
wire \Mux22~15_combout ;
wire \Mux22~12_combout ;
wire \Mux22~13_combout ;
wire \Mux22~16_combout ;
wire \register[17][4]~feeder_combout ;
wire \register[17][4]~q ;
wire \Mux59~0_combout ;
wire \Mux59~1_combout ;
wire \Mux59~7_combout ;
wire \Mux59~8_combout ;
wire \Mux59~2_combout ;
wire \register[22][4]~q ;
wire \Mux59~3_combout ;
wire \Mux59~4_combout ;
wire \Mux59~5_combout ;
wire \Mux59~6_combout ;
wire \Mux59~12_combout ;
wire \Mux59~13_combout ;
wire \register[2][4]~q ;
wire \Mux59~15_combout ;
wire \Mux59~16_combout ;
wire \Mux59~17_combout ;
wire \Mux59~18_combout ;
wire \Mux59~10_combout ;
wire \Mux59~11_combout ;
wire \Mux0~7_combout ;
wire \Mux0~8_combout ;
wire \register[17][31]~q ;
wire \Mux0~0_combout ;
wire \Mux0~1_combout ;
wire \register[20][31]~q ;
wire \Mux0~4_combout ;
wire \Mux0~5_combout ;
wire \Mux0~2_combout ;
wire \Mux0~3_combout ;
wire \Mux0~6_combout ;
wire \register[4][31]~q ;
wire \Mux0~12_combout ;
wire \Mux0~13_combout ;
wire \Mux0~14_combout ;
wire \Mux0~15_combout ;
wire \Mux0~16_combout ;
wire \register[11][31]~feeder_combout ;
wire \register[11][31]~q ;
wire \Mux0~10_combout ;
wire \Mux0~11_combout ;
wire \register[12][31]~q ;
wire \Mux0~17_combout ;
wire \Mux0~18_combout ;
wire \Mux2~0_combout ;
wire \Mux2~1_combout ;
wire \register[30][29]~q ;
wire \Mux2~3_combout ;
wire \register[24][29]~q ;
wire \Mux2~4_combout ;
wire \Mux2~5_combout ;
wire \Mux2~6_combout ;
wire \Mux2~7_combout ;
wire \Mux2~8_combout ;
wire \Mux2~17_combout ;
wire \Mux2~18_combout ;
wire \register[8][29]~q ;
wire \Mux2~10_combout ;
wire \Mux2~11_combout ;
wire \register[1][29]~q ;
wire \Mux2~14_combout ;
wire \Mux2~15_combout ;
wire \Mux2~13_combout ;
wire \Mux2~16_combout ;
wire \register[24][30]~q ;
wire \Mux1~4_combout ;
wire \Mux1~5_combout ;
wire \register[22][30]~q ;
wire \Mux1~2_combout ;
wire \register[26][30]~q ;
wire \Mux1~3_combout ;
wire \Mux1~6_combout ;
wire \register[17][30]~q ;
wire \Mux1~0_combout ;
wire \Mux1~1_combout ;
wire \Mux1~7_combout ;
wire \Mux1~8_combout ;
wire \register[4][30]~q ;
wire \Mux1~10_combout ;
wire \Mux1~11_combout ;
wire \Mux1~17_combout ;
wire \Mux1~18_combout ;
wire \Mux1~14_combout ;
wire \Mux1~15_combout ;
wire \Mux1~12_combout ;
wire \Mux1~13_combout ;
wire \Mux1~16_combout ;
wire \register[17][28]~feeder_combout ;
wire \register[17][28]~q ;
wire \Mux3~0_combout ;
wire \Mux3~1_combout ;
wire \Mux3~7_combout ;
wire \Mux3~8_combout ;
wire \Mux3~2_combout ;
wire \Mux3~3_combout ;
wire \register[16][28]~q ;
wire \Mux3~4_combout ;
wire \Mux3~5_combout ;
wire \Mux3~6_combout ;
wire \Mux3~12_combout ;
wire \Mux3~13_combout ;
wire \Mux3~15_combout ;
wire \Mux3~16_combout ;
wire \register[13][28]~q ;
wire \Mux3~17_combout ;
wire \Mux3~18_combout ;
wire \register[6][28]~q ;
wire \Mux3~10_combout ;
wire \Mux3~11_combout ;
wire \register[19][27]~q ;
wire \Mux4~7_combout ;
wire \Mux4~8_combout ;
wire \Mux4~0_combout ;
wire \Mux4~1_combout ;
wire \Mux4~4_combout ;
wire \Mux4~5_combout ;
wire \Mux4~2_combout ;
wire \Mux4~3_combout ;
wire \Mux4~6_combout ;
wire \register[4][27]~q ;
wire \Mux4~12_combout ;
wire \Mux4~13_combout ;
wire \register[2][27]~q ;
wire \Mux4~14_combout ;
wire \Mux4~15_combout ;
wire \Mux4~16_combout ;
wire \Mux4~10_combout ;
wire \Mux4~11_combout ;
wire \register[12][27]~q ;
wire \Mux4~17_combout ;
wire \Mux4~18_combout ;
wire \Mux5~7_combout ;
wire \Mux5~8_combout ;
wire \Mux5~0_combout ;
wire \Mux5~1_combout ;
wire \Mux5~2_combout ;
wire \Mux5~3_combout ;
wire \register[16][26]~q ;
wire \Mux5~4_combout ;
wire \Mux5~5_combout ;
wire \Mux5~6_combout ;
wire \Mux5~17_combout ;
wire \Mux5~18_combout ;
wire \Mux5~10_combout ;
wire \Mux5~11_combout ;
wire \register[2][26]~feeder_combout ;
wire \register[2][26]~q ;
wire \Mux5~14_combout ;
wire \Mux5~15_combout ;
wire \Mux5~12_combout ;
wire \Mux5~13_combout ;
wire \Mux5~16_combout ;
wire \Mux6~0_combout ;
wire \Mux6~1_combout ;
wire \Mux6~7_combout ;
wire \Mux6~8_combout ;
wire \Mux6~2_combout ;
wire \Mux6~3_combout ;
wire \register[24][25]~q ;
wire \register[16][25]~feeder_combout ;
wire \register[16][25]~q ;
wire \Mux6~4_combout ;
wire \Mux6~5_combout ;
wire \Mux6~6_combout ;
wire \Mux6~10_combout ;
wire \Mux6~11_combout ;
wire \register[4][25]~q ;
wire \Mux6~12_combout ;
wire \Mux6~13_combout ;
wire \Mux6~15_combout ;
wire \Mux6~16_combout ;
wire \register[13][25]~q ;
wire \Mux6~17_combout ;
wire \Mux6~18_combout ;
wire \Mux7~7_combout ;
wire \Mux7~8_combout ;
wire \register[28][24]~q ;
wire \Mux7~4_combout ;
wire \Mux7~5_combout ;
wire \register[18][24]~q ;
wire \Mux7~2_combout ;
wire \Mux7~3_combout ;
wire \Mux7~6_combout ;
wire \Mux7~0_combout ;
wire \register[21][24]~feeder_combout ;
wire \register[21][24]~q ;
wire \Mux7~1_combout ;
wire \register[5][24]~q ;
wire \Mux7~10_combout ;
wire \Mux7~11_combout ;
wire \Mux7~17_combout ;
wire \Mux7~18_combout ;
wire \Mux7~14_combout ;
wire \Mux7~15_combout ;
wire \Mux7~12_combout ;
wire \Mux7~13_combout ;
wire \Mux7~16_combout ;
wire \Mux8~7_combout ;
wire \Mux8~8_combout ;
wire \register[17][23]~feeder_combout ;
wire \register[17][23]~q ;
wire \Mux8~0_combout ;
wire \Mux8~1_combout ;
wire \register[18][23]~feeder_combout ;
wire \register[18][23]~q ;
wire \register[26][23]~q ;
wire \Mux8~2_combout ;
wire \Mux8~3_combout ;
wire \register[16][23]~feeder_combout ;
wire \register[16][23]~q ;
wire \Mux8~4_combout ;
wire \Mux8~5_combout ;
wire \Mux8~6_combout ;
wire \Mux8~17_combout ;
wire \Mux8~18_combout ;
wire \Mux8~10_combout ;
wire \Mux8~11_combout ;
wire \register[3][23]~q ;
wire \Mux8~14_combout ;
wire \Mux8~15_combout ;
wire \Mux8~12_combout ;
wire \Mux8~13_combout ;
wire \Mux8~16_combout ;
wire \Mux9~4_combout ;
wire \Mux9~5_combout ;
wire \Mux9~2_combout ;
wire \register[26][22]~q ;
wire \Mux9~3_combout ;
wire \Mux9~6_combout ;
wire \Mux9~7_combout ;
wire \register[23][22]~q ;
wire \Mux9~8_combout ;
wire \Mux9~0_combout ;
wire \Mux9~1_combout ;
wire \Mux9~10_combout ;
wire \register[6][22]~feeder_combout ;
wire \register[6][22]~q ;
wire \Mux9~11_combout ;
wire \Mux9~17_combout ;
wire \Mux9~18_combout ;
wire \Mux9~15_combout ;
wire \Mux9~13_combout ;
wire \Mux9~16_combout ;
wire \Mux10~7_combout ;
wire \Mux10~8_combout ;
wire \Mux10~0_combout ;
wire \Mux10~1_combout ;
wire \register[16][21]~feeder_combout ;
wire \register[16][21]~q ;
wire \Mux10~4_combout ;
wire \Mux10~5_combout ;
wire \Mux10~2_combout ;
wire \Mux10~3_combout ;
wire \Mux10~6_combout ;
wire \Mux10~17_combout ;
wire \Mux10~18_combout ;
wire \register[10][21]~q ;
wire \Mux10~10_combout ;
wire \Mux10~11_combout ;
wire \Mux10~13_combout ;
wire \Mux10~14_combout ;
wire \Mux10~15_combout ;
wire \Mux10~16_combout ;
wire \Mux11~7_combout ;
wire \Mux11~8_combout ;
wire \Mux11~0_combout ;
wire \Mux11~1_combout ;
wire \register[16][20]~q ;
wire \Mux11~4_combout ;
wire \Mux11~5_combout ;
wire \register[18][20]~q ;
wire \Mux11~2_combout ;
wire \Mux11~3_combout ;
wire \Mux11~6_combout ;
wire \register[8][20]~q ;
wire \Mux11~12_combout ;
wire \Mux11~13_combout ;
wire \Mux11~14_combout ;
wire \Mux11~15_combout ;
wire \Mux11~16_combout ;
wire \Mux11~17_combout ;
wire \Mux11~18_combout ;
wire \register[4][20]~q ;
wire \Mux11~10_combout ;
wire \Mux11~11_combout ;
wire \Mux12~0_combout ;
wire \Mux12~1_combout ;
wire \Mux12~7_combout ;
wire \register[27][19]~feeder_combout ;
wire \register[27][19]~q ;
wire \Mux12~8_combout ;
wire \register[18][19]~q ;
wire \Mux12~2_combout ;
wire \Mux12~3_combout ;
wire \Mux12~4_combout ;
wire \Mux12~5_combout ;
wire \Mux12~6_combout ;
wire \Mux12~17_combout ;
wire \Mux12~18_combout ;
wire \Mux12~13_combout ;
wire \register[2][19]~feeder_combout ;
wire \register[2][19]~q ;
wire \Mux12~14_combout ;
wire \Mux12~15_combout ;
wire \Mux12~16_combout ;
wire \Mux12~10_combout ;
wire \Mux12~11_combout ;
wire \Mux13~7_combout ;
wire \Mux13~8_combout ;
wire \Mux13~0_combout ;
wire \Mux13~1_combout ;
wire \Mux13~2_combout ;
wire \Mux13~3_combout ;
wire \register[28][18]~q ;
wire \Mux13~5_combout ;
wire \Mux13~6_combout ;
wire \Mux13~13_combout ;
wire \register[1][18]~q ;
wire \Mux13~14_combout ;
wire \Mux13~15_combout ;
wire \Mux13~16_combout ;
wire \register[4][18]~q ;
wire \register[5][18]~q ;
wire \Mux13~10_combout ;
wire \Mux13~11_combout ;
wire \Mux13~17_combout ;
wire \Mux13~18_combout ;
wire \register[19][17]~q ;
wire \Mux14~7_combout ;
wire \Mux14~8_combout ;
wire \Mux14~0_combout ;
wire \Mux14~1_combout ;
wire \register[22][17]~q ;
wire \register[26][17]~q ;
wire \Mux14~2_combout ;
wire \Mux14~3_combout ;
wire \Mux14~4_combout ;
wire \Mux14~5_combout ;
wire \Mux14~6_combout ;
wire \Mux14~17_combout ;
wire \Mux14~18_combout ;
wire \register[10][17]~q ;
wire \Mux14~10_combout ;
wire \Mux14~11_combout ;
wire \Mux14~14_combout ;
wire \Mux14~15_combout ;
wire \Mux14~12_combout ;
wire \Mux14~13_combout ;
wire \Mux14~16_combout ;
wire \Mux31~7_combout ;
wire \Mux31~8_combout ;
wire \Mux31~0_combout ;
wire \Mux31~1_combout ;
wire \Mux31~4_combout ;
wire \Mux31~5_combout ;
wire \register[22][0]~feeder_combout ;
wire \register[22][0]~q ;
wire \Mux31~2_combout ;
wire \Mux31~3_combout ;
wire \Mux31~6_combout ;
wire \Mux31~13_combout ;
wire \register[1][0]~q ;
wire \Mux31~14_combout ;
wire \Mux31~15_combout ;
wire \Mux31~16_combout ;
wire \Mux31~10_combout ;
wire \Mux31~11_combout ;
wire \Mux31~17_combout ;
wire \Mux31~18_combout ;


// Location: FF_X67_Y39_N29
dffeas \register[28][30] (
	.clk(!CLK),
	.d(\register[28][30]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~57_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\register[28][30]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \register[28][30] .is_wysiwyg = "true";
defparam \register[28][30] .power_up = "low";
// synopsys translate_on

// Location: FF_X69_Y33_N9
dffeas \register[3][29] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\register~66_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~48_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\register[3][29]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \register[3][29] .is_wysiwyg = "true";
defparam \register[3][29] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X69_Y33_N8
cycloneive_lcell_comb \Mux34~14 (
// Equation(s):
// \Mux34~14_combout  = (Selector9 & ((plif_ifidinstr_l_17 & (\register[3][29]~q )) # (!plif_ifidinstr_l_17 & ((\register[1][29]~q ))))) # (!Selector9 & (((\register[1][29]~q ))))

	.dataa(Selector9),
	.datab(plif_ifidinstr_l_17),
	.datac(\register[3][29]~q ),
	.datad(\register[1][29]~q ),
	.cin(gnd),
	.combout(\Mux34~14_combout ),
	.cout());
// synopsys translate_off
defparam \Mux34~14 .lut_mask = 16'hF780;
defparam \Mux34~14 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X67_Y39_N21
dffeas \register[30][28] (
	.clk(!CLK),
	.d(\register[30][28]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~56_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\register[30][28]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \register[30][28] .is_wysiwyg = "true";
defparam \register[30][28] .power_up = "low";
// synopsys translate_on

// Location: FF_X65_Y35_N21
dffeas \register[24][28] (
	.clk(!CLK),
	.d(\register[24][28]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~34_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\register[24][28]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \register[24][28] .is_wysiwyg = "true";
defparam \register[24][28] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X65_Y39_N16
cycloneive_lcell_comb \Mux35~4 (
// Equation(s):
// \Mux35~4_combout  = (Selector7 & ((\register[24][28]~q ) # ((Selector8)))) # (!Selector7 & (((\register[16][28]~q  & !Selector8))))

	.dataa(Selector7),
	.datab(\register[24][28]~q ),
	.datac(\register[16][28]~q ),
	.datad(Selector8),
	.cin(gnd),
	.combout(\Mux35~4_combout ),
	.cout());
// synopsys translate_off
defparam \Mux35~4 .lut_mask = 16'hAAD8;
defparam \Mux35~4 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X65_Y33_N21
dffeas \register[3][28] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\register~67_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~48_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\register[3][28]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \register[3][28] .is_wysiwyg = "true";
defparam \register[3][28] .power_up = "low";
// synopsys translate_on

// Location: FF_X65_Y33_N15
dffeas \register[1][28] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\register~67_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~49_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\register[1][28]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \register[1][28] .is_wysiwyg = "true";
defparam \register[1][28] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X65_Y33_N14
cycloneive_lcell_comb \Mux35~14 (
// Equation(s):
// \Mux35~14_combout  = (Selector10 & ((Selector91 & (\register[3][28]~q )) # (!Selector91 & ((\register[1][28]~q )))))

	.dataa(Selector91),
	.datab(\register[3][28]~q ),
	.datac(\register[1][28]~q ),
	.datad(Selector10),
	.cin(gnd),
	.combout(\Mux35~14_combout ),
	.cout());
// synopsys translate_off
defparam \Mux35~14 .lut_mask = 16'hD800;
defparam \Mux35~14 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X69_Y31_N31
dffeas \register[4][24] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\register~71_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~60_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\register[4][24]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \register[4][24] .is_wysiwyg = "true";
defparam \register[4][24] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X69_Y31_N30
cycloneive_lcell_comb \Mux39~12 (
// Equation(s):
// \Mux39~12_combout  = (Selector91 & (((Selector10)))) # (!Selector91 & ((Selector10 & (\register[5][24]~q )) # (!Selector10 & ((\register[4][24]~q )))))

	.dataa(Selector91),
	.datab(\register[5][24]~q ),
	.datac(\register[4][24]~q ),
	.datad(Selector10),
	.cin(gnd),
	.combout(\Mux39~12_combout ),
	.cout());
// synopsys translate_off
defparam \Mux39~12 .lut_mask = 16'hEE50;
defparam \Mux39~12 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X69_Y33_N31
dffeas \register[1][23] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\register~72_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~49_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\register[1][23]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \register[1][23] .is_wysiwyg = "true";
defparam \register[1][23] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X69_Y33_N30
cycloneive_lcell_comb \Mux40~14 (
// Equation(s):
// \Mux40~14_combout  = (Selector9 & ((plif_ifidinstr_l_17 & ((\register[3][23]~q ))) # (!plif_ifidinstr_l_17 & (\register[1][23]~q )))) # (!Selector9 & (((\register[1][23]~q ))))

	.dataa(Selector9),
	.datab(plif_ifidinstr_l_17),
	.datac(\register[1][23]~q ),
	.datad(\register[3][23]~q ),
	.cin(gnd),
	.combout(\Mux40~14_combout ),
	.cout());
// synopsys translate_off
defparam \Mux40~14 .lut_mask = 16'hF870;
defparam \Mux40~14 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X68_Y34_N27
dffeas \register[28][21] (
	.clk(!CLK),
	.d(\register[28][21]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~57_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\register[28][21]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \register[28][21] .is_wysiwyg = "true";
defparam \register[28][21] .power_up = "low";
// synopsys translate_on

// Location: FF_X67_Y32_N13
dffeas \register[5][21] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\register~74_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~59_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\register[5][21]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \register[5][21] .is_wysiwyg = "true";
defparam \register[5][21] .power_up = "low";
// synopsys translate_on

// Location: FF_X66_Y40_N27
dffeas \register[8][21] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\register~74_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~46_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\register[8][21]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \register[8][21] .is_wysiwyg = "true";
defparam \register[8][21] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X66_Y40_N26
cycloneive_lcell_comb \Mux42~12 (
// Equation(s):
// \Mux42~12_combout  = (Selector91 & ((Selector10) # ((\register[10][21]~q )))) # (!Selector91 & (!Selector10 & (\register[8][21]~q )))

	.dataa(Selector91),
	.datab(Selector10),
	.datac(\register[8][21]~q ),
	.datad(\register[10][21]~q ),
	.cin(gnd),
	.combout(\Mux42~12_combout ),
	.cout());
// synopsys translate_off
defparam \Mux42~12 .lut_mask = 16'hBA98;
defparam \Mux42~12 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X69_Y39_N11
dffeas \register[26][20] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\register~75_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~54_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\register[26][20]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \register[26][20] .is_wysiwyg = "true";
defparam \register[26][20] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X69_Y39_N10
cycloneive_lcell_comb \Mux43~2 (
// Equation(s):
// \Mux43~2_combout  = (Selector8 & (((Selector7)))) # (!Selector8 & ((Selector7 & ((\register[26][20]~q ))) # (!Selector7 & (\register[18][20]~q ))))

	.dataa(Selector8),
	.datab(\register[18][20]~q ),
	.datac(\register[26][20]~q ),
	.datad(Selector7),
	.cin(gnd),
	.combout(\Mux43~2_combout ),
	.cout());
// synopsys translate_off
defparam \Mux43~2 .lut_mask = 16'hFA44;
defparam \Mux43~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X66_Y39_N11
dffeas \register[24][20] (
	.clk(!CLK),
	.d(\register[24][20]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~34_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\register[24][20]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \register[24][20] .is_wysiwyg = "true";
defparam \register[24][20] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X65_Y39_N0
cycloneive_lcell_comb \Mux43~4 (
// Equation(s):
// \Mux43~4_combout  = (Selector7 & ((\register[24][20]~q ) # ((Selector8)))) # (!Selector7 & (((\register[16][20]~q  & !Selector8))))

	.dataa(Selector7),
	.datab(\register[24][20]~q ),
	.datac(\register[16][20]~q ),
	.datad(Selector8),
	.cin(gnd),
	.combout(\Mux43~4_combout ),
	.cout());
// synopsys translate_off
defparam \Mux43~4 .lut_mask = 16'hAAD8;
defparam \Mux43~4 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X67_Y32_N15
dffeas \register[4][19] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\register~76_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~60_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\register[4][19]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \register[4][19] .is_wysiwyg = "true";
defparam \register[4][19] .power_up = "low";
// synopsys translate_on

// Location: FF_X59_Y36_N11
dffeas \register[13][19] (
	.clk(!CLK),
	.d(\register[13][19]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~62_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\register[13][19]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \register[13][19] .is_wysiwyg = "true";
defparam \register[13][19] .power_up = "low";
// synopsys translate_on

// Location: FF_X66_Y40_N31
dffeas \register[8][18] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\register~77_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~46_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\register[8][18]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \register[8][18] .is_wysiwyg = "true";
defparam \register[8][18] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X67_Y32_N4
cycloneive_lcell_comb \Mux45~12 (
// Equation(s):
// \Mux45~12_combout  = (Selector91 & (((Selector10)))) # (!Selector91 & ((Selector10 & ((\register[5][18]~q ))) # (!Selector10 & (\register[4][18]~q ))))

	.dataa(\register[4][18]~q ),
	.datab(Selector91),
	.datac(\register[5][18]~q ),
	.datad(Selector10),
	.cin(gnd),
	.combout(\Mux45~12_combout ),
	.cout());
// synopsys translate_off
defparam \Mux45~12 .lut_mask = 16'hFC22;
defparam \Mux45~12 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X59_Y36_N13
dffeas \register[13][18] (
	.clk(!CLK),
	.d(\register[13][18]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~62_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\register[13][18]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \register[13][18] .is_wysiwyg = "true";
defparam \register[13][18] .power_up = "low";
// synopsys translate_on

// Location: FF_X61_Y40_N11
dffeas \register[28][17] (
	.clk(!CLK),
	.d(\register[28][17]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~57_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\register[28][17]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \register[28][17] .is_wysiwyg = "true";
defparam \register[28][17] .power_up = "low";
// synopsys translate_on

// Location: FF_X66_Y40_N1
dffeas \register[8][17] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\register~78_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~46_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\register[8][17]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \register[8][17] .is_wysiwyg = "true";
defparam \register[8][17] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X66_Y40_N0
cycloneive_lcell_comb \Mux46~12 (
// Equation(s):
// \Mux46~12_combout  = (Selector91 & ((Selector10) # ((\register[10][17]~q )))) # (!Selector91 & (!Selector10 & (\register[8][17]~q )))

	.dataa(Selector91),
	.datab(Selector10),
	.datac(\register[8][17]~q ),
	.datad(\register[10][17]~q ),
	.cin(gnd),
	.combout(\Mux46~12_combout ),
	.cout());
// synopsys translate_off
defparam \Mux46~12 .lut_mask = 16'hBA98;
defparam \Mux46~12 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X67_Y37_N11
dffeas \register[18][16] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\register~79_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~33_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\register[18][16]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \register[18][16] .is_wysiwyg = "true";
defparam \register[18][16] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X67_Y37_N10
cycloneive_lcell_comb \Mux47~2 (
// Equation(s):
// \Mux47~2_combout  = (Selector8 & (((Selector7)))) # (!Selector8 & ((Selector7 & (\register[26][16]~q )) # (!Selector7 & ((\register[18][16]~q )))))

	.dataa(Selector8),
	.datab(\register[26][16]~q ),
	.datac(\register[18][16]~q ),
	.datad(Selector7),
	.cin(gnd),
	.combout(\Mux47~2_combout ),
	.cout());
// synopsys translate_off
defparam \Mux47~2 .lut_mask = 16'hEE50;
defparam \Mux47~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y40_N16
cycloneive_lcell_comb \Mux48~12 (
// Equation(s):
// \Mux48~12_combout  = (Selector91 & (((\register[10][15]~q ) # (Selector10)))) # (!Selector91 & (\register[8][15]~q  & ((!Selector10))))

	.dataa(\register[8][15]~q ),
	.datab(Selector91),
	.datac(\register[10][15]~q ),
	.datad(Selector10),
	.cin(gnd),
	.combout(\Mux48~12_combout ),
	.cout());
// synopsys translate_off
defparam \Mux48~12 .lut_mask = 16'hCCE2;
defparam \Mux48~12 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X68_Y39_N27
dffeas \register[22][13] (
	.clk(!CLK),
	.d(\register[22][13]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~55_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\register[22][13]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \register[22][13] .is_wysiwyg = "true";
defparam \register[22][13] .power_up = "low";
// synopsys translate_on

// Location: FF_X69_Y37_N7
dffeas \register[22][12] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\register~83_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~55_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\register[22][12]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \register[22][12] .is_wysiwyg = "true";
defparam \register[22][12] .power_up = "low";
// synopsys translate_on

// Location: FF_X62_Y41_N13
dffeas \register[10][10] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\register~85_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~45_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\register[10][10]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \register[10][10] .is_wysiwyg = "true";
defparam \register[10][10] .power_up = "low";
// synopsys translate_on

// Location: FF_X68_Y37_N27
dffeas \register[26][8] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\register~87_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~54_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\register[26][8]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \register[26][8] .is_wysiwyg = "true";
defparam \register[26][8] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X68_Y37_N26
cycloneive_lcell_comb \Mux55~2 (
// Equation(s):
// \Mux55~2_combout  = (Selector7 & (((\register[26][8]~q ) # (Selector8)))) # (!Selector7 & (\register[18][8]~q  & ((!Selector8))))

	.dataa(Selector7),
	.datab(\register[18][8]~q ),
	.datac(\register[26][8]~q ),
	.datad(Selector8),
	.cin(gnd),
	.combout(\Mux55~2_combout ),
	.cout());
// synopsys translate_off
defparam \Mux55~2 .lut_mask = 16'hAAE4;
defparam \Mux55~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X65_Y39_N31
dffeas \register[20][8] (
	.clk(!CLK),
	.d(\register[20][8]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~35_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\register[20][8]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \register[20][8] .is_wysiwyg = "true";
defparam \register[20][8] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X67_Y38_N20
cycloneive_lcell_comb \Mux56~12 (
// Equation(s):
// \Mux56~12_combout  = (Selector10 & (Selector91)) # (!Selector10 & ((Selector91 & (\register[10][7]~q )) # (!Selector91 & ((\register[8][7]~q )))))

	.dataa(Selector10),
	.datab(Selector91),
	.datac(\register[10][7]~q ),
	.datad(\register[8][7]~q ),
	.cin(gnd),
	.combout(\Mux56~12_combout ),
	.cout());
// synopsys translate_off
defparam \Mux56~12 .lut_mask = 16'hD9C8;
defparam \Mux56~12 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X69_Y37_N21
dffeas \register[18][6] (
	.clk(!CLK),
	.d(\register[18][6]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~33_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\register[18][6]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \register[18][6] .is_wysiwyg = "true";
defparam \register[18][6] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X68_Y37_N22
cycloneive_lcell_comb \Mux57~2 (
// Equation(s):
// \Mux57~2_combout  = (Selector7 & ((Selector8) # ((\register[26][6]~q )))) # (!Selector7 & (!Selector8 & ((\register[18][6]~q ))))

	.dataa(Selector7),
	.datab(Selector8),
	.datac(\register[26][6]~q ),
	.datad(\register[18][6]~q ),
	.cin(gnd),
	.combout(\Mux57~2_combout ),
	.cout());
// synopsys translate_off
defparam \Mux57~2 .lut_mask = 16'hB9A8;
defparam \Mux57~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X70_Y38_N13
dffeas \register[16][5] (
	.clk(!CLK),
	.d(\register[16][5]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~36_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\register[16][5]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \register[16][5] .is_wysiwyg = "true";
defparam \register[16][5] .power_up = "low";
// synopsys translate_on

// Location: FF_X67_Y39_N1
dffeas \register[28][5] (
	.clk(!CLK),
	.d(\register[28][5]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~57_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\register[28][5]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \register[28][5] .is_wysiwyg = "true";
defparam \register[28][5] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X62_Y40_N8
cycloneive_lcell_comb \Mux58~12 (
// Equation(s):
// \Mux58~12_combout  = (Selector91 & (((\register[10][5]~q ) # (Selector10)))) # (!Selector91 & (\register[8][5]~q  & ((!Selector10))))

	.dataa(Selector91),
	.datab(\register[8][5]~q ),
	.datac(\register[10][5]~q ),
	.datad(Selector10),
	.cin(gnd),
	.combout(\Mux58~12_combout ),
	.cout());
// synopsys translate_off
defparam \Mux58~12 .lut_mask = 16'hAAE4;
defparam \Mux58~12 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X70_Y34_N5
dffeas \register[3][2] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\register~91_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~48_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\register[3][2]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \register[3][2] .is_wysiwyg = "true";
defparam \register[3][2] .power_up = "low";
// synopsys translate_on

// Location: FF_X70_Y34_N19
dffeas \register[1][2] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\register~91_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~49_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\register[1][2]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \register[1][2] .is_wysiwyg = "true";
defparam \register[1][2] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X70_Y34_N18
cycloneive_lcell_comb \Mux29~14 (
// Equation(s):
// \Mux29~14_combout  = (Selector4 & ((plif_ifidinstr_l_22 & (\register[3][2]~q )) # (!plif_ifidinstr_l_22 & ((\register[1][2]~q ))))) # (!Selector4 & (((\register[1][2]~q ))))

	.dataa(Selector4),
	.datab(\register[3][2]~q ),
	.datac(\register[1][2]~q ),
	.datad(plif_ifidinstr_l_22),
	.cin(gnd),
	.combout(\Mux29~14_combout ),
	.cout());
// synopsys translate_off
defparam \Mux29~14 .lut_mask = 16'hD8F0;
defparam \Mux29~14 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X70_Y35_N13
dffeas \register[24][1] (
	.clk(!CLK),
	.d(\register[24][1]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~34_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\register[24][1]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \register[24][1] .is_wysiwyg = "true";
defparam \register[24][1] .power_up = "low";
// synopsys translate_on

// Location: FF_X66_Y36_N7
dffeas \register[20][0] (
	.clk(!CLK),
	.d(\register[20][0]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~35_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\register[20][0]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \register[20][0] .is_wysiwyg = "true";
defparam \register[20][0] .power_up = "low";
// synopsys translate_on

// Location: FF_X63_Y41_N23
dffeas \register[8][0] (
	.clk(!CLK),
	.d(\register[8][0]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~46_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\register[8][0]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \register[8][0] .is_wysiwyg = "true";
defparam \register[8][0] .power_up = "low";
// synopsys translate_on

// Location: FF_X66_Y33_N23
dffeas \register[28][4] (
	.clk(!CLK),
	.d(\register[28][4]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~57_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\register[28][4]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \register[28][4] .is_wysiwyg = "true";
defparam \register[28][4] .power_up = "low";
// synopsys translate_on

// Location: FF_X70_Y34_N13
dffeas \register[3][4] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\register~94_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~48_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\register[3][4]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \register[3][4] .is_wysiwyg = "true";
defparam \register[3][4] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X70_Y34_N4
cycloneive_lcell_comb \Mux61~14 (
// Equation(s):
// \Mux61~14_combout  = (Selector10 & ((Selector91 & ((\register[3][2]~q ))) # (!Selector91 & (\register[1][2]~q ))))

	.dataa(Selector91),
	.datab(\register[1][2]~q ),
	.datac(\register[3][2]~q ),
	.datad(Selector10),
	.cin(gnd),
	.combout(\Mux61~14_combout ),
	.cout());
// synopsys translate_off
defparam \Mux61~14 .lut_mask = 16'hE400;
defparam \Mux61~14 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X70_Y38_N20
cycloneive_lcell_comb \Mux24~4 (
// Equation(s):
// \Mux24~4_combout  = (Selector3 & (((Selector2)))) # (!Selector3 & ((Selector2 & (\register[24][7]~q )) # (!Selector2 & ((\register[16][7]~q )))))

	.dataa(Selector3),
	.datab(\register[24][7]~q ),
	.datac(Selector2),
	.datad(\register[16][7]~q ),
	.cin(gnd),
	.combout(\Mux24~4_combout ),
	.cout());
// synopsys translate_off
defparam \Mux24~4 .lut_mask = 16'hE5E0;
defparam \Mux24~4 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X69_Y37_N30
cycloneive_lcell_comb \Mux25~2 (
// Equation(s):
// \Mux25~2_combout  = (Selector2 & (((Selector3)))) # (!Selector2 & ((Selector3 & ((\register[22][6]~q ))) # (!Selector3 & (\register[18][6]~q ))))

	.dataa(Selector2),
	.datab(\register[18][6]~q ),
	.datac(\register[22][6]~q ),
	.datad(Selector3),
	.cin(gnd),
	.combout(\Mux25~2_combout ),
	.cout());
// synopsys translate_off
defparam \Mux25~2 .lut_mask = 16'hFA44;
defparam \Mux25~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X70_Y34_N20
cycloneive_lcell_comb \Mux60~14 (
// Equation(s):
// \Mux60~14_combout  = (Selector10 & ((Selector91 & ((\register[3][3]~q ))) # (!Selector91 & (\register[1][3]~q ))))

	.dataa(\register[1][3]~q ),
	.datab(Selector91),
	.datac(\register[3][3]~q ),
	.datad(Selector10),
	.cin(gnd),
	.combout(\Mux60~14_combout ),
	.cout());
// synopsys translate_off
defparam \Mux60~14 .lut_mask = 16'hE200;
defparam \Mux60~14 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X65_Y37_N16
cycloneive_lcell_comb \Mux15~4 (
// Equation(s):
// \Mux15~4_combout  = (Selector3 & (((\register[20][16]~q ) # (Selector2)))) # (!Selector3 & (\register[16][16]~q  & ((!Selector2))))

	.dataa(Selector3),
	.datab(\register[16][16]~q ),
	.datac(\register[20][16]~q ),
	.datad(Selector2),
	.cin(gnd),
	.combout(\Mux15~4_combout ),
	.cout());
// synopsys translate_off
defparam \Mux15~4 .lut_mask = 16'hAAE4;
defparam \Mux15~4 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X65_Y33_N0
cycloneive_lcell_comb \Mux16~14 (
// Equation(s):
// \Mux16~14_combout  = (Selector5 & ((Selector41 & ((\register[3][15]~q ))) # (!Selector41 & (\register[1][15]~q ))))

	.dataa(\register[1][15]~q ),
	.datab(Selector5),
	.datac(\register[3][15]~q ),
	.datad(Selector41),
	.cin(gnd),
	.combout(\Mux16~14_combout ),
	.cout());
// synopsys translate_off
defparam \Mux16~14 .lut_mask = 16'hC088;
defparam \Mux16~14 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X70_Y34_N16
cycloneive_lcell_comb \Mux17~14 (
// Equation(s):
// \Mux17~14_combout  = (Selector4 & ((plif_ifidinstr_l_22 & ((\register[3][14]~q ))) # (!plif_ifidinstr_l_22 & (\register[1][14]~q )))) # (!Selector4 & (\register[1][14]~q ))

	.dataa(Selector4),
	.datab(\register[1][14]~q ),
	.datac(\register[3][14]~q ),
	.datad(plif_ifidinstr_l_22),
	.cin(gnd),
	.combout(\Mux17~14_combout ),
	.cout());
// synopsys translate_off
defparam \Mux17~14 .lut_mask = 16'hE4CC;
defparam \Mux17~14 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X69_Y37_N6
cycloneive_lcell_comb \Mux19~2 (
// Equation(s):
// \Mux19~2_combout  = (Selector2 & (((Selector3)))) # (!Selector2 & ((Selector3 & ((\register[22][12]~q ))) # (!Selector3 & (\register[18][12]~q ))))

	.dataa(Selector2),
	.datab(\register[18][12]~q ),
	.datac(\register[22][12]~q ),
	.datad(Selector3),
	.cin(gnd),
	.combout(\Mux19~2_combout ),
	.cout());
// synopsys translate_off
defparam \Mux19~2 .lut_mask = 16'hFA44;
defparam \Mux19~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y41_N12
cycloneive_lcell_comb \Mux21~12 (
// Equation(s):
// \Mux21~12_combout  = (Selector41 & (((\register[10][10]~q ) # (Selector5)))) # (!Selector41 & (\register[8][10]~q  & ((!Selector5))))

	.dataa(Selector41),
	.datab(\register[8][10]~q ),
	.datac(\register[10][10]~q ),
	.datad(Selector5),
	.cin(gnd),
	.combout(\Mux21~12_combout ),
	.cout());
// synopsys translate_off
defparam \Mux21~12 .lut_mask = 16'hAAE4;
defparam \Mux21~12 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X68_Y37_N16
cycloneive_lcell_comb \Mux22~2 (
// Equation(s):
// \Mux22~2_combout  = (Selector2 & ((Selector3) # ((\register[26][9]~q )))) # (!Selector2 & (!Selector3 & ((\register[18][9]~q ))))

	.dataa(Selector2),
	.datab(Selector3),
	.datac(\register[26][9]~q ),
	.datad(\register[18][9]~q ),
	.cin(gnd),
	.combout(\Mux22~2_combout ),
	.cout());
// synopsys translate_off
defparam \Mux22~2 .lut_mask = 16'hB9A8;
defparam \Mux22~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X70_Y34_N12
cycloneive_lcell_comb \Mux59~14 (
// Equation(s):
// \Mux59~14_combout  = (Selector10 & ((Selector91 & (\register[3][4]~q )) # (!Selector91 & ((\register[1][4]~q )))))

	.dataa(Selector10),
	.datab(Selector91),
	.datac(\register[3][4]~q ),
	.datad(\register[1][4]~q ),
	.cin(gnd),
	.combout(\Mux59~14_combout ),
	.cout());
// synopsys translate_off
defparam \Mux59~14 .lut_mask = 16'hA280;
defparam \Mux59~14 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X69_Y35_N6
cycloneive_lcell_comb \Mux2~2 (
// Equation(s):
// \Mux2~2_combout  = (Selector3 & (((Selector2)))) # (!Selector3 & ((Selector2 & (\register[26][29]~q )) # (!Selector2 & ((\register[18][29]~q )))))

	.dataa(\register[26][29]~q ),
	.datab(Selector3),
	.datac(\register[18][29]~q ),
	.datad(Selector2),
	.cin(gnd),
	.combout(\Mux2~2_combout ),
	.cout());
// synopsys translate_off
defparam \Mux2~2 .lut_mask = 16'hEE30;
defparam \Mux2~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X69_Y31_N12
cycloneive_lcell_comb \Mux2~12 (
// Equation(s):
// \Mux2~12_combout  = (Selector5 & (((\register[5][29]~q ) # (Selector41)))) # (!Selector5 & (\register[4][29]~q  & ((!Selector41))))

	.dataa(Selector5),
	.datab(\register[4][29]~q ),
	.datac(\register[5][29]~q ),
	.datad(Selector41),
	.cin(gnd),
	.combout(\Mux2~12_combout ),
	.cout());
// synopsys translate_off
defparam \Mux2~12 .lut_mask = 16'hAAE4;
defparam \Mux2~12 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X65_Y33_N20
cycloneive_lcell_comb \Mux3~14 (
// Equation(s):
// \Mux3~14_combout  = (Selector5 & ((Selector41 & ((\register[3][28]~q ))) # (!Selector41 & (\register[1][28]~q ))))

	.dataa(\register[1][28]~q ),
	.datab(Selector5),
	.datac(\register[3][28]~q ),
	.datad(Selector41),
	.cin(gnd),
	.combout(\Mux3~14_combout ),
	.cout());
// synopsys translate_off
defparam \Mux3~14 .lut_mask = 16'hC088;
defparam \Mux3~14 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X65_Y36_N28
cycloneive_lcell_comb \Mux6~14 (
// Equation(s):
// \Mux6~14_combout  = (plif_ifidinstr_l_22 & ((Selector4 & ((\register[3][25]~q ))) # (!Selector4 & (\register[1][25]~q )))) # (!plif_ifidinstr_l_22 & (\register[1][25]~q ))

	.dataa(\register[1][25]~q ),
	.datab(plif_ifidinstr_l_22),
	.datac(\register[3][25]~q ),
	.datad(Selector4),
	.cin(gnd),
	.combout(\Mux6~14_combout ),
	.cout());
// synopsys translate_off
defparam \Mux6~14 .lut_mask = 16'hE2AA;
defparam \Mux6~14 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y40_N14
cycloneive_lcell_comb \Mux9~12 (
// Equation(s):
// \Mux9~12_combout  = (Selector41 & ((Selector5) # ((\register[10][22]~q )))) # (!Selector41 & (!Selector5 & (\register[8][22]~q )))

	.dataa(Selector41),
	.datab(Selector5),
	.datac(\register[8][22]~q ),
	.datad(\register[10][22]~q ),
	.cin(gnd),
	.combout(\Mux9~12_combout ),
	.cout());
// synopsys translate_off
defparam \Mux9~12 .lut_mask = 16'hBA98;
defparam \Mux9~12 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X69_Y33_N4
cycloneive_lcell_comb \Mux9~14 (
// Equation(s):
// \Mux9~14_combout  = (Selector4 & ((plif_ifidinstr_l_22 & (\register[3][22]~q )) # (!plif_ifidinstr_l_22 & ((\register[1][22]~q ))))) # (!Selector4 & (((\register[1][22]~q ))))

	.dataa(Selector4),
	.datab(plif_ifidinstr_l_22),
	.datac(\register[3][22]~q ),
	.datad(\register[1][22]~q ),
	.cin(gnd),
	.combout(\Mux9~14_combout ),
	.cout());
// synopsys translate_off
defparam \Mux9~14 .lut_mask = 16'hF780;
defparam \Mux9~14 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X67_Y32_N12
cycloneive_lcell_comb \Mux10~12 (
// Equation(s):
// \Mux10~12_combout  = (Selector41 & (Selector5)) # (!Selector41 & ((Selector5 & (\register[5][21]~q )) # (!Selector5 & ((\register[4][21]~q )))))

	.dataa(Selector41),
	.datab(Selector5),
	.datac(\register[5][21]~q ),
	.datad(\register[4][21]~q ),
	.cin(gnd),
	.combout(\Mux10~12_combout ),
	.cout());
// synopsys translate_off
defparam \Mux10~12 .lut_mask = 16'hD9C8;
defparam \Mux10~12 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X67_Y32_N14
cycloneive_lcell_comb \Mux12~12 (
// Equation(s):
// \Mux12~12_combout  = (Selector41 & (Selector5)) # (!Selector41 & ((Selector5 & ((\register[5][19]~q ))) # (!Selector5 & (\register[4][19]~q ))))

	.dataa(Selector41),
	.datab(Selector5),
	.datac(\register[4][19]~q ),
	.datad(\register[5][19]~q ),
	.cin(gnd),
	.combout(\Mux12~12_combout ),
	.cout());
// synopsys translate_off
defparam \Mux12~12 .lut_mask = 16'hDC98;
defparam \Mux12~12 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X65_Y39_N2
cycloneive_lcell_comb \Mux13~4 (
// Equation(s):
// \Mux13~4_combout  = (Selector2 & (((Selector3)))) # (!Selector2 & ((Selector3 & ((\register[20][18]~q ))) # (!Selector3 & (\register[16][18]~q ))))

	.dataa(Selector2),
	.datab(\register[16][18]~q ),
	.datac(\register[20][18]~q ),
	.datad(Selector3),
	.cin(gnd),
	.combout(\Mux13~4_combout ),
	.cout());
// synopsys translate_off
defparam \Mux13~4 .lut_mask = 16'hFA44;
defparam \Mux13~4 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X66_Y40_N30
cycloneive_lcell_comb \Mux13~12 (
// Equation(s):
// \Mux13~12_combout  = (Selector5 & (((Selector41)))) # (!Selector5 & ((Selector41 & (\register[10][18]~q )) # (!Selector41 & ((\register[8][18]~q )))))

	.dataa(\register[10][18]~q ),
	.datab(Selector5),
	.datac(\register[8][18]~q ),
	.datad(Selector41),
	.cin(gnd),
	.combout(\Mux13~12_combout ),
	.cout());
// synopsys translate_off
defparam \Mux13~12 .lut_mask = 16'hEE30;
defparam \Mux13~12 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X63_Y41_N30
cycloneive_lcell_comb \Mux31~12 (
// Equation(s):
// \Mux31~12_combout  = (Selector5 & (((Selector41)))) # (!Selector5 & ((Selector41 & ((\register[10][0]~q ))) # (!Selector41 & (\register[8][0]~q ))))

	.dataa(\register[8][0]~q ),
	.datab(\register[10][0]~q ),
	.datac(Selector5),
	.datad(Selector41),
	.cin(gnd),
	.combout(\Mux31~12_combout ),
	.cout());
// synopsys translate_off
defparam \Mux31~12 .lut_mask = 16'hFC0A;
defparam \Mux31~12 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X67_Y39_N28
cycloneive_lcell_comb \register[28][30]~feeder (
// Equation(s):
// \register[28][30]~feeder_combout  = \register~65_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(\register~65_combout ),
	.cin(gnd),
	.combout(\register[28][30]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \register[28][30]~feeder .lut_mask = 16'hFF00;
defparam \register[28][30]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X67_Y39_N20
cycloneive_lcell_comb \register[30][28]~feeder (
// Equation(s):
// \register[30][28]~feeder_combout  = \register~67_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(\register~67_combout ),
	.datad(gnd),
	.cin(gnd),
	.combout(\register[30][28]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \register[30][28]~feeder .lut_mask = 16'hF0F0;
defparam \register[30][28]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X65_Y35_N20
cycloneive_lcell_comb \register[24][28]~feeder (
// Equation(s):
// \register[24][28]~feeder_combout  = \register~67_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(\register~67_combout ),
	.cin(gnd),
	.combout(\register[24][28]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \register[24][28]~feeder .lut_mask = 16'hFF00;
defparam \register[24][28]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X68_Y34_N26
cycloneive_lcell_comb \register[28][21]~feeder (
// Equation(s):
// \register[28][21]~feeder_combout  = \register~74_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(\register~74_combout ),
	.cin(gnd),
	.combout(\register[28][21]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \register[28][21]~feeder .lut_mask = 16'hFF00;
defparam \register[28][21]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X66_Y39_N10
cycloneive_lcell_comb \register[24][20]~feeder (
// Equation(s):
// \register[24][20]~feeder_combout  = \register~75_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(\register~75_combout ),
	.datad(gnd),
	.cin(gnd),
	.combout(\register[24][20]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \register[24][20]~feeder .lut_mask = 16'hF0F0;
defparam \register[24][20]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y36_N10
cycloneive_lcell_comb \register[13][19]~feeder (
// Equation(s):
// \register[13][19]~feeder_combout  = \register~76_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(\register~76_combout ),
	.cin(gnd),
	.combout(\register[13][19]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \register[13][19]~feeder .lut_mask = 16'hFF00;
defparam \register[13][19]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y36_N12
cycloneive_lcell_comb \register[13][18]~feeder (
// Equation(s):
// \register[13][18]~feeder_combout  = \register~77_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(\register~77_combout ),
	.datad(gnd),
	.cin(gnd),
	.combout(\register[13][18]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \register[13][18]~feeder .lut_mask = 16'hF0F0;
defparam \register[13][18]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y40_N10
cycloneive_lcell_comb \register[28][17]~feeder (
// Equation(s):
// \register[28][17]~feeder_combout  = \register~78_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(\register~78_combout ),
	.datad(gnd),
	.cin(gnd),
	.combout(\register[28][17]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \register[28][17]~feeder .lut_mask = 16'hF0F0;
defparam \register[28][17]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X68_Y39_N26
cycloneive_lcell_comb \register[22][13]~feeder (
// Equation(s):
// \register[22][13]~feeder_combout  = \register~82_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(\register~82_combout ),
	.datad(gnd),
	.cin(gnd),
	.combout(\register[22][13]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \register[22][13]~feeder .lut_mask = 16'hF0F0;
defparam \register[22][13]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X65_Y39_N30
cycloneive_lcell_comb \register[20][8]~feeder (
// Equation(s):
// \register[20][8]~feeder_combout  = \register~87_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(\register~87_combout ),
	.cin(gnd),
	.combout(\register[20][8]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \register[20][8]~feeder .lut_mask = 16'hFF00;
defparam \register[20][8]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X69_Y37_N20
cycloneive_lcell_comb \register[18][6]~feeder (
// Equation(s):
// \register[18][6]~feeder_combout  = \register~89_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(\register~89_combout ),
	.datad(gnd),
	.cin(gnd),
	.combout(\register[18][6]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \register[18][6]~feeder .lut_mask = 16'hF0F0;
defparam \register[18][6]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X67_Y39_N0
cycloneive_lcell_comb \register[28][5]~feeder (
// Equation(s):
// \register[28][5]~feeder_combout  = \register~90_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(\register~90_combout ),
	.cin(gnd),
	.combout(\register[28][5]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \register[28][5]~feeder .lut_mask = 16'hFF00;
defparam \register[28][5]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X70_Y38_N12
cycloneive_lcell_comb \register[16][5]~feeder (
// Equation(s):
// \register[16][5]~feeder_combout  = \register~90_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(\register~90_combout ),
	.datad(gnd),
	.cin(gnd),
	.combout(\register[16][5]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \register[16][5]~feeder .lut_mask = 16'hF0F0;
defparam \register[16][5]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X70_Y35_N12
cycloneive_lcell_comb \register[24][1]~feeder (
// Equation(s):
// \register[24][1]~feeder_combout  = \register~92_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(\register~92_combout ),
	.datad(gnd),
	.cin(gnd),
	.combout(\register[24][1]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \register[24][1]~feeder .lut_mask = 16'hF0F0;
defparam \register[24][1]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X63_Y41_N22
cycloneive_lcell_comb \register[8][0]~feeder (
// Equation(s):
// \register[8][0]~feeder_combout  = \register~93_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(\register~93_combout ),
	.cin(gnd),
	.combout(\register[8][0]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \register[8][0]~feeder .lut_mask = 16'hFF00;
defparam \register[8][0]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X66_Y36_N6
cycloneive_lcell_comb \register[20][0]~feeder (
// Equation(s):
// \register[20][0]~feeder_combout  = \register~93_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(\register~93_combout ),
	.cin(gnd),
	.combout(\register[20][0]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \register[20][0]~feeder .lut_mask = 16'hFF00;
defparam \register[20][0]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X66_Y33_N22
cycloneive_lcell_comb \register[28][4]~feeder (
// Equation(s):
// \register[28][4]~feeder_combout  = \register~94_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(\register~94_combout ),
	.datad(gnd),
	.cin(gnd),
	.combout(\register[28][4]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \register[28][4]~feeder .lut_mask = 16'hF0F0;
defparam \register[28][4]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y37_N2
cycloneive_lcell_comb \Decoder0~20 (
// Equation(s):
// Decoder0 = (!plif_memwbwsel_l_2 & !plif_memwbwsel_l_1)

	.dataa(gnd),
	.datab(gnd),
	.datac(plif_memwbwsel_l_2),
	.datad(plif_memwbwsel_l_1),
	.cin(gnd),
	.combout(Decoder0),
	.cout());
// synopsys translate_off
defparam \Decoder0~20 .lut_mask = 16'h000F;
defparam \Decoder0~20 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X67_Y35_N0
cycloneive_lcell_comb \Mux32~9 (
// Equation(s):
// Mux32 = (Selector10 & ((\Mux32~6_combout  & (\Mux32~8_combout )) # (!\Mux32~6_combout  & ((\Mux32~1_combout ))))) # (!Selector10 & (((\Mux32~6_combout ))))

	.dataa(\Mux32~8_combout ),
	.datab(Selector10),
	.datac(\Mux32~1_combout ),
	.datad(\Mux32~6_combout ),
	.cin(gnd),
	.combout(Mux32),
	.cout());
// synopsys translate_off
defparam \Mux32~9 .lut_mask = 16'hBBC0;
defparam \Mux32~9 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X67_Y35_N26
cycloneive_lcell_comb \Mux32~19 (
// Equation(s):
// Mux321 = (Selector8 & ((\Mux32~16_combout  & ((\Mux32~18_combout ))) # (!\Mux32~16_combout  & (\Mux32~11_combout )))) # (!Selector8 & (((\Mux32~16_combout ))))

	.dataa(Selector8),
	.datab(\Mux32~11_combout ),
	.datac(\Mux32~18_combout ),
	.datad(\Mux32~16_combout ),
	.cin(gnd),
	.combout(Mux321),
	.cout());
// synopsys translate_off
defparam \Mux32~19 .lut_mask = 16'hF588;
defparam \Mux32~19 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y39_N2
cycloneive_lcell_comb \Mux33~9 (
// Equation(s):
// Mux33 = (\Mux33~6_combout  & ((\Mux33~8_combout ) # ((!Selector10)))) # (!\Mux33~6_combout  & (((\Mux33~1_combout  & Selector10))))

	.dataa(\Mux33~6_combout ),
	.datab(\Mux33~8_combout ),
	.datac(\Mux33~1_combout ),
	.datad(Selector10),
	.cin(gnd),
	.combout(Mux33),
	.cout());
// synopsys translate_off
defparam \Mux33~9 .lut_mask = 16'hD8AA;
defparam \Mux33~9 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y39_N20
cycloneive_lcell_comb \Mux33~19 (
// Equation(s):
// Mux331 = (Selector7 & ((\Mux33~16_combout  & (\Mux33~18_combout )) # (!\Mux33~16_combout  & ((\Mux33~11_combout ))))) # (!Selector7 & (((\Mux33~16_combout ))))

	.dataa(Selector7),
	.datab(\Mux33~18_combout ),
	.datac(\Mux33~11_combout ),
	.datad(\Mux33~16_combout ),
	.cin(gnd),
	.combout(Mux331),
	.cout());
// synopsys translate_off
defparam \Mux33~19 .lut_mask = 16'hDDA0;
defparam \Mux33~19 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y32_N26
cycloneive_lcell_comb \Mux34~9 (
// Equation(s):
// Mux34 = (Selector10 & ((\Mux34~6_combout  & (\Mux34~8_combout )) # (!\Mux34~6_combout  & ((\Mux34~1_combout ))))) # (!Selector10 & (((\Mux34~6_combout ))))

	.dataa(\Mux34~8_combout ),
	.datab(Selector10),
	.datac(\Mux34~1_combout ),
	.datad(\Mux34~6_combout ),
	.cin(gnd),
	.combout(Mux34),
	.cout());
// synopsys translate_off
defparam \Mux34~9 .lut_mask = 16'hBBC0;
defparam \Mux34~9 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y32_N18
cycloneive_lcell_comb \Mux34~19 (
// Equation(s):
// Mux341 = (Selector8 & ((\Mux34~16_combout  & (\Mux34~18_combout )) # (!\Mux34~16_combout  & ((\Mux34~11_combout ))))) # (!Selector8 & (((\Mux34~16_combout ))))

	.dataa(\Mux34~18_combout ),
	.datab(Selector8),
	.datac(\Mux34~11_combout ),
	.datad(\Mux34~16_combout ),
	.cin(gnd),
	.combout(Mux341),
	.cout());
// synopsys translate_off
defparam \Mux34~19 .lut_mask = 16'hBBC0;
defparam \Mux34~19 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X67_Y35_N18
cycloneive_lcell_comb \Mux35~9 (
// Equation(s):
// Mux35 = (Selector10 & ((\Mux35~6_combout  & (\Mux35~8_combout )) # (!\Mux35~6_combout  & ((\Mux35~1_combout ))))) # (!Selector10 & (((\Mux35~6_combout ))))

	.dataa(Selector10),
	.datab(\Mux35~8_combout ),
	.datac(\Mux35~1_combout ),
	.datad(\Mux35~6_combout ),
	.cin(gnd),
	.combout(Mux35),
	.cout());
// synopsys translate_off
defparam \Mux35~9 .lut_mask = 16'hDDA0;
defparam \Mux35~9 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X67_Y35_N22
cycloneive_lcell_comb \Mux35~19 (
// Equation(s):
// Mux351 = (Selector7 & ((\Mux35~16_combout  & (\Mux35~18_combout )) # (!\Mux35~16_combout  & ((\Mux35~11_combout ))))) # (!Selector7 & (((\Mux35~16_combout ))))

	.dataa(\Mux35~18_combout ),
	.datab(Selector7),
	.datac(\Mux35~16_combout ),
	.datad(\Mux35~11_combout ),
	.cin(gnd),
	.combout(Mux351),
	.cout());
// synopsys translate_off
defparam \Mux35~19 .lut_mask = 16'hBCB0;
defparam \Mux35~19 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y39_N14
cycloneive_lcell_comb \Mux36~9 (
// Equation(s):
// Mux36 = (Selector10 & ((\Mux36~6_combout  & (\Mux36~8_combout )) # (!\Mux36~6_combout  & ((\Mux36~1_combout ))))) # (!Selector10 & (((\Mux36~6_combout ))))

	.dataa(\Mux36~8_combout ),
	.datab(Selector10),
	.datac(\Mux36~1_combout ),
	.datad(\Mux36~6_combout ),
	.cin(gnd),
	.combout(Mux36),
	.cout());
// synopsys translate_off
defparam \Mux36~9 .lut_mask = 16'hBBC0;
defparam \Mux36~9 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y39_N0
cycloneive_lcell_comb \Mux36~19 (
// Equation(s):
// Mux361 = (Selector8 & ((\Mux36~16_combout  & ((\Mux36~18_combout ))) # (!\Mux36~16_combout  & (\Mux36~11_combout )))) # (!Selector8 & (((\Mux36~16_combout ))))

	.dataa(Selector8),
	.datab(\Mux36~11_combout ),
	.datac(\Mux36~18_combout ),
	.datad(\Mux36~16_combout ),
	.cin(gnd),
	.combout(Mux361),
	.cout());
// synopsys translate_off
defparam \Mux36~19 .lut_mask = 16'hF588;
defparam \Mux36~19 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y32_N0
cycloneive_lcell_comb \Mux37~9 (
// Equation(s):
// Mux37 = (Selector10 & ((\Mux37~6_combout  & ((\Mux37~8_combout ))) # (!\Mux37~6_combout  & (\Mux37~1_combout )))) # (!Selector10 & (((\Mux37~6_combout ))))

	.dataa(Selector10),
	.datab(\Mux37~1_combout ),
	.datac(\Mux37~8_combout ),
	.datad(\Mux37~6_combout ),
	.cin(gnd),
	.combout(Mux37),
	.cout());
// synopsys translate_off
defparam \Mux37~9 .lut_mask = 16'hF588;
defparam \Mux37~9 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y32_N14
cycloneive_lcell_comb \Mux37~19 (
// Equation(s):
// Mux371 = (Selector7 & ((\Mux37~16_combout  & ((\Mux37~18_combout ))) # (!\Mux37~16_combout  & (\Mux37~11_combout )))) # (!Selector7 & (((\Mux37~16_combout ))))

	.dataa(\Mux37~11_combout ),
	.datab(Selector7),
	.datac(\Mux37~16_combout ),
	.datad(\Mux37~18_combout ),
	.cin(gnd),
	.combout(Mux371),
	.cout());
// synopsys translate_off
defparam \Mux37~19 .lut_mask = 16'hF838;
defparam \Mux37~19 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X65_Y32_N2
cycloneive_lcell_comb \Mux38~9 (
// Equation(s):
// Mux38 = (Selector10 & ((\Mux38~6_combout  & ((\Mux38~8_combout ))) # (!\Mux38~6_combout  & (\Mux38~1_combout )))) # (!Selector10 & (((\Mux38~6_combout ))))

	.dataa(Selector10),
	.datab(\Mux38~1_combout ),
	.datac(\Mux38~8_combout ),
	.datad(\Mux38~6_combout ),
	.cin(gnd),
	.combout(Mux38),
	.cout());
// synopsys translate_off
defparam \Mux38~9 .lut_mask = 16'hF588;
defparam \Mux38~9 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X65_Y32_N14
cycloneive_lcell_comb \Mux38~19 (
// Equation(s):
// Mux381 = (Selector8 & ((\Mux38~16_combout  & (\Mux38~18_combout )) # (!\Mux38~16_combout  & ((\Mux38~11_combout ))))) # (!Selector8 & (((\Mux38~16_combout ))))

	.dataa(\Mux38~18_combout ),
	.datab(Selector8),
	.datac(\Mux38~11_combout ),
	.datad(\Mux38~16_combout ),
	.cin(gnd),
	.combout(Mux381),
	.cout());
// synopsys translate_off
defparam \Mux38~19 .lut_mask = 16'hBBC0;
defparam \Mux38~19 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X65_Y34_N4
cycloneive_lcell_comb \Mux39~9 (
// Equation(s):
// Mux39 = (Selector10 & ((\Mux39~6_combout  & ((\Mux39~8_combout ))) # (!\Mux39~6_combout  & (\Mux39~1_combout )))) # (!Selector10 & (((\Mux39~6_combout ))))

	.dataa(\Mux39~1_combout ),
	.datab(Selector10),
	.datac(\Mux39~6_combout ),
	.datad(\Mux39~8_combout ),
	.cin(gnd),
	.combout(Mux39),
	.cout());
// synopsys translate_off
defparam \Mux39~9 .lut_mask = 16'hF838;
defparam \Mux39~9 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X65_Y32_N0
cycloneive_lcell_comb \Mux39~19 (
// Equation(s):
// Mux391 = (\Mux39~16_combout  & (((\Mux39~18_combout )) # (!Selector7))) # (!\Mux39~16_combout  & (Selector7 & ((\Mux39~11_combout ))))

	.dataa(\Mux39~16_combout ),
	.datab(Selector7),
	.datac(\Mux39~18_combout ),
	.datad(\Mux39~11_combout ),
	.cin(gnd),
	.combout(Mux391),
	.cout());
// synopsys translate_off
defparam \Mux39~19 .lut_mask = 16'hE6A2;
defparam \Mux39~19 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X67_Y30_N4
cycloneive_lcell_comb \Mux40~9 (
// Equation(s):
// Mux40 = (Selector10 & ((\Mux40~6_combout  & (\Mux40~8_combout )) # (!\Mux40~6_combout  & ((\Mux40~1_combout ))))) # (!Selector10 & (((\Mux40~6_combout ))))

	.dataa(\Mux40~8_combout ),
	.datab(Selector10),
	.datac(\Mux40~1_combout ),
	.datad(\Mux40~6_combout ),
	.cin(gnd),
	.combout(Mux40),
	.cout());
// synopsys translate_off
defparam \Mux40~9 .lut_mask = 16'hBBC0;
defparam \Mux40~9 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X67_Y30_N20
cycloneive_lcell_comb \Mux40~19 (
// Equation(s):
// Mux401 = (Selector8 & ((\Mux40~16_combout  & (\Mux40~18_combout )) # (!\Mux40~16_combout  & ((\Mux40~11_combout ))))) # (!Selector8 & (\Mux40~16_combout ))

	.dataa(Selector8),
	.datab(\Mux40~16_combout ),
	.datac(\Mux40~18_combout ),
	.datad(\Mux40~11_combout ),
	.cin(gnd),
	.combout(Mux401),
	.cout());
// synopsys translate_off
defparam \Mux40~19 .lut_mask = 16'hE6C4;
defparam \Mux40~19 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X67_Y30_N28
cycloneive_lcell_comb \Mux41~9 (
// Equation(s):
// Mux41 = (Selector10 & ((\Mux41~6_combout  & ((\Mux41~8_combout ))) # (!\Mux41~6_combout  & (\Mux41~1_combout )))) # (!Selector10 & (((\Mux41~6_combout ))))

	.dataa(Selector10),
	.datab(\Mux41~1_combout ),
	.datac(\Mux41~6_combout ),
	.datad(\Mux41~8_combout ),
	.cin(gnd),
	.combout(Mux41),
	.cout());
// synopsys translate_off
defparam \Mux41~9 .lut_mask = 16'hF858;
defparam \Mux41~9 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X67_Y30_N12
cycloneive_lcell_comb \Mux41~19 (
// Equation(s):
// Mux411 = (\Mux41~16_combout  & ((\Mux41~18_combout ) # ((!Selector7)))) # (!\Mux41~16_combout  & (((Selector7 & \Mux41~11_combout ))))

	.dataa(\Mux41~18_combout ),
	.datab(\Mux41~16_combout ),
	.datac(Selector7),
	.datad(\Mux41~11_combout ),
	.cin(gnd),
	.combout(Mux411),
	.cout());
// synopsys translate_off
defparam \Mux41~19 .lut_mask = 16'hBC8C;
defparam \Mux41~19 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X68_Y34_N24
cycloneive_lcell_comb \Mux42~9 (
// Equation(s):
// Mux42 = (Selector10 & ((\Mux42~6_combout  & ((\Mux42~8_combout ))) # (!\Mux42~6_combout  & (\Mux42~1_combout )))) # (!Selector10 & (\Mux42~6_combout ))

	.dataa(Selector10),
	.datab(\Mux42~6_combout ),
	.datac(\Mux42~1_combout ),
	.datad(\Mux42~8_combout ),
	.cin(gnd),
	.combout(Mux42),
	.cout());
// synopsys translate_off
defparam \Mux42~9 .lut_mask = 16'hEC64;
defparam \Mux42~9 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X68_Y34_N22
cycloneive_lcell_comb \Mux42~19 (
// Equation(s):
// Mux421 = (\Mux42~16_combout  & ((\Mux42~18_combout ) # ((!Selector8)))) # (!\Mux42~16_combout  & (((\Mux42~11_combout  & Selector8))))

	.dataa(\Mux42~18_combout ),
	.datab(\Mux42~11_combout ),
	.datac(\Mux42~16_combout ),
	.datad(Selector8),
	.cin(gnd),
	.combout(Mux421),
	.cout());
// synopsys translate_off
defparam \Mux42~19 .lut_mask = 16'hACF0;
defparam \Mux42~19 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y39_N26
cycloneive_lcell_comb \Mux43~9 (
// Equation(s):
// Mux43 = (\Mux43~6_combout  & (((\Mux43~8_combout )) # (!Selector10))) # (!\Mux43~6_combout  & (Selector10 & ((\Mux43~1_combout ))))

	.dataa(\Mux43~6_combout ),
	.datab(Selector10),
	.datac(\Mux43~8_combout ),
	.datad(\Mux43~1_combout ),
	.cin(gnd),
	.combout(Mux43),
	.cout());
// synopsys translate_off
defparam \Mux43~9 .lut_mask = 16'hE6A2;
defparam \Mux43~9 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y39_N28
cycloneive_lcell_comb \Mux43~19 (
// Equation(s):
// Mux431 = (\Mux43~16_combout  & (((\Mux43~18_combout )) # (!Selector7))) # (!\Mux43~16_combout  & (Selector7 & (\Mux43~11_combout )))

	.dataa(\Mux43~16_combout ),
	.datab(Selector7),
	.datac(\Mux43~11_combout ),
	.datad(\Mux43~18_combout ),
	.cin(gnd),
	.combout(Mux431),
	.cout());
// synopsys translate_off
defparam \Mux43~19 .lut_mask = 16'hEA62;
defparam \Mux43~19 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y39_N16
cycloneive_lcell_comb \Mux44~9 (
// Equation(s):
// Mux44 = (Selector10 & ((\Mux44~6_combout  & (\Mux44~8_combout )) # (!\Mux44~6_combout  & ((\Mux44~1_combout ))))) # (!Selector10 & (((\Mux44~6_combout ))))

	.dataa(\Mux44~8_combout ),
	.datab(Selector10),
	.datac(\Mux44~1_combout ),
	.datad(\Mux44~6_combout ),
	.cin(gnd),
	.combout(Mux44),
	.cout());
// synopsys translate_off
defparam \Mux44~9 .lut_mask = 16'hBBC0;
defparam \Mux44~9 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y39_N4
cycloneive_lcell_comb \Mux44~19 (
// Equation(s):
// Mux441 = (Selector8 & ((\Mux44~16_combout  & (\Mux44~18_combout )) # (!\Mux44~16_combout  & ((\Mux44~11_combout ))))) # (!Selector8 & (((\Mux44~16_combout ))))

	.dataa(\Mux44~18_combout ),
	.datab(\Mux44~11_combout ),
	.datac(Selector8),
	.datad(\Mux44~16_combout ),
	.cin(gnd),
	.combout(Mux441),
	.cout());
// synopsys translate_off
defparam \Mux44~19 .lut_mask = 16'hAFC0;
defparam \Mux44~19 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X66_Y39_N24
cycloneive_lcell_comb \Mux45~9 (
// Equation(s):
// Mux45 = (\Mux45~6_combout  & (((\Mux45~8_combout )) # (!Selector10))) # (!\Mux45~6_combout  & (Selector10 & (\Mux45~1_combout )))

	.dataa(\Mux45~6_combout ),
	.datab(Selector10),
	.datac(\Mux45~1_combout ),
	.datad(\Mux45~8_combout ),
	.cin(gnd),
	.combout(Mux45),
	.cout());
// synopsys translate_off
defparam \Mux45~9 .lut_mask = 16'hEA62;
defparam \Mux45~9 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X66_Y39_N12
cycloneive_lcell_comb \Mux45~19 (
// Equation(s):
// Mux451 = (Selector7 & ((\Mux45~16_combout  & ((\Mux45~18_combout ))) # (!\Mux45~16_combout  & (\Mux45~11_combout )))) # (!Selector7 & (((\Mux45~16_combout ))))

	.dataa(Selector7),
	.datab(\Mux45~11_combout ),
	.datac(\Mux45~18_combout ),
	.datad(\Mux45~16_combout ),
	.cin(gnd),
	.combout(Mux451),
	.cout());
// synopsys translate_off
defparam \Mux45~19 .lut_mask = 16'hF588;
defparam \Mux45~19 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X67_Y40_N20
cycloneive_lcell_comb \Mux46~9 (
// Equation(s):
// Mux46 = (Selector10 & ((\Mux46~6_combout  & (\Mux46~8_combout )) # (!\Mux46~6_combout  & ((\Mux46~1_combout ))))) # (!Selector10 & (\Mux46~6_combout ))

	.dataa(Selector10),
	.datab(\Mux46~6_combout ),
	.datac(\Mux46~8_combout ),
	.datad(\Mux46~1_combout ),
	.cin(gnd),
	.combout(Mux46),
	.cout());
// synopsys translate_off
defparam \Mux46~9 .lut_mask = 16'hE6C4;
defparam \Mux46~9 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X67_Y40_N14
cycloneive_lcell_comb \Mux46~19 (
// Equation(s):
// Mux461 = (Selector8 & ((\Mux46~16_combout  & ((\Mux46~18_combout ))) # (!\Mux46~16_combout  & (\Mux46~11_combout )))) # (!Selector8 & (((\Mux46~16_combout ))))

	.dataa(Selector8),
	.datab(\Mux46~11_combout ),
	.datac(\Mux46~18_combout ),
	.datad(\Mux46~16_combout ),
	.cin(gnd),
	.combout(Mux461),
	.cout());
// synopsys translate_off
defparam \Mux46~19 .lut_mask = 16'hF588;
defparam \Mux46~19 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X67_Y40_N10
cycloneive_lcell_comb \Mux47~9 (
// Equation(s):
// Mux47 = (Selector10 & ((\Mux47~6_combout  & (\Mux47~8_combout )) # (!\Mux47~6_combout  & ((\Mux47~1_combout ))))) # (!Selector10 & (((\Mux47~6_combout ))))

	.dataa(Selector10),
	.datab(\Mux47~8_combout ),
	.datac(\Mux47~6_combout ),
	.datad(\Mux47~1_combout ),
	.cin(gnd),
	.combout(Mux47),
	.cout());
// synopsys translate_off
defparam \Mux47~9 .lut_mask = 16'hDAD0;
defparam \Mux47~9 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X67_Y40_N26
cycloneive_lcell_comb \Mux47~19 (
// Equation(s):
// Mux471 = (Selector7 & ((\Mux47~16_combout  & ((\Mux47~18_combout ))) # (!\Mux47~16_combout  & (\Mux47~11_combout )))) # (!Selector7 & (((\Mux47~16_combout ))))

	.dataa(\Mux47~11_combout ),
	.datab(Selector7),
	.datac(\Mux47~18_combout ),
	.datad(\Mux47~16_combout ),
	.cin(gnd),
	.combout(Mux471),
	.cout());
// synopsys translate_off
defparam \Mux47~19 .lut_mask = 16'hF388;
defparam \Mux47~19 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X70_Y35_N10
cycloneive_lcell_comb \Mux48~9 (
// Equation(s):
// Mux48 = (Selector10 & ((\Mux48~6_combout  & (\Mux48~8_combout )) # (!\Mux48~6_combout  & ((\Mux48~1_combout ))))) # (!Selector10 & (\Mux48~6_combout ))

	.dataa(Selector10),
	.datab(\Mux48~6_combout ),
	.datac(\Mux48~8_combout ),
	.datad(\Mux48~1_combout ),
	.cin(gnd),
	.combout(Mux48),
	.cout());
// synopsys translate_off
defparam \Mux48~9 .lut_mask = 16'hE6C4;
defparam \Mux48~9 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X70_Y35_N14
cycloneive_lcell_comb \Mux48~19 (
// Equation(s):
// Mux481 = (Selector8 & ((\Mux48~16_combout  & ((\Mux48~18_combout ))) # (!\Mux48~16_combout  & (\Mux48~11_combout )))) # (!Selector8 & (((\Mux48~16_combout ))))

	.dataa(Selector8),
	.datab(\Mux48~11_combout ),
	.datac(\Mux48~18_combout ),
	.datad(\Mux48~16_combout ),
	.cin(gnd),
	.combout(Mux481),
	.cout());
// synopsys translate_off
defparam \Mux48~19 .lut_mask = 16'hF588;
defparam \Mux48~19 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X66_Y30_N30
cycloneive_lcell_comb \Mux49~9 (
// Equation(s):
// Mux49 = (Selector10 & ((\Mux49~6_combout  & (\Mux49~8_combout )) # (!\Mux49~6_combout  & ((\Mux49~1_combout ))))) # (!Selector10 & (((\Mux49~6_combout ))))

	.dataa(Selector10),
	.datab(\Mux49~8_combout ),
	.datac(\Mux49~1_combout ),
	.datad(\Mux49~6_combout ),
	.cin(gnd),
	.combout(Mux49),
	.cout());
// synopsys translate_off
defparam \Mux49~9 .lut_mask = 16'hDDA0;
defparam \Mux49~9 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X66_Y30_N26
cycloneive_lcell_comb \Mux49~19 (
// Equation(s):
// Mux491 = (\Mux49~16_combout  & (((\Mux49~18_combout )) # (!Selector7))) # (!\Mux49~16_combout  & (Selector7 & (\Mux49~11_combout )))

	.dataa(\Mux49~16_combout ),
	.datab(Selector7),
	.datac(\Mux49~11_combout ),
	.datad(\Mux49~18_combout ),
	.cin(gnd),
	.combout(Mux491),
	.cout());
// synopsys translate_off
defparam \Mux49~19 .lut_mask = 16'hEA62;
defparam \Mux49~19 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X65_Y38_N16
cycloneive_lcell_comb \Mux50~9 (
// Equation(s):
// Mux50 = (Selector10 & ((\Mux50~6_combout  & ((\Mux50~8_combout ))) # (!\Mux50~6_combout  & (\Mux50~1_combout )))) # (!Selector10 & (((\Mux50~6_combout ))))

	.dataa(\Mux50~1_combout ),
	.datab(\Mux50~8_combout ),
	.datac(Selector10),
	.datad(\Mux50~6_combout ),
	.cin(gnd),
	.combout(Mux50),
	.cout());
// synopsys translate_off
defparam \Mux50~9 .lut_mask = 16'hCFA0;
defparam \Mux50~9 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X65_Y36_N10
cycloneive_lcell_comb \Mux50~19 (
// Equation(s):
// Mux501 = (Selector8 & ((\Mux50~16_combout  & (\Mux50~18_combout )) # (!\Mux50~16_combout  & ((\Mux50~11_combout ))))) # (!Selector8 & (((\Mux50~16_combout ))))

	.dataa(\Mux50~18_combout ),
	.datab(\Mux50~11_combout ),
	.datac(Selector8),
	.datad(\Mux50~16_combout ),
	.cin(gnd),
	.combout(Mux501),
	.cout());
// synopsys translate_off
defparam \Mux50~19 .lut_mask = 16'hAFC0;
defparam \Mux50~19 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y30_N16
cycloneive_lcell_comb \Mux51~9 (
// Equation(s):
// Mux51 = (Selector10 & ((\Mux51~6_combout  & (\Mux51~8_combout )) # (!\Mux51~6_combout  & ((\Mux51~1_combout ))))) # (!Selector10 & (((\Mux51~6_combout ))))

	.dataa(\Mux51~8_combout ),
	.datab(Selector10),
	.datac(\Mux51~1_combout ),
	.datad(\Mux51~6_combout ),
	.cin(gnd),
	.combout(Mux51),
	.cout());
// synopsys translate_off
defparam \Mux51~9 .lut_mask = 16'hBBC0;
defparam \Mux51~9 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y30_N26
cycloneive_lcell_comb \Mux51~19 (
// Equation(s):
// Mux511 = (Selector7 & ((\Mux51~16_combout  & ((\Mux51~18_combout ))) # (!\Mux51~16_combout  & (\Mux51~11_combout )))) # (!Selector7 & (((\Mux51~16_combout ))))

	.dataa(Selector7),
	.datab(\Mux51~11_combout ),
	.datac(\Mux51~18_combout ),
	.datad(\Mux51~16_combout ),
	.cin(gnd),
	.combout(Mux511),
	.cout());
// synopsys translate_off
defparam \Mux51~19 .lut_mask = 16'hF588;
defparam \Mux51~19 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y40_N4
cycloneive_lcell_comb \Mux52~9 (
// Equation(s):
// Mux52 = (Selector10 & ((\Mux52~6_combout  & ((\Mux52~8_combout ))) # (!\Mux52~6_combout  & (\Mux52~1_combout )))) # (!Selector10 & (((\Mux52~6_combout ))))

	.dataa(\Mux52~1_combout ),
	.datab(\Mux52~8_combout ),
	.datac(Selector10),
	.datad(\Mux52~6_combout ),
	.cin(gnd),
	.combout(Mux52),
	.cout());
// synopsys translate_off
defparam \Mux52~9 .lut_mask = 16'hCFA0;
defparam \Mux52~9 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X66_Y33_N6
cycloneive_lcell_comb \Mux52~19 (
// Equation(s):
// Mux521 = (Selector8 & ((\Mux52~16_combout  & ((\Mux52~18_combout ))) # (!\Mux52~16_combout  & (\Mux52~11_combout )))) # (!Selector8 & (((\Mux52~16_combout ))))

	.dataa(Selector8),
	.datab(\Mux52~11_combout ),
	.datac(\Mux52~18_combout ),
	.datad(\Mux52~16_combout ),
	.cin(gnd),
	.combout(Mux521),
	.cout());
// synopsys translate_off
defparam \Mux52~19 .lut_mask = 16'hF588;
defparam \Mux52~19 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X68_Y40_N8
cycloneive_lcell_comb \Mux53~9 (
// Equation(s):
// Mux53 = (Selector10 & ((\Mux53~6_combout  & (\Mux53~8_combout )) # (!\Mux53~6_combout  & ((\Mux53~1_combout ))))) # (!Selector10 & (\Mux53~6_combout ))

	.dataa(Selector10),
	.datab(\Mux53~6_combout ),
	.datac(\Mux53~8_combout ),
	.datad(\Mux53~1_combout ),
	.cin(gnd),
	.combout(Mux53),
	.cout());
// synopsys translate_off
defparam \Mux53~9 .lut_mask = 16'hE6C4;
defparam \Mux53~9 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X68_Y40_N12
cycloneive_lcell_comb \Mux53~19 (
// Equation(s):
// Mux531 = (Selector7 & ((\Mux53~16_combout  & ((\Mux53~18_combout ))) # (!\Mux53~16_combout  & (\Mux53~11_combout )))) # (!Selector7 & (((\Mux53~16_combout ))))

	.dataa(Selector7),
	.datab(\Mux53~11_combout ),
	.datac(\Mux53~18_combout ),
	.datad(\Mux53~16_combout ),
	.cin(gnd),
	.combout(Mux531),
	.cout());
// synopsys translate_off
defparam \Mux53~19 .lut_mask = 16'hF588;
defparam \Mux53~19 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X68_Y40_N2
cycloneive_lcell_comb \Mux54~9 (
// Equation(s):
// Mux54 = (Selector10 & ((\Mux54~6_combout  & (\Mux54~8_combout )) # (!\Mux54~6_combout  & ((\Mux54~1_combout ))))) # (!Selector10 & (\Mux54~6_combout ))

	.dataa(Selector10),
	.datab(\Mux54~6_combout ),
	.datac(\Mux54~8_combout ),
	.datad(\Mux54~1_combout ),
	.cin(gnd),
	.combout(Mux54),
	.cout());
// synopsys translate_off
defparam \Mux54~9 .lut_mask = 16'hE6C4;
defparam \Mux54~9 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X68_Y40_N22
cycloneive_lcell_comb \Mux54~19 (
// Equation(s):
// Mux541 = (Selector8 & ((\Mux54~16_combout  & (\Mux54~18_combout )) # (!\Mux54~16_combout  & ((\Mux54~11_combout ))))) # (!Selector8 & (((\Mux54~16_combout ))))

	.dataa(\Mux54~18_combout ),
	.datab(Selector8),
	.datac(\Mux54~11_combout ),
	.datad(\Mux54~16_combout ),
	.cin(gnd),
	.combout(Mux541),
	.cout());
// synopsys translate_off
defparam \Mux54~19 .lut_mask = 16'hBBC0;
defparam \Mux54~19 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X69_Y36_N28
cycloneive_lcell_comb \Mux55~9 (
// Equation(s):
// Mux55 = (Selector10 & ((\Mux55~6_combout  & ((\Mux55~8_combout ))) # (!\Mux55~6_combout  & (\Mux55~1_combout )))) # (!Selector10 & (((\Mux55~6_combout ))))

	.dataa(Selector10),
	.datab(\Mux55~1_combout ),
	.datac(\Mux55~6_combout ),
	.datad(\Mux55~8_combout ),
	.cin(gnd),
	.combout(Mux55),
	.cout());
// synopsys translate_off
defparam \Mux55~9 .lut_mask = 16'hF858;
defparam \Mux55~9 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X66_Y33_N26
cycloneive_lcell_comb \Mux55~19 (
// Equation(s):
// Mux551 = (Selector7 & ((\Mux55~16_combout  & (\Mux55~18_combout )) # (!\Mux55~16_combout  & ((\Mux55~11_combout ))))) # (!Selector7 & (((\Mux55~16_combout ))))

	.dataa(Selector7),
	.datab(\Mux55~18_combout ),
	.datac(\Mux55~11_combout ),
	.datad(\Mux55~16_combout ),
	.cin(gnd),
	.combout(Mux551),
	.cout());
// synopsys translate_off
defparam \Mux55~19 .lut_mask = 16'hDDA0;
defparam \Mux55~19 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X66_Y35_N18
cycloneive_lcell_comb \Mux56~9 (
// Equation(s):
// Mux56 = (Selector10 & ((\Mux56~6_combout  & (\Mux56~8_combout )) # (!\Mux56~6_combout  & ((\Mux56~1_combout ))))) # (!Selector10 & (((\Mux56~6_combout ))))

	.dataa(\Mux56~8_combout ),
	.datab(Selector10),
	.datac(\Mux56~1_combout ),
	.datad(\Mux56~6_combout ),
	.cin(gnd),
	.combout(Mux56),
	.cout());
// synopsys translate_off
defparam \Mux56~9 .lut_mask = 16'hBBC0;
defparam \Mux56~9 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X67_Y39_N4
cycloneive_lcell_comb \Mux56~19 (
// Equation(s):
// Mux561 = (Selector8 & ((\Mux56~16_combout  & ((\Mux56~18_combout ))) # (!\Mux56~16_combout  & (\Mux56~11_combout )))) # (!Selector8 & (\Mux56~16_combout ))

	.dataa(Selector8),
	.datab(\Mux56~16_combout ),
	.datac(\Mux56~11_combout ),
	.datad(\Mux56~18_combout ),
	.cin(gnd),
	.combout(Mux561),
	.cout());
// synopsys translate_off
defparam \Mux56~19 .lut_mask = 16'hEC64;
defparam \Mux56~19 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X65_Y30_N6
cycloneive_lcell_comb \Mux57~9 (
// Equation(s):
// Mux57 = (Selector10 & ((\Mux57~6_combout  & (\Mux57~8_combout )) # (!\Mux57~6_combout  & ((\Mux57~1_combout ))))) # (!Selector10 & (((\Mux57~6_combout ))))

	.dataa(Selector10),
	.datab(\Mux57~8_combout ),
	.datac(\Mux57~6_combout ),
	.datad(\Mux57~1_combout ),
	.cin(gnd),
	.combout(Mux57),
	.cout());
// synopsys translate_off
defparam \Mux57~9 .lut_mask = 16'hDAD0;
defparam \Mux57~9 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X65_Y30_N30
cycloneive_lcell_comb \Mux57~19 (
// Equation(s):
// Mux571 = (Selector7 & ((\Mux57~16_combout  & ((\Mux57~18_combout ))) # (!\Mux57~16_combout  & (\Mux57~11_combout )))) # (!Selector7 & (((\Mux57~16_combout ))))

	.dataa(Selector7),
	.datab(\Mux57~11_combout ),
	.datac(\Mux57~16_combout ),
	.datad(\Mux57~18_combout ),
	.cin(gnd),
	.combout(Mux571),
	.cout());
// synopsys translate_off
defparam \Mux57~19 .lut_mask = 16'hF858;
defparam \Mux57~19 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X65_Y30_N0
cycloneive_lcell_comb \Mux58~9 (
// Equation(s):
// Mux58 = (Selector10 & ((\Mux58~6_combout  & (\Mux58~8_combout )) # (!\Mux58~6_combout  & ((\Mux58~1_combout ))))) # (!Selector10 & (((\Mux58~6_combout ))))

	.dataa(Selector10),
	.datab(\Mux58~8_combout ),
	.datac(\Mux58~1_combout ),
	.datad(\Mux58~6_combout ),
	.cin(gnd),
	.combout(Mux58),
	.cout());
// synopsys translate_off
defparam \Mux58~9 .lut_mask = 16'hDDA0;
defparam \Mux58~9 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X65_Y30_N10
cycloneive_lcell_comb \Mux58~19 (
// Equation(s):
// Mux581 = (Selector8 & ((\Mux58~16_combout  & ((\Mux58~18_combout ))) # (!\Mux58~16_combout  & (\Mux58~11_combout )))) # (!Selector8 & (((\Mux58~16_combout ))))

	.dataa(\Mux58~11_combout ),
	.datab(Selector8),
	.datac(\Mux58~18_combout ),
	.datad(\Mux58~16_combout ),
	.cin(gnd),
	.combout(Mux581),
	.cout());
// synopsys translate_off
defparam \Mux58~19 .lut_mask = 16'hF388;
defparam \Mux58~19 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X63_Y32_N0
cycloneive_lcell_comb \Mux29~9 (
// Equation(s):
// Mux29 = (Selector5 & ((\Mux29~6_combout  & (\Mux29~8_combout )) # (!\Mux29~6_combout  & ((\Mux29~1_combout ))))) # (!Selector5 & (((\Mux29~6_combout ))))

	.dataa(\Mux29~8_combout ),
	.datab(Selector5),
	.datac(\Mux29~1_combout ),
	.datad(\Mux29~6_combout ),
	.cin(gnd),
	.combout(Mux29),
	.cout());
// synopsys translate_off
defparam \Mux29~9 .lut_mask = 16'hBBC0;
defparam \Mux29~9 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X63_Y32_N14
cycloneive_lcell_comb \Mux29~19 (
// Equation(s):
// Mux291 = (Selector3 & ((\Mux29~16_combout  & ((\Mux29~18_combout ))) # (!\Mux29~16_combout  & (\Mux29~11_combout )))) # (!Selector3 & (((\Mux29~16_combout ))))

	.dataa(\Mux29~11_combout ),
	.datab(Selector3),
	.datac(\Mux29~18_combout ),
	.datad(\Mux29~16_combout ),
	.cin(gnd),
	.combout(Mux291),
	.cout());
// synopsys translate_off
defparam \Mux29~19 .lut_mask = 16'hF388;
defparam \Mux29~19 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X65_Y31_N2
cycloneive_lcell_comb \Mux30~9 (
// Equation(s):
// Mux30 = (Selector5 & ((\Mux30~6_combout  & ((\Mux30~8_combout ))) # (!\Mux30~6_combout  & (\Mux30~1_combout )))) # (!Selector5 & (((\Mux30~6_combout ))))

	.dataa(\Mux30~1_combout ),
	.datab(Selector5),
	.datac(\Mux30~6_combout ),
	.datad(\Mux30~8_combout ),
	.cin(gnd),
	.combout(Mux30),
	.cout());
// synopsys translate_off
defparam \Mux30~9 .lut_mask = 16'hF838;
defparam \Mux30~9 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X65_Y31_N4
cycloneive_lcell_comb \Mux30~19 (
// Equation(s):
// Mux301 = (Selector2 & ((\Mux30~16_combout  & ((\Mux30~18_combout ))) # (!\Mux30~16_combout  & (\Mux30~11_combout )))) # (!Selector2 & (\Mux30~16_combout ))

	.dataa(Selector2),
	.datab(\Mux30~16_combout ),
	.datac(\Mux30~11_combout ),
	.datad(\Mux30~18_combout ),
	.cin(gnd),
	.combout(Mux301),
	.cout());
// synopsys translate_off
defparam \Mux30~19 .lut_mask = 16'hEC64;
defparam \Mux30~19 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y35_N12
cycloneive_lcell_comb \Mux63~9 (
// Equation(s):
// Mux63 = (Selector10 & ((\Mux63~6_combout  & ((\Mux63~8_combout ))) # (!\Mux63~6_combout  & (\Mux63~1_combout )))) # (!Selector10 & (((\Mux63~6_combout ))))

	.dataa(\Mux63~1_combout ),
	.datab(Selector10),
	.datac(\Mux63~8_combout ),
	.datad(\Mux63~6_combout ),
	.cin(gnd),
	.combout(Mux63),
	.cout());
// synopsys translate_off
defparam \Mux63~9 .lut_mask = 16'hF388;
defparam \Mux63~9 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y35_N8
cycloneive_lcell_comb \Mux63~19 (
// Equation(s):
// Mux631 = (Selector7 & ((\Mux63~16_combout  & ((\Mux63~18_combout ))) # (!\Mux63~16_combout  & (\Mux63~11_combout )))) # (!Selector7 & (((\Mux63~16_combout ))))

	.dataa(Selector7),
	.datab(\Mux63~11_combout ),
	.datac(\Mux63~16_combout ),
	.datad(\Mux63~18_combout ),
	.cin(gnd),
	.combout(Mux631),
	.cout());
// synopsys translate_off
defparam \Mux63~19 .lut_mask = 16'hF858;
defparam \Mux63~19 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X66_Y35_N8
cycloneive_lcell_comb \Mux62~9 (
// Equation(s):
// Mux62 = (\Mux62~6_combout  & (((\Mux62~8_combout )) # (!Selector10))) # (!\Mux62~6_combout  & (Selector10 & (\Mux62~1_combout )))

	.dataa(\Mux62~6_combout ),
	.datab(Selector10),
	.datac(\Mux62~1_combout ),
	.datad(\Mux62~8_combout ),
	.cin(gnd),
	.combout(Mux62),
	.cout());
// synopsys translate_off
defparam \Mux62~9 .lut_mask = 16'hEA62;
defparam \Mux62~9 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y35_N4
cycloneive_lcell_comb \Mux62~19 (
// Equation(s):
// Mux621 = (Selector8 & ((\Mux62~16_combout  & ((\Mux62~18_combout ))) # (!\Mux62~16_combout  & (\Mux62~11_combout )))) # (!Selector8 & (((\Mux62~16_combout ))))

	.dataa(\Mux62~11_combout ),
	.datab(\Mux62~18_combout ),
	.datac(Selector8),
	.datad(\Mux62~16_combout ),
	.cin(gnd),
	.combout(Mux621),
	.cout());
// synopsys translate_off
defparam \Mux62~19 .lut_mask = 16'hCFA0;
defparam \Mux62~19 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y34_N12
cycloneive_lcell_comb \Mux27~9 (
// Equation(s):
// Mux27 = (Selector5 & ((\Mux27~6_combout  & ((\Mux27~8_combout ))) # (!\Mux27~6_combout  & (\Mux27~1_combout )))) # (!Selector5 & (((\Mux27~6_combout ))))

	.dataa(Selector5),
	.datab(\Mux27~1_combout ),
	.datac(\Mux27~8_combout ),
	.datad(\Mux27~6_combout ),
	.cin(gnd),
	.combout(Mux27),
	.cout());
// synopsys translate_off
defparam \Mux27~9 .lut_mask = 16'hF588;
defparam \Mux27~9 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y34_N10
cycloneive_lcell_comb \Mux27~19 (
// Equation(s):
// Mux271 = (Selector3 & ((\Mux27~16_combout  & ((\Mux27~18_combout ))) # (!\Mux27~16_combout  & (\Mux27~11_combout )))) # (!Selector3 & (((\Mux27~16_combout ))))

	.dataa(\Mux27~11_combout ),
	.datab(\Mux27~18_combout ),
	.datac(Selector3),
	.datad(\Mux27~16_combout ),
	.cin(gnd),
	.combout(Mux271),
	.cout());
// synopsys translate_off
defparam \Mux27~19 .lut_mask = 16'hCFA0;
defparam \Mux27~19 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X70_Y37_N4
cycloneive_lcell_comb \Mux28~9 (
// Equation(s):
// Mux28 = (Selector5 & ((\Mux28~6_combout  & (\Mux28~8_combout )) # (!\Mux28~6_combout  & ((\Mux28~1_combout ))))) # (!Selector5 & (\Mux28~6_combout ))

	.dataa(Selector5),
	.datab(\Mux28~6_combout ),
	.datac(\Mux28~8_combout ),
	.datad(\Mux28~1_combout ),
	.cin(gnd),
	.combout(Mux28),
	.cout());
// synopsys translate_off
defparam \Mux28~9 .lut_mask = 16'hE6C4;
defparam \Mux28~9 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X70_Y37_N30
cycloneive_lcell_comb \Mux28~19 (
// Equation(s):
// Mux281 = (Selector2 & ((\Mux28~16_combout  & (\Mux28~18_combout )) # (!\Mux28~16_combout  & ((\Mux28~11_combout ))))) # (!Selector2 & (((\Mux28~16_combout ))))

	.dataa(Selector2),
	.datab(\Mux28~18_combout ),
	.datac(\Mux28~16_combout ),
	.datad(\Mux28~11_combout ),
	.cin(gnd),
	.combout(Mux281),
	.cout());
// synopsys translate_off
defparam \Mux28~19 .lut_mask = 16'hDAD0;
defparam \Mux28~19 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y35_N30
cycloneive_lcell_comb \Mux61~9 (
// Equation(s):
// Mux61 = (Selector10 & ((\Mux61~6_combout  & (\Mux61~8_combout )) # (!\Mux61~6_combout  & ((\Mux61~1_combout ))))) # (!Selector10 & (((\Mux61~6_combout ))))

	.dataa(Selector10),
	.datab(\Mux61~8_combout ),
	.datac(\Mux61~1_combout ),
	.datad(\Mux61~6_combout ),
	.cin(gnd),
	.combout(Mux61),
	.cout());
// synopsys translate_off
defparam \Mux61~9 .lut_mask = 16'hDDA0;
defparam \Mux61~9 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y35_N20
cycloneive_lcell_comb \Mux61~19 (
// Equation(s):
// Mux611 = (Selector7 & ((\Mux61~16_combout  & (\Mux61~18_combout )) # (!\Mux61~16_combout  & ((\Mux61~11_combout ))))) # (!Selector7 & (((\Mux61~16_combout ))))

	.dataa(Selector7),
	.datab(\Mux61~18_combout ),
	.datac(\Mux61~11_combout ),
	.datad(\Mux61~16_combout ),
	.cin(gnd),
	.combout(Mux611),
	.cout());
// synopsys translate_off
defparam \Mux61~19 .lut_mask = 16'hDDA0;
defparam \Mux61~19 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X68_Y36_N2
cycloneive_lcell_comb \Mux23~9 (
// Equation(s):
// Mux23 = (Selector5 & ((\Mux23~6_combout  & (\Mux23~8_combout )) # (!\Mux23~6_combout  & ((\Mux23~1_combout ))))) # (!Selector5 & (((\Mux23~6_combout ))))

	.dataa(\Mux23~8_combout ),
	.datab(Selector5),
	.datac(\Mux23~6_combout ),
	.datad(\Mux23~1_combout ),
	.cin(gnd),
	.combout(Mux23),
	.cout());
// synopsys translate_off
defparam \Mux23~9 .lut_mask = 16'hBCB0;
defparam \Mux23~9 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X68_Y36_N22
cycloneive_lcell_comb \Mux23~19 (
// Equation(s):
// Mux231 = (Selector3 & ((\Mux23~16_combout  & (\Mux23~18_combout )) # (!\Mux23~16_combout  & ((\Mux23~11_combout ))))) # (!Selector3 & (((\Mux23~16_combout ))))

	.dataa(\Mux23~18_combout ),
	.datab(Selector3),
	.datac(\Mux23~11_combout ),
	.datad(\Mux23~16_combout ),
	.cin(gnd),
	.combout(Mux231),
	.cout());
// synopsys translate_off
defparam \Mux23~19 .lut_mask = 16'hBBC0;
defparam \Mux23~19 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y40_N16
cycloneive_lcell_comb \Mux24~9 (
// Equation(s):
// Mux24 = (Selector5 & ((\Mux24~6_combout  & (\Mux24~8_combout )) # (!\Mux24~6_combout  & ((\Mux24~1_combout ))))) # (!Selector5 & (((\Mux24~6_combout ))))

	.dataa(Selector5),
	.datab(\Mux24~8_combout ),
	.datac(\Mux24~1_combout ),
	.datad(\Mux24~6_combout ),
	.cin(gnd),
	.combout(Mux24),
	.cout());
// synopsys translate_off
defparam \Mux24~9 .lut_mask = 16'hDDA0;
defparam \Mux24~9 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y40_N14
cycloneive_lcell_comb \Mux24~19 (
// Equation(s):
// Mux241 = (Selector2 & ((\Mux24~16_combout  & (\Mux24~18_combout )) # (!\Mux24~16_combout  & ((\Mux24~11_combout ))))) # (!Selector2 & (((\Mux24~16_combout ))))

	.dataa(\Mux24~18_combout ),
	.datab(\Mux24~11_combout ),
	.datac(Selector2),
	.datad(\Mux24~16_combout ),
	.cin(gnd),
	.combout(Mux241),
	.cout());
// synopsys translate_off
defparam \Mux24~19 .lut_mask = 16'hAFC0;
defparam \Mux24~19 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X67_Y36_N22
cycloneive_lcell_comb \Mux25~9 (
// Equation(s):
// Mux25 = (\Mux25~6_combout  & ((\Mux25~8_combout ) # ((!Selector5)))) # (!\Mux25~6_combout  & (((Selector5 & \Mux25~1_combout ))))

	.dataa(\Mux25~8_combout ),
	.datab(\Mux25~6_combout ),
	.datac(Selector5),
	.datad(\Mux25~1_combout ),
	.cin(gnd),
	.combout(Mux25),
	.cout());
// synopsys translate_off
defparam \Mux25~9 .lut_mask = 16'hBC8C;
defparam \Mux25~9 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X67_Y36_N0
cycloneive_lcell_comb \Mux25~19 (
// Equation(s):
// Mux251 = (Selector3 & ((\Mux25~16_combout  & (\Mux25~18_combout )) # (!\Mux25~16_combout  & ((\Mux25~11_combout ))))) # (!Selector3 & (((\Mux25~16_combout ))))

	.dataa(\Mux25~18_combout ),
	.datab(\Mux25~11_combout ),
	.datac(Selector3),
	.datad(\Mux25~16_combout ),
	.cin(gnd),
	.combout(Mux251),
	.cout());
// synopsys translate_off
defparam \Mux25~19 .lut_mask = 16'hAFC0;
defparam \Mux25~19 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X70_Y38_N0
cycloneive_lcell_comb \Mux26~9 (
// Equation(s):
// Mux26 = (Selector5 & ((\Mux26~6_combout  & (\Mux26~8_combout )) # (!\Mux26~6_combout  & ((\Mux26~1_combout ))))) # (!Selector5 & (((\Mux26~6_combout ))))

	.dataa(Selector5),
	.datab(\Mux26~8_combout ),
	.datac(\Mux26~6_combout ),
	.datad(\Mux26~1_combout ),
	.cin(gnd),
	.combout(Mux26),
	.cout());
// synopsys translate_off
defparam \Mux26~9 .lut_mask = 16'hDAD0;
defparam \Mux26~9 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X67_Y36_N28
cycloneive_lcell_comb \Mux26~19 (
// Equation(s):
// Mux261 = (\Mux26~16_combout  & (((\Mux26~18_combout )) # (!Selector2))) # (!\Mux26~16_combout  & (Selector2 & ((\Mux26~11_combout ))))

	.dataa(\Mux26~16_combout ),
	.datab(Selector2),
	.datac(\Mux26~18_combout ),
	.datad(\Mux26~11_combout ),
	.cin(gnd),
	.combout(Mux261),
	.cout());
// synopsys translate_off
defparam \Mux26~19 .lut_mask = 16'hE6A2;
defparam \Mux26~19 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y36_N20
cycloneive_lcell_comb \Mux60~9 (
// Equation(s):
// Mux60 = (Selector10 & ((\Mux60~6_combout  & (\Mux60~8_combout )) # (!\Mux60~6_combout  & ((\Mux60~1_combout ))))) # (!Selector10 & (((\Mux60~6_combout ))))

	.dataa(\Mux60~8_combout ),
	.datab(Selector10),
	.datac(\Mux60~1_combout ),
	.datad(\Mux60~6_combout ),
	.cin(gnd),
	.combout(Mux60),
	.cout());
// synopsys translate_off
defparam \Mux60~9 .lut_mask = 16'hBBC0;
defparam \Mux60~9 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y36_N12
cycloneive_lcell_comb \Mux60~19 (
// Equation(s):
// Mux601 = (Selector8 & ((\Mux60~16_combout  & ((\Mux60~18_combout ))) # (!\Mux60~16_combout  & (\Mux60~11_combout )))) # (!Selector8 & (((\Mux60~16_combout ))))

	.dataa(\Mux60~11_combout ),
	.datab(Selector8),
	.datac(\Mux60~18_combout ),
	.datad(\Mux60~16_combout ),
	.cin(gnd),
	.combout(Mux601),
	.cout());
// synopsys translate_off
defparam \Mux60~19 .lut_mask = 16'hF388;
defparam \Mux60~19 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X63_Y36_N14
cycloneive_lcell_comb \Mux15~9 (
// Equation(s):
// Mux15 = (\Mux15~6_combout  & (((\Mux15~8_combout )) # (!Selector5))) # (!\Mux15~6_combout  & (Selector5 & ((\Mux15~1_combout ))))

	.dataa(\Mux15~6_combout ),
	.datab(Selector5),
	.datac(\Mux15~8_combout ),
	.datad(\Mux15~1_combout ),
	.cin(gnd),
	.combout(Mux15),
	.cout());
// synopsys translate_off
defparam \Mux15~9 .lut_mask = 16'hE6A2;
defparam \Mux15~9 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X65_Y35_N0
cycloneive_lcell_comb \Mux15~19 (
// Equation(s):
// Mux151 = (Selector3 & ((\Mux15~16_combout  & ((\Mux15~18_combout ))) # (!\Mux15~16_combout  & (\Mux15~11_combout )))) # (!Selector3 & (((\Mux15~16_combout ))))

	.dataa(Selector3),
	.datab(\Mux15~11_combout ),
	.datac(\Mux15~18_combout ),
	.datad(\Mux15~16_combout ),
	.cin(gnd),
	.combout(Mux151),
	.cout());
// synopsys translate_off
defparam \Mux15~19 .lut_mask = 16'hF588;
defparam \Mux15~19 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y40_N14
cycloneive_lcell_comb \Mux16~9 (
// Equation(s):
// Mux16 = (Selector5 & ((\Mux16~6_combout  & ((\Mux16~8_combout ))) # (!\Mux16~6_combout  & (\Mux16~1_combout )))) # (!Selector5 & (((\Mux16~6_combout ))))

	.dataa(\Mux16~1_combout ),
	.datab(\Mux16~8_combout ),
	.datac(Selector5),
	.datad(\Mux16~6_combout ),
	.cin(gnd),
	.combout(Mux16),
	.cout());
// synopsys translate_off
defparam \Mux16~9 .lut_mask = 16'hCFA0;
defparam \Mux16~9 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y40_N6
cycloneive_lcell_comb \Mux16~19 (
// Equation(s):
// Mux161 = (Selector2 & ((\Mux16~16_combout  & (\Mux16~18_combout )) # (!\Mux16~16_combout  & ((\Mux16~11_combout ))))) # (!Selector2 & (((\Mux16~16_combout ))))

	.dataa(Selector2),
	.datab(\Mux16~18_combout ),
	.datac(\Mux16~11_combout ),
	.datad(\Mux16~16_combout ),
	.cin(gnd),
	.combout(Mux161),
	.cout());
// synopsys translate_off
defparam \Mux16~19 .lut_mask = 16'hDDA0;
defparam \Mux16~19 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X66_Y30_N4
cycloneive_lcell_comb \Mux17~9 (
// Equation(s):
// Mux17 = (\Mux17~6_combout  & (((\Mux17~8_combout )) # (!Selector5))) # (!\Mux17~6_combout  & (Selector5 & ((\Mux17~1_combout ))))

	.dataa(\Mux17~6_combout ),
	.datab(Selector5),
	.datac(\Mux17~8_combout ),
	.datad(\Mux17~1_combout ),
	.cin(gnd),
	.combout(Mux17),
	.cout());
// synopsys translate_off
defparam \Mux17~9 .lut_mask = 16'hE6A2;
defparam \Mux17~9 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X65_Y37_N0
cycloneive_lcell_comb \Mux17~19 (
// Equation(s):
// Mux171 = (Selector3 & ((\Mux17~16_combout  & (\Mux17~18_combout )) # (!\Mux17~16_combout  & ((\Mux17~11_combout ))))) # (!Selector3 & (((\Mux17~16_combout ))))

	.dataa(\Mux17~18_combout ),
	.datab(Selector3),
	.datac(\Mux17~16_combout ),
	.datad(\Mux17~11_combout ),
	.cin(gnd),
	.combout(Mux171),
	.cout());
// synopsys translate_off
defparam \Mux17~19 .lut_mask = 16'hBCB0;
defparam \Mux17~19 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X63_Y38_N16
cycloneive_lcell_comb \Mux18~9 (
// Equation(s):
// Mux18 = (\Mux18~6_combout  & ((\Mux18~8_combout ) # ((!Selector5)))) # (!\Mux18~6_combout  & (((\Mux18~1_combout  & Selector5))))

	.dataa(\Mux18~8_combout ),
	.datab(\Mux18~6_combout ),
	.datac(\Mux18~1_combout ),
	.datad(Selector5),
	.cin(gnd),
	.combout(Mux18),
	.cout());
// synopsys translate_off
defparam \Mux18~9 .lut_mask = 16'hB8CC;
defparam \Mux18~9 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X63_Y38_N12
cycloneive_lcell_comb \Mux18~19 (
// Equation(s):
// Mux181 = (Selector2 & ((\Mux18~16_combout  & ((\Mux18~18_combout ))) # (!\Mux18~16_combout  & (\Mux18~11_combout )))) # (!Selector2 & (((\Mux18~16_combout ))))

	.dataa(\Mux18~11_combout ),
	.datab(Selector2),
	.datac(\Mux18~18_combout ),
	.datad(\Mux18~16_combout ),
	.cin(gnd),
	.combout(Mux181),
	.cout());
// synopsys translate_off
defparam \Mux18~19 .lut_mask = 16'hF388;
defparam \Mux18~19 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y30_N12
cycloneive_lcell_comb \Mux19~9 (
// Equation(s):
// Mux19 = (Selector5 & ((\Mux19~6_combout  & ((\Mux19~8_combout ))) # (!\Mux19~6_combout  & (\Mux19~1_combout )))) # (!Selector5 & (((\Mux19~6_combout ))))

	.dataa(\Mux19~1_combout ),
	.datab(Selector5),
	.datac(\Mux19~8_combout ),
	.datad(\Mux19~6_combout ),
	.cin(gnd),
	.combout(Mux19),
	.cout());
// synopsys translate_off
defparam \Mux19~9 .lut_mask = 16'hF388;
defparam \Mux19~9 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X69_Y34_N14
cycloneive_lcell_comb \Mux19~19 (
// Equation(s):
// Mux191 = (Selector3 & ((\Mux19~16_combout  & (\Mux19~18_combout )) # (!\Mux19~16_combout  & ((\Mux19~11_combout ))))) # (!Selector3 & (((\Mux19~16_combout ))))

	.dataa(\Mux19~18_combout ),
	.datab(\Mux19~11_combout ),
	.datac(Selector3),
	.datad(\Mux19~16_combout ),
	.cin(gnd),
	.combout(Mux191),
	.cout());
// synopsys translate_off
defparam \Mux19~19 .lut_mask = 16'hAFC0;
defparam \Mux19~19 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X63_Y38_N2
cycloneive_lcell_comb \Mux20~9 (
// Equation(s):
// Mux20 = (Selector5 & ((\Mux20~6_combout  & (\Mux20~8_combout )) # (!\Mux20~6_combout  & ((\Mux20~1_combout ))))) # (!Selector5 & (((\Mux20~6_combout ))))

	.dataa(Selector5),
	.datab(\Mux20~8_combout ),
	.datac(\Mux20~1_combout ),
	.datad(\Mux20~6_combout ),
	.cin(gnd),
	.combout(Mux20),
	.cout());
// synopsys translate_off
defparam \Mux20~9 .lut_mask = 16'hDDA0;
defparam \Mux20~9 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X63_Y38_N6
cycloneive_lcell_comb \Mux20~19 (
// Equation(s):
// Mux201 = (\Mux20~16_combout  & ((\Mux20~18_combout ) # ((!Selector2)))) # (!\Mux20~16_combout  & (((Selector2 & \Mux20~11_combout ))))

	.dataa(\Mux20~18_combout ),
	.datab(\Mux20~16_combout ),
	.datac(Selector2),
	.datad(\Mux20~11_combout ),
	.cin(gnd),
	.combout(Mux201),
	.cout());
// synopsys translate_off
defparam \Mux20~19 .lut_mask = 16'hBC8C;
defparam \Mux20~19 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X66_Y36_N8
cycloneive_lcell_comb \Mux21~9 (
// Equation(s):
// Mux21 = (\Mux21~6_combout  & (((\Mux21~8_combout ) # (!Selector5)))) # (!\Mux21~6_combout  & (\Mux21~1_combout  & (Selector5)))

	.dataa(\Mux21~1_combout ),
	.datab(\Mux21~6_combout ),
	.datac(Selector5),
	.datad(\Mux21~8_combout ),
	.cin(gnd),
	.combout(Mux21),
	.cout());
// synopsys translate_off
defparam \Mux21~9 .lut_mask = 16'hEC2C;
defparam \Mux21~9 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X66_Y36_N2
cycloneive_lcell_comb \Mux21~19 (
// Equation(s):
// Mux211 = (Selector3 & ((\Mux21~16_combout  & ((\Mux21~18_combout ))) # (!\Mux21~16_combout  & (\Mux21~11_combout )))) # (!Selector3 & (((\Mux21~16_combout ))))

	.dataa(Selector3),
	.datab(\Mux21~11_combout ),
	.datac(\Mux21~18_combout ),
	.datad(\Mux21~16_combout ),
	.cin(gnd),
	.combout(Mux211),
	.cout());
// synopsys translate_off
defparam \Mux21~19 .lut_mask = 16'hF588;
defparam \Mux21~19 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y41_N24
cycloneive_lcell_comb \Mux22~9 (
// Equation(s):
// Mux22 = (Selector5 & ((\Mux22~6_combout  & (\Mux22~8_combout )) # (!\Mux22~6_combout  & ((\Mux22~1_combout ))))) # (!Selector5 & (((\Mux22~6_combout ))))

	.dataa(\Mux22~8_combout ),
	.datab(Selector5),
	.datac(\Mux22~1_combout ),
	.datad(\Mux22~6_combout ),
	.cin(gnd),
	.combout(Mux22),
	.cout());
// synopsys translate_off
defparam \Mux22~9 .lut_mask = 16'hBBC0;
defparam \Mux22~9 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y41_N14
cycloneive_lcell_comb \Mux22~19 (
// Equation(s):
// Mux221 = (Selector2 & ((\Mux22~16_combout  & (\Mux22~18_combout )) # (!\Mux22~16_combout  & ((\Mux22~11_combout ))))) # (!Selector2 & (((\Mux22~16_combout ))))

	.dataa(Selector2),
	.datab(\Mux22~18_combout ),
	.datac(\Mux22~11_combout ),
	.datad(\Mux22~16_combout ),
	.cin(gnd),
	.combout(Mux221),
	.cout());
// synopsys translate_off
defparam \Mux22~19 .lut_mask = 16'hDDA0;
defparam \Mux22~19 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y41_N24
cycloneive_lcell_comb \Mux59~9 (
// Equation(s):
// Mux59 = (Selector10 & ((\Mux59~6_combout  & ((\Mux59~8_combout ))) # (!\Mux59~6_combout  & (\Mux59~1_combout )))) # (!Selector10 & (((\Mux59~6_combout ))))

	.dataa(Selector10),
	.datab(\Mux59~1_combout ),
	.datac(\Mux59~8_combout ),
	.datad(\Mux59~6_combout ),
	.cin(gnd),
	.combout(Mux59),
	.cout());
// synopsys translate_off
defparam \Mux59~9 .lut_mask = 16'hF588;
defparam \Mux59~9 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y41_N4
cycloneive_lcell_comb \Mux59~19 (
// Equation(s):
// Mux591 = (\Mux59~16_combout  & (((\Mux59~18_combout )) # (!Selector7))) # (!\Mux59~16_combout  & (Selector7 & ((\Mux59~11_combout ))))

	.dataa(\Mux59~16_combout ),
	.datab(Selector7),
	.datac(\Mux59~18_combout ),
	.datad(\Mux59~11_combout ),
	.cin(gnd),
	.combout(Mux591),
	.cout());
// synopsys translate_off
defparam \Mux59~19 .lut_mask = 16'hE6A2;
defparam \Mux59~19 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y33_N0
cycloneive_lcell_comb \Mux0~9 (
// Equation(s):
// Mux0 = (Selector5 & ((\Mux0~6_combout  & (\Mux0~8_combout )) # (!\Mux0~6_combout  & ((\Mux0~1_combout ))))) # (!Selector5 & (((\Mux0~6_combout ))))

	.dataa(\Mux0~8_combout ),
	.datab(Selector5),
	.datac(\Mux0~1_combout ),
	.datad(\Mux0~6_combout ),
	.cin(gnd),
	.combout(Mux0),
	.cout());
// synopsys translate_off
defparam \Mux0~9 .lut_mask = 16'hBBC0;
defparam \Mux0~9 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y33_N4
cycloneive_lcell_comb \Mux0~19 (
// Equation(s):
// Mux01 = (\Mux0~16_combout  & (((\Mux0~18_combout )) # (!Selector2))) # (!\Mux0~16_combout  & (Selector2 & (\Mux0~11_combout )))

	.dataa(\Mux0~16_combout ),
	.datab(Selector2),
	.datac(\Mux0~11_combout ),
	.datad(\Mux0~18_combout ),
	.cin(gnd),
	.combout(Mux01),
	.cout());
// synopsys translate_off
defparam \Mux0~19 .lut_mask = 16'hEA62;
defparam \Mux0~19 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y33_N28
cycloneive_lcell_comb \Mux2~9 (
// Equation(s):
// Mux2 = (Selector5 & ((\Mux2~6_combout  & ((\Mux2~8_combout ))) # (!\Mux2~6_combout  & (\Mux2~1_combout )))) # (!Selector5 & (((\Mux2~6_combout ))))

	.dataa(\Mux2~1_combout ),
	.datab(Selector5),
	.datac(\Mux2~6_combout ),
	.datad(\Mux2~8_combout ),
	.cin(gnd),
	.combout(Mux2),
	.cout());
// synopsys translate_off
defparam \Mux2~9 .lut_mask = 16'hF838;
defparam \Mux2~9 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y33_N18
cycloneive_lcell_comb \Mux2~19 (
// Equation(s):
// Mux210 = (Selector2 & ((\Mux2~16_combout  & (\Mux2~18_combout )) # (!\Mux2~16_combout  & ((\Mux2~11_combout ))))) # (!Selector2 & (((\Mux2~16_combout ))))

	.dataa(\Mux2~18_combout ),
	.datab(Selector2),
	.datac(\Mux2~11_combout ),
	.datad(\Mux2~16_combout ),
	.cin(gnd),
	.combout(Mux210),
	.cout());
// synopsys translate_off
defparam \Mux2~19 .lut_mask = 16'hBBC0;
defparam \Mux2~19 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X65_Y35_N10
cycloneive_lcell_comb \Mux1~9 (
// Equation(s):
// Mux1 = (Selector5 & ((\Mux1~6_combout  & ((\Mux1~8_combout ))) # (!\Mux1~6_combout  & (\Mux1~1_combout )))) # (!Selector5 & (\Mux1~6_combout ))

	.dataa(Selector5),
	.datab(\Mux1~6_combout ),
	.datac(\Mux1~1_combout ),
	.datad(\Mux1~8_combout ),
	.cin(gnd),
	.combout(Mux1),
	.cout());
// synopsys translate_off
defparam \Mux1~9 .lut_mask = 16'hEC64;
defparam \Mux1~9 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X65_Y37_N24
cycloneive_lcell_comb \Mux1~19 (
// Equation(s):
// Mux11 = (Selector3 & ((\Mux1~16_combout  & ((\Mux1~18_combout ))) # (!\Mux1~16_combout  & (\Mux1~11_combout )))) # (!Selector3 & (((\Mux1~16_combout ))))

	.dataa(Selector3),
	.datab(\Mux1~11_combout ),
	.datac(\Mux1~18_combout ),
	.datad(\Mux1~16_combout ),
	.cin(gnd),
	.combout(Mux11),
	.cout());
// synopsys translate_off
defparam \Mux1~19 .lut_mask = 16'hF588;
defparam \Mux1~19 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X63_Y39_N18
cycloneive_lcell_comb \Mux3~9 (
// Equation(s):
// Mux3 = (Selector5 & ((\Mux3~6_combout  & ((\Mux3~8_combout ))) # (!\Mux3~6_combout  & (\Mux3~1_combout )))) # (!Selector5 & (((\Mux3~6_combout ))))

	.dataa(\Mux3~1_combout ),
	.datab(Selector5),
	.datac(\Mux3~8_combout ),
	.datad(\Mux3~6_combout ),
	.cin(gnd),
	.combout(Mux3),
	.cout());
// synopsys translate_off
defparam \Mux3~9 .lut_mask = 16'hF388;
defparam \Mux3~9 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X63_Y39_N8
cycloneive_lcell_comb \Mux3~19 (
// Equation(s):
// Mux31 = (\Mux3~16_combout  & (((\Mux3~18_combout )) # (!Selector3))) # (!\Mux3~16_combout  & (Selector3 & ((\Mux3~11_combout ))))

	.dataa(\Mux3~16_combout ),
	.datab(Selector3),
	.datac(\Mux3~18_combout ),
	.datad(\Mux3~11_combout ),
	.cin(gnd),
	.combout(Mux31),
	.cout());
// synopsys translate_off
defparam \Mux3~19 .lut_mask = 16'hE6A2;
defparam \Mux3~19 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X63_Y39_N14
cycloneive_lcell_comb \Mux4~9 (
// Equation(s):
// Mux4 = (Selector5 & ((\Mux4~6_combout  & (\Mux4~8_combout )) # (!\Mux4~6_combout  & ((\Mux4~1_combout ))))) # (!Selector5 & (((\Mux4~6_combout ))))

	.dataa(\Mux4~8_combout ),
	.datab(Selector5),
	.datac(\Mux4~1_combout ),
	.datad(\Mux4~6_combout ),
	.cin(gnd),
	.combout(Mux4),
	.cout());
// synopsys translate_off
defparam \Mux4~9 .lut_mask = 16'hBBC0;
defparam \Mux4~9 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X63_Y39_N2
cycloneive_lcell_comb \Mux4~19 (
// Equation(s):
// Mux410 = (Selector2 & ((\Mux4~16_combout  & ((\Mux4~18_combout ))) # (!\Mux4~16_combout  & (\Mux4~11_combout )))) # (!Selector2 & (\Mux4~16_combout ))

	.dataa(Selector2),
	.datab(\Mux4~16_combout ),
	.datac(\Mux4~11_combout ),
	.datad(\Mux4~18_combout ),
	.cin(gnd),
	.combout(Mux410),
	.cout());
// synopsys translate_off
defparam \Mux4~19 .lut_mask = 16'hEC64;
defparam \Mux4~19 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X63_Y32_N18
cycloneive_lcell_comb \Mux5~9 (
// Equation(s):
// Mux5 = (Selector5 & ((\Mux5~6_combout  & (\Mux5~8_combout )) # (!\Mux5~6_combout  & ((\Mux5~1_combout ))))) # (!Selector5 & (((\Mux5~6_combout ))))

	.dataa(\Mux5~8_combout ),
	.datab(Selector5),
	.datac(\Mux5~1_combout ),
	.datad(\Mux5~6_combout ),
	.cin(gnd),
	.combout(Mux5),
	.cout());
// synopsys translate_off
defparam \Mux5~9 .lut_mask = 16'hBBC0;
defparam \Mux5~9 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X63_Y32_N26
cycloneive_lcell_comb \Mux5~19 (
// Equation(s):
// Mux510 = (Selector3 & ((\Mux5~16_combout  & (\Mux5~18_combout )) # (!\Mux5~16_combout  & ((\Mux5~11_combout ))))) # (!Selector3 & (((\Mux5~16_combout ))))

	.dataa(\Mux5~18_combout ),
	.datab(Selector3),
	.datac(\Mux5~11_combout ),
	.datad(\Mux5~16_combout ),
	.cin(gnd),
	.combout(Mux510),
	.cout());
// synopsys translate_off
defparam \Mux5~19 .lut_mask = 16'hBBC0;
defparam \Mux5~19 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X65_Y31_N12
cycloneive_lcell_comb \Mux6~9 (
// Equation(s):
// Mux6 = (Selector5 & ((\Mux6~6_combout  & ((\Mux6~8_combout ))) # (!\Mux6~6_combout  & (\Mux6~1_combout )))) # (!Selector5 & (((\Mux6~6_combout ))))

	.dataa(\Mux6~1_combout ),
	.datab(Selector5),
	.datac(\Mux6~8_combout ),
	.datad(\Mux6~6_combout ),
	.cin(gnd),
	.combout(Mux6),
	.cout());
// synopsys translate_off
defparam \Mux6~9 .lut_mask = 16'hF388;
defparam \Mux6~9 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X65_Y31_N22
cycloneive_lcell_comb \Mux6~19 (
// Equation(s):
// Mux64 = (\Mux6~16_combout  & (((\Mux6~18_combout ) # (!Selector2)))) # (!\Mux6~16_combout  & (\Mux6~11_combout  & (Selector2)))

	.dataa(\Mux6~11_combout ),
	.datab(\Mux6~16_combout ),
	.datac(Selector2),
	.datad(\Mux6~18_combout ),
	.cin(gnd),
	.combout(Mux64),
	.cout());
// synopsys translate_off
defparam \Mux6~19 .lut_mask = 16'hEC2C;
defparam \Mux6~19 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y34_N2
cycloneive_lcell_comb \Mux7~9 (
// Equation(s):
// Mux7 = (Selector5 & ((\Mux7~6_combout  & (\Mux7~8_combout )) # (!\Mux7~6_combout  & ((\Mux7~1_combout ))))) # (!Selector5 & (((\Mux7~6_combout ))))

	.dataa(Selector5),
	.datab(\Mux7~8_combout ),
	.datac(\Mux7~6_combout ),
	.datad(\Mux7~1_combout ),
	.cin(gnd),
	.combout(Mux7),
	.cout());
// synopsys translate_off
defparam \Mux7~9 .lut_mask = 16'hDAD0;
defparam \Mux7~9 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y34_N14
cycloneive_lcell_comb \Mux7~19 (
// Equation(s):
// Mux71 = (Selector3 & ((\Mux7~16_combout  & ((\Mux7~18_combout ))) # (!\Mux7~16_combout  & (\Mux7~11_combout )))) # (!Selector3 & (((\Mux7~16_combout ))))

	.dataa(\Mux7~11_combout ),
	.datab(Selector3),
	.datac(\Mux7~18_combout ),
	.datad(\Mux7~16_combout ),
	.cin(gnd),
	.combout(Mux71),
	.cout());
// synopsys translate_off
defparam \Mux7~19 .lut_mask = 16'hF388;
defparam \Mux7~19 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X70_Y37_N26
cycloneive_lcell_comb \Mux8~9 (
// Equation(s):
// Mux8 = (Selector5 & ((\Mux8~6_combout  & (\Mux8~8_combout )) # (!\Mux8~6_combout  & ((\Mux8~1_combout ))))) # (!Selector5 & (((\Mux8~6_combout ))))

	.dataa(\Mux8~8_combout ),
	.datab(\Mux8~1_combout ),
	.datac(Selector5),
	.datad(\Mux8~6_combout ),
	.cin(gnd),
	.combout(Mux8),
	.cout());
// synopsys translate_off
defparam \Mux8~9 .lut_mask = 16'hAFC0;
defparam \Mux8~9 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X70_Y37_N8
cycloneive_lcell_comb \Mux8~19 (
// Equation(s):
// Mux81 = (Selector2 & ((\Mux8~16_combout  & (\Mux8~18_combout )) # (!\Mux8~16_combout  & ((\Mux8~11_combout ))))) # (!Selector2 & (((\Mux8~16_combout ))))

	.dataa(Selector2),
	.datab(\Mux8~18_combout ),
	.datac(\Mux8~11_combout ),
	.datad(\Mux8~16_combout ),
	.cin(gnd),
	.combout(Mux81),
	.cout());
// synopsys translate_off
defparam \Mux8~19 .lut_mask = 16'hDDA0;
defparam \Mux8~19 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X68_Y36_N16
cycloneive_lcell_comb \Mux9~9 (
// Equation(s):
// Mux9 = (\Mux9~6_combout  & (((\Mux9~8_combout )) # (!Selector5))) # (!\Mux9~6_combout  & (Selector5 & ((\Mux9~1_combout ))))

	.dataa(\Mux9~6_combout ),
	.datab(Selector5),
	.datac(\Mux9~8_combout ),
	.datad(\Mux9~1_combout ),
	.cin(gnd),
	.combout(Mux9),
	.cout());
// synopsys translate_off
defparam \Mux9~9 .lut_mask = 16'hE6A2;
defparam \Mux9~9 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X68_Y36_N30
cycloneive_lcell_comb \Mux9~19 (
// Equation(s):
// Mux91 = (Selector3 & ((\Mux9~16_combout  & ((\Mux9~18_combout ))) # (!\Mux9~16_combout  & (\Mux9~11_combout )))) # (!Selector3 & (((\Mux9~16_combout ))))

	.dataa(\Mux9~11_combout ),
	.datab(Selector3),
	.datac(\Mux9~18_combout ),
	.datad(\Mux9~16_combout ),
	.cin(gnd),
	.combout(Mux91),
	.cout());
// synopsys translate_off
defparam \Mux9~19 .lut_mask = 16'hF388;
defparam \Mux9~19 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y38_N8
cycloneive_lcell_comb \Mux10~9 (
// Equation(s):
// Mux10 = (Selector5 & ((\Mux10~6_combout  & (\Mux10~8_combout )) # (!\Mux10~6_combout  & ((\Mux10~1_combout ))))) # (!Selector5 & (((\Mux10~6_combout ))))

	.dataa(\Mux10~8_combout ),
	.datab(Selector5),
	.datac(\Mux10~1_combout ),
	.datad(\Mux10~6_combout ),
	.cin(gnd),
	.combout(Mux10),
	.cout());
// synopsys translate_off
defparam \Mux10~9 .lut_mask = 16'hBBC0;
defparam \Mux10~9 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y38_N10
cycloneive_lcell_comb \Mux10~19 (
// Equation(s):
// Mux101 = (Selector2 & ((\Mux10~16_combout  & (\Mux10~18_combout )) # (!\Mux10~16_combout  & ((\Mux10~11_combout ))))) # (!Selector2 & (((\Mux10~16_combout ))))

	.dataa(Selector2),
	.datab(\Mux10~18_combout ),
	.datac(\Mux10~11_combout ),
	.datad(\Mux10~16_combout ),
	.cin(gnd),
	.combout(Mux101),
	.cout());
// synopsys translate_off
defparam \Mux10~19 .lut_mask = 16'hDDA0;
defparam \Mux10~19 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y40_N2
cycloneive_lcell_comb \Mux11~9 (
// Equation(s):
// Mux111 = (Selector5 & ((\Mux11~6_combout  & (\Mux11~8_combout )) # (!\Mux11~6_combout  & ((\Mux11~1_combout ))))) # (!Selector5 & (((\Mux11~6_combout ))))

	.dataa(Selector5),
	.datab(\Mux11~8_combout ),
	.datac(\Mux11~1_combout ),
	.datad(\Mux11~6_combout ),
	.cin(gnd),
	.combout(Mux111),
	.cout());
// synopsys translate_off
defparam \Mux11~9 .lut_mask = 16'hDDA0;
defparam \Mux11~9 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y40_N22
cycloneive_lcell_comb \Mux11~19 (
// Equation(s):
// Mux112 = (Selector3 & ((\Mux11~16_combout  & (\Mux11~18_combout )) # (!\Mux11~16_combout  & ((\Mux11~11_combout ))))) # (!Selector3 & (\Mux11~16_combout ))

	.dataa(Selector3),
	.datab(\Mux11~16_combout ),
	.datac(\Mux11~18_combout ),
	.datad(\Mux11~11_combout ),
	.cin(gnd),
	.combout(Mux112),
	.cout());
// synopsys translate_off
defparam \Mux11~19 .lut_mask = 16'hE6C4;
defparam \Mux11~19 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X67_Y36_N2
cycloneive_lcell_comb \Mux12~9 (
// Equation(s):
// Mux12 = (Selector5 & ((\Mux12~6_combout  & ((\Mux12~8_combout ))) # (!\Mux12~6_combout  & (\Mux12~1_combout )))) # (!Selector5 & (((\Mux12~6_combout ))))

	.dataa(\Mux12~1_combout ),
	.datab(\Mux12~8_combout ),
	.datac(Selector5),
	.datad(\Mux12~6_combout ),
	.cin(gnd),
	.combout(Mux12),
	.cout());
// synopsys translate_off
defparam \Mux12~9 .lut_mask = 16'hCFA0;
defparam \Mux12~9 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X67_Y36_N14
cycloneive_lcell_comb \Mux12~19 (
// Equation(s):
// Mux121 = (Selector2 & ((\Mux12~16_combout  & (\Mux12~18_combout )) # (!\Mux12~16_combout  & ((\Mux12~11_combout ))))) # (!Selector2 & (((\Mux12~16_combout ))))

	.dataa(\Mux12~18_combout ),
	.datab(Selector2),
	.datac(\Mux12~16_combout ),
	.datad(\Mux12~11_combout ),
	.cin(gnd),
	.combout(Mux121),
	.cout());
// synopsys translate_off
defparam \Mux12~19 .lut_mask = 16'hBCB0;
defparam \Mux12~19 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X63_Y36_N24
cycloneive_lcell_comb \Mux13~9 (
// Equation(s):
// Mux13 = (Selector5 & ((\Mux13~6_combout  & (\Mux13~8_combout )) # (!\Mux13~6_combout  & ((\Mux13~1_combout ))))) # (!Selector5 & (((\Mux13~6_combout ))))

	.dataa(\Mux13~8_combout ),
	.datab(Selector5),
	.datac(\Mux13~1_combout ),
	.datad(\Mux13~6_combout ),
	.cin(gnd),
	.combout(Mux13),
	.cout());
// synopsys translate_off
defparam \Mux13~9 .lut_mask = 16'hBBC0;
defparam \Mux13~9 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X63_Y36_N16
cycloneive_lcell_comb \Mux13~19 (
// Equation(s):
// Mux131 = (Selector3 & ((\Mux13~16_combout  & ((\Mux13~18_combout ))) # (!\Mux13~16_combout  & (\Mux13~11_combout )))) # (!Selector3 & (\Mux13~16_combout ))

	.dataa(Selector3),
	.datab(\Mux13~16_combout ),
	.datac(\Mux13~11_combout ),
	.datad(\Mux13~18_combout ),
	.cin(gnd),
	.combout(Mux131),
	.cout());
// synopsys translate_off
defparam \Mux13~19 .lut_mask = 16'hEC64;
defparam \Mux13~19 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y40_N0
cycloneive_lcell_comb \Mux14~9 (
// Equation(s):
// Mux14 = (Selector5 & ((\Mux14~6_combout  & (\Mux14~8_combout )) # (!\Mux14~6_combout  & ((\Mux14~1_combout ))))) # (!Selector5 & (((\Mux14~6_combout ))))

	.dataa(Selector5),
	.datab(\Mux14~8_combout ),
	.datac(\Mux14~1_combout ),
	.datad(\Mux14~6_combout ),
	.cin(gnd),
	.combout(Mux14),
	.cout());
// synopsys translate_off
defparam \Mux14~9 .lut_mask = 16'hDDA0;
defparam \Mux14~9 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y40_N8
cycloneive_lcell_comb \Mux14~19 (
// Equation(s):
// Mux141 = (Selector2 & ((\Mux14~16_combout  & (\Mux14~18_combout )) # (!\Mux14~16_combout  & ((\Mux14~11_combout ))))) # (!Selector2 & (((\Mux14~16_combout ))))

	.dataa(Selector2),
	.datab(\Mux14~18_combout ),
	.datac(\Mux14~11_combout ),
	.datad(\Mux14~16_combout ),
	.cin(gnd),
	.combout(Mux141),
	.cout());
// synopsys translate_off
defparam \Mux14~19 .lut_mask = 16'hDDA0;
defparam \Mux14~19 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y40_N8
cycloneive_lcell_comb \Mux31~9 (
// Equation(s):
// Mux311 = (Selector5 & ((\Mux31~6_combout  & (\Mux31~8_combout )) # (!\Mux31~6_combout  & ((\Mux31~1_combout ))))) # (!Selector5 & (((\Mux31~6_combout ))))

	.dataa(Selector5),
	.datab(\Mux31~8_combout ),
	.datac(\Mux31~1_combout ),
	.datad(\Mux31~6_combout ),
	.cin(gnd),
	.combout(Mux311),
	.cout());
// synopsys translate_off
defparam \Mux31~9 .lut_mask = 16'hDDA0;
defparam \Mux31~9 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y40_N30
cycloneive_lcell_comb \Mux31~19 (
// Equation(s):
// Mux312 = (Selector3 & ((\Mux31~16_combout  & ((\Mux31~18_combout ))) # (!\Mux31~16_combout  & (\Mux31~11_combout )))) # (!Selector3 & (\Mux31~16_combout ))

	.dataa(Selector3),
	.datab(\Mux31~16_combout ),
	.datac(\Mux31~11_combout ),
	.datad(\Mux31~18_combout ),
	.cin(gnd),
	.combout(Mux312),
	.cout());
// synopsys translate_off
defparam \Mux31~19 .lut_mask = 16'hEC64;
defparam \Mux31~19 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y35_N12
cycloneive_lcell_comb \register~64 (
// Equation(s):
// \register~64_combout  = (WideOr01 & ((\wdat[31]~0_combout ) # ((plif_memwbrtnaddr_l_31 & plif_memwbregsrc_l_1))))

	.dataa(plif_memwbrtnaddr_l_31),
	.datab(WideOr0),
	.datac(wdat_31),
	.datad(plif_memwbregsrc_l_1),
	.cin(gnd),
	.combout(\register~64_combout ),
	.cout());
// synopsys translate_off
defparam \register~64 .lut_mask = 16'hC8C0;
defparam \register~64 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X66_Y37_N30
cycloneive_lcell_comb \Decoder0~32 (
// Equation(s):
// \Decoder0~32_combout  = (plif_memwbwsel_l_4 & (plif_memwbwsel_l_1 & (plif_memwbregen_l & !plif_memwbwsel_l_3)))

	.dataa(plif_memwbwsel_l_4),
	.datab(plif_memwbwsel_l_1),
	.datac(plif_memwbregen_l),
	.datad(plif_memwbwsel_l_3),
	.cin(gnd),
	.combout(\Decoder0~32_combout ),
	.cout());
// synopsys translate_off
defparam \Decoder0~32 .lut_mask = 16'h0080;
defparam \Decoder0~32 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y37_N10
cycloneive_lcell_comb \Decoder0~37 (
// Equation(s):
// \Decoder0~37_combout  = (plif_memwbwsel_l_0 & (plif_memwbwsel_l_2 & \Decoder0~32_combout ))

	.dataa(gnd),
	.datab(plif_memwbwsel_l_0),
	.datac(plif_memwbwsel_l_2),
	.datad(\Decoder0~32_combout ),
	.cin(gnd),
	.combout(\Decoder0~37_combout ),
	.cout());
// synopsys translate_off
defparam \Decoder0~37 .lut_mask = 16'hC000;
defparam \Decoder0~37 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X60_Y35_N9
dffeas \register[23][31] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\register~64_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~37_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\register[23][31]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \register[23][31] .is_wysiwyg = "true";
defparam \register[23][31] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X62_Y37_N30
cycloneive_lcell_comb \Decoder0~40 (
// Equation(s):
// \Decoder0~40_combout  = (\Decoder0~29_combout  & (plif_memwbwsel_l_0 & (plif_memwbwsel_l_2 & plif_memwbwsel_l_4)))

	.dataa(\Decoder0~29_combout ),
	.datab(plif_memwbwsel_l_0),
	.datac(plif_memwbwsel_l_2),
	.datad(plif_memwbwsel_l_4),
	.cin(gnd),
	.combout(\Decoder0~40_combout ),
	.cout());
// synopsys translate_off
defparam \Decoder0~40 .lut_mask = 16'h8000;
defparam \Decoder0~40 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X61_Y33_N15
dffeas \register[31][31] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\register~64_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~40_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\register[31][31]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \register[31][31] .is_wysiwyg = "true";
defparam \register[31][31] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X62_Y39_N4
cycloneive_lcell_comb \register[27][31]~feeder (
// Equation(s):
// \register[27][31]~feeder_combout  = \register~64_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(\register~64_combout ),
	.cin(gnd),
	.combout(\register[27][31]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \register[27][31]~feeder .lut_mask = 16'hFF00;
defparam \register[27][31]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y37_N6
cycloneive_lcell_comb \Decoder0~29 (
// Equation(s):
// \Decoder0~29_combout  = (plif_memwbwsel_l_3 & (plif_memwbwsel_l_1 & plif_memwbregen_l))

	.dataa(plif_memwbwsel_l_3),
	.datab(gnd),
	.datac(plif_memwbwsel_l_1),
	.datad(plif_memwbregen_l),
	.cin(gnd),
	.combout(\Decoder0~29_combout ),
	.cout());
// synopsys translate_off
defparam \Decoder0~29 .lut_mask = 16'hA000;
defparam \Decoder0~29 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y37_N0
cycloneive_lcell_comb \Decoder0~38 (
// Equation(s):
// \Decoder0~38_combout  = (!plif_memwbwsel_l_2 & (plif_memwbwsel_l_4 & (plif_memwbwsel_l_0 & \Decoder0~29_combout )))

	.dataa(plif_memwbwsel_l_2),
	.datab(plif_memwbwsel_l_4),
	.datac(plif_memwbwsel_l_0),
	.datad(\Decoder0~29_combout ),
	.cin(gnd),
	.combout(\Decoder0~38_combout ),
	.cout());
// synopsys translate_off
defparam \Decoder0~38 .lut_mask = 16'h4000;
defparam \Decoder0~38 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X62_Y39_N5
dffeas \register[27][31] (
	.clk(!CLK),
	.d(\register[27][31]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~38_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\register[27][31]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \register[27][31] .is_wysiwyg = "true";
defparam \register[27][31] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X66_Y37_N12
cycloneive_lcell_comb \Decoder0~39 (
// Equation(s):
// \Decoder0~39_combout  = (plif_memwbwsel_l_0 & (\Decoder0~32_combout  & !plif_memwbwsel_l_2))

	.dataa(gnd),
	.datab(plif_memwbwsel_l_0),
	.datac(\Decoder0~32_combout ),
	.datad(plif_memwbwsel_l_2),
	.cin(gnd),
	.combout(\Decoder0~39_combout ),
	.cout());
// synopsys translate_off
defparam \Decoder0~39 .lut_mask = 16'h00C0;
defparam \Decoder0~39 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X60_Y35_N11
dffeas \register[19][31] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\register~64_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~39_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\register[19][31]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \register[19][31] .is_wysiwyg = "true";
defparam \register[19][31] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X60_Y35_N10
cycloneive_lcell_comb \Mux32~7 (
// Equation(s):
// \Mux32~7_combout  = (Selector8 & (((Selector7)))) # (!Selector8 & ((Selector7 & (\register[27][31]~q )) # (!Selector7 & ((\register[19][31]~q )))))

	.dataa(Selector8),
	.datab(\register[27][31]~q ),
	.datac(\register[19][31]~q ),
	.datad(Selector7),
	.cin(gnd),
	.combout(\Mux32~7_combout ),
	.cout());
// synopsys translate_off
defparam \Mux32~7 .lut_mask = 16'hEE50;
defparam \Mux32~7 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X67_Y35_N30
cycloneive_lcell_comb \Mux32~8 (
// Equation(s):
// \Mux32~8_combout  = (\Mux32~7_combout  & (((\register[31][31]~q ) # (!Selector8)))) # (!\Mux32~7_combout  & (\register[23][31]~q  & ((Selector8))))

	.dataa(\register[23][31]~q ),
	.datab(\register[31][31]~q ),
	.datac(\Mux32~7_combout ),
	.datad(Selector8),
	.cin(gnd),
	.combout(\Mux32~8_combout ),
	.cout());
// synopsys translate_off
defparam \Mux32~8 .lut_mask = 16'hCAF0;
defparam \Mux32~8 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y38_N12
cycloneive_lcell_comb \register[29][31]~feeder (
// Equation(s):
// \register[29][31]~feeder_combout  = \register~64_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(\register~64_combout ),
	.cin(gnd),
	.combout(\register[29][31]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \register[29][31]~feeder .lut_mask = 16'hFF00;
defparam \register[29][31]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X66_Y37_N16
cycloneive_lcell_comb \Decoder0~27 (
// Equation(s):
// \Decoder0~27_combout  = (plif_memwbwsel_l_4 & (!plif_memwbwsel_l_1 & (plif_memwbregen_l & plif_memwbwsel_l_3)))

	.dataa(plif_memwbwsel_l_4),
	.datab(plif_memwbwsel_l_1),
	.datac(plif_memwbregen_l),
	.datad(plif_memwbwsel_l_3),
	.cin(gnd),
	.combout(\Decoder0~27_combout ),
	.cout());
// synopsys translate_off
defparam \Decoder0~27 .lut_mask = 16'h2000;
defparam \Decoder0~27 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X65_Y34_N6
cycloneive_lcell_comb \Decoder0~28 (
// Equation(s):
// \Decoder0~28_combout  = (plif_memwbwsel_l_2 & (plif_memwbwsel_l_0 & \Decoder0~27_combout ))

	.dataa(plif_memwbwsel_l_2),
	.datab(gnd),
	.datac(plif_memwbwsel_l_0),
	.datad(\Decoder0~27_combout ),
	.cin(gnd),
	.combout(\Decoder0~28_combout ),
	.cout());
// synopsys translate_off
defparam \Decoder0~28 .lut_mask = 16'hA000;
defparam \Decoder0~28 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X61_Y38_N13
dffeas \register[29][31] (
	.clk(!CLK),
	.d(\register[29][31]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~28_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\register[29][31]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \register[29][31] .is_wysiwyg = "true";
defparam \register[29][31] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X66_Y37_N20
cycloneive_lcell_comb \Decoder0~21 (
// Equation(s):
// \Decoder0~21_combout  = (!plif_memwbwsel_l_1 & (plif_memwbregen_l & plif_memwbwsel_l_2))

	.dataa(gnd),
	.datab(plif_memwbwsel_l_1),
	.datac(plif_memwbregen_l),
	.datad(plif_memwbwsel_l_2),
	.cin(gnd),
	.combout(\Decoder0~21_combout ),
	.cout());
// synopsys translate_off
defparam \Decoder0~21 .lut_mask = 16'h3000;
defparam \Decoder0~21 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X66_Y37_N14
cycloneive_lcell_comb \Decoder0~22 (
// Equation(s):
// \Decoder0~22_combout  = (plif_memwbwsel_l_4 & (plif_memwbwsel_l_0 & (!plif_memwbwsel_l_3 & \Decoder0~21_combout )))

	.dataa(plif_memwbwsel_l_4),
	.datab(plif_memwbwsel_l_0),
	.datac(plif_memwbwsel_l_3),
	.datad(\Decoder0~21_combout ),
	.cin(gnd),
	.combout(\Decoder0~22_combout ),
	.cout());
// synopsys translate_off
defparam \Decoder0~22 .lut_mask = 16'h0800;
defparam \Decoder0~22 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X61_Y35_N13
dffeas \register[21][31] (
	.clk(!CLK),
	.d(\register~64_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~22_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\register[21][31]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \register[21][31] .is_wysiwyg = "true";
defparam \register[21][31] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X61_Y37_N28
cycloneive_lcell_comb \register[25][31]~feeder (
// Equation(s):
// \register[25][31]~feeder_combout  = \register~64_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(\register~64_combout ),
	.datad(gnd),
	.cin(gnd),
	.combout(\register[25][31]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \register[25][31]~feeder .lut_mask = 16'hF0F0;
defparam \register[25][31]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y37_N8
cycloneive_lcell_comb \Decoder0~23 (
// Equation(s):
// \Decoder0~23_combout  = (plif_memwbwsel_l_3 & plif_memwbregen_l)

	.dataa(gnd),
	.datab(plif_memwbwsel_l_3),
	.datac(plif_memwbregen_l),
	.datad(gnd),
	.cin(gnd),
	.combout(\Decoder0~23_combout ),
	.cout());
// synopsys translate_off
defparam \Decoder0~23 .lut_mask = 16'hC0C0;
defparam \Decoder0~23 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y37_N6
cycloneive_lcell_comb \Decoder0~24 (
// Equation(s):
// \Decoder0~24_combout  = (plif_memwbwsel_l_0 & (Decoder0 & (plif_memwbwsel_l_4 & \Decoder0~23_combout )))

	.dataa(plif_memwbwsel_l_0),
	.datab(Decoder0),
	.datac(plif_memwbwsel_l_4),
	.datad(\Decoder0~23_combout ),
	.cin(gnd),
	.combout(\Decoder0~24_combout ),
	.cout());
// synopsys translate_off
defparam \Decoder0~24 .lut_mask = 16'h8000;
defparam \Decoder0~24 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X61_Y37_N29
dffeas \register[25][31] (
	.clk(!CLK),
	.d(\register[25][31]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~24_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\register[25][31]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \register[25][31] .is_wysiwyg = "true";
defparam \register[25][31] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X61_Y37_N30
cycloneive_lcell_comb \Mux32~0 (
// Equation(s):
// \Mux32~0_combout  = (Selector8 & (((Selector7)))) # (!Selector8 & ((Selector7 & ((\register[25][31]~q ))) # (!Selector7 & (\register[17][31]~q ))))

	.dataa(\register[17][31]~q ),
	.datab(\register[25][31]~q ),
	.datac(Selector8),
	.datad(Selector7),
	.cin(gnd),
	.combout(\Mux32~0_combout ),
	.cout());
// synopsys translate_off
defparam \Mux32~0 .lut_mask = 16'hFC0A;
defparam \Mux32~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y37_N0
cycloneive_lcell_comb \Mux32~1 (
// Equation(s):
// \Mux32~1_combout  = (Selector8 & ((\Mux32~0_combout  & (\register[29][31]~q )) # (!\Mux32~0_combout  & ((\register[21][31]~q ))))) # (!Selector8 & (((\Mux32~0_combout ))))

	.dataa(\register[29][31]~q ),
	.datab(\register[21][31]~q ),
	.datac(Selector8),
	.datad(\Mux32~0_combout ),
	.cin(gnd),
	.combout(\Mux32~1_combout ),
	.cout());
// synopsys translate_off
defparam \Mux32~1 .lut_mask = 16'hAFC0;
defparam \Mux32~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y37_N0
cycloneive_lcell_comb \Decoder0~34 (
// Equation(s):
// \Decoder0~34_combout  = (!plif_memwbwsel_l_0 & (Decoder0 & (plif_memwbwsel_l_4 & \Decoder0~23_combout )))

	.dataa(plif_memwbwsel_l_0),
	.datab(Decoder0),
	.datac(plif_memwbwsel_l_4),
	.datad(\Decoder0~23_combout ),
	.cin(gnd),
	.combout(\Decoder0~34_combout ),
	.cout());
// synopsys translate_off
defparam \Decoder0~34 .lut_mask = 16'h4000;
defparam \Decoder0~34 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X65_Y35_N17
dffeas \register[24][31] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\register~64_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~34_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\register[24][31]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \register[24][31] .is_wysiwyg = "true";
defparam \register[24][31] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X58_Y37_N10
cycloneive_lcell_comb \Decoder0~25 (
// Equation(s):
// \Decoder0~25_combout  = (plif_memwbregen_l & (plif_memwbwsel_l_4 & (!plif_memwbwsel_l_3 & Decoder0)))

	.dataa(plif_memwbregen_l),
	.datab(plif_memwbwsel_l_4),
	.datac(plif_memwbwsel_l_3),
	.datad(Decoder0),
	.cin(gnd),
	.combout(\Decoder0~25_combout ),
	.cout());
// synopsys translate_off
defparam \Decoder0~25 .lut_mask = 16'h0800;
defparam \Decoder0~25 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y37_N30
cycloneive_lcell_comb \Decoder0~36 (
// Equation(s):
// \Decoder0~36_combout  = (!plif_memwbwsel_l_0 & \Decoder0~25_combout )

	.dataa(plif_memwbwsel_l_0),
	.datab(gnd),
	.datac(gnd),
	.datad(\Decoder0~25_combout ),
	.cin(gnd),
	.combout(\Decoder0~36_combout ),
	.cout());
// synopsys translate_off
defparam \Decoder0~36 .lut_mask = 16'h5500;
defparam \Decoder0~36 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X65_Y35_N27
dffeas \register[16][31] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\register~64_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~36_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\register[16][31]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \register[16][31] .is_wysiwyg = "true";
defparam \register[16][31] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X65_Y35_N26
cycloneive_lcell_comb \Mux32~4 (
// Equation(s):
// \Mux32~4_combout  = (Selector8 & ((\register[20][31]~q ) # ((Selector7)))) # (!Selector8 & (((\register[16][31]~q  & !Selector7))))

	.dataa(\register[20][31]~q ),
	.datab(Selector8),
	.datac(\register[16][31]~q ),
	.datad(Selector7),
	.cin(gnd),
	.combout(\Mux32~4_combout ),
	.cout());
// synopsys translate_off
defparam \Mux32~4 .lut_mask = 16'hCCB8;
defparam \Mux32~4 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X66_Y35_N12
cycloneive_lcell_comb \register[28][31]~feeder (
// Equation(s):
// \register[28][31]~feeder_combout  = \register~64_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(\register~64_combout ),
	.cin(gnd),
	.combout(\register[28][31]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \register[28][31]~feeder .lut_mask = 16'hFF00;
defparam \register[28][31]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X66_Y37_N28
cycloneive_lcell_comb \Decoder0~57 (
// Equation(s):
// \Decoder0~57_combout  = (\Decoder0~27_combout  & (!plif_memwbwsel_l_0 & plif_memwbwsel_l_2))

	.dataa(\Decoder0~27_combout ),
	.datab(plif_memwbwsel_l_0),
	.datac(gnd),
	.datad(plif_memwbwsel_l_2),
	.cin(gnd),
	.combout(\Decoder0~57_combout ),
	.cout());
// synopsys translate_off
defparam \Decoder0~57 .lut_mask = 16'h2200;
defparam \Decoder0~57 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X66_Y35_N13
dffeas \register[28][31] (
	.clk(!CLK),
	.d(\register[28][31]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~57_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\register[28][31]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \register[28][31] .is_wysiwyg = "true";
defparam \register[28][31] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X66_Y35_N26
cycloneive_lcell_comb \Mux32~5 (
// Equation(s):
// \Mux32~5_combout  = (Selector7 & ((\Mux32~4_combout  & ((\register[28][31]~q ))) # (!\Mux32~4_combout  & (\register[24][31]~q )))) # (!Selector7 & (((\Mux32~4_combout ))))

	.dataa(Selector7),
	.datab(\register[24][31]~q ),
	.datac(\Mux32~4_combout ),
	.datad(\register[28][31]~q ),
	.cin(gnd),
	.combout(\Mux32~5_combout ),
	.cout());
// synopsys translate_off
defparam \Mux32~5 .lut_mask = 16'hF858;
defparam \Mux32~5 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X68_Y35_N12
cycloneive_lcell_comb \register[26][31]~feeder (
// Equation(s):
// \register[26][31]~feeder_combout  = \register~64_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(\register~64_combout ),
	.cin(gnd),
	.combout(\register[26][31]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \register[26][31]~feeder .lut_mask = 16'hFF00;
defparam \register[26][31]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y37_N28
cycloneive_lcell_comb \Decoder0~30 (
// Equation(s):
// \Decoder0~30_combout  = (!plif_memwbwsel_l_0 & (!plif_memwbwsel_l_2 & plif_memwbwsel_l_4))

	.dataa(gnd),
	.datab(plif_memwbwsel_l_0),
	.datac(plif_memwbwsel_l_2),
	.datad(plif_memwbwsel_l_4),
	.cin(gnd),
	.combout(\Decoder0~30_combout ),
	.cout());
// synopsys translate_off
defparam \Decoder0~30 .lut_mask = 16'h0300;
defparam \Decoder0~30 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X66_Y37_N24
cycloneive_lcell_comb \Decoder0~54 (
// Equation(s):
// \Decoder0~54_combout  = (plif_memwbregen_l & (plif_memwbwsel_l_3 & (plif_memwbwsel_l_1 & \Decoder0~30_combout )))

	.dataa(plif_memwbregen_l),
	.datab(plif_memwbwsel_l_3),
	.datac(plif_memwbwsel_l_1),
	.datad(\Decoder0~30_combout ),
	.cin(gnd),
	.combout(\Decoder0~54_combout ),
	.cout());
// synopsys translate_off
defparam \Decoder0~54 .lut_mask = 16'h8000;
defparam \Decoder0~54 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X68_Y35_N13
dffeas \register[26][31] (
	.clk(!CLK),
	.d(\register[26][31]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~54_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\register[26][31]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \register[26][31] .is_wysiwyg = "true";
defparam \register[26][31] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X62_Y37_N24
cycloneive_lcell_comb \Decoder0~33 (
// Equation(s):
// \Decoder0~33_combout  = (!plif_memwbwsel_l_3 & (\Decoder0~30_combout  & (plif_memwbwsel_l_1 & plif_memwbregen_l)))

	.dataa(plif_memwbwsel_l_3),
	.datab(\Decoder0~30_combout ),
	.datac(plif_memwbwsel_l_1),
	.datad(plif_memwbregen_l),
	.cin(gnd),
	.combout(\Decoder0~33_combout ),
	.cout());
// synopsys translate_off
defparam \Decoder0~33 .lut_mask = 16'h4000;
defparam \Decoder0~33 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X69_Y35_N19
dffeas \register[18][31] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\register~64_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~33_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\register[18][31]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \register[18][31] .is_wysiwyg = "true";
defparam \register[18][31] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X67_Y37_N4
cycloneive_lcell_comb \Decoder0~55 (
// Equation(s):
// \Decoder0~55_combout  = (!plif_memwbwsel_l_0 & (plif_memwbwsel_l_2 & \Decoder0~32_combout ))

	.dataa(plif_memwbwsel_l_0),
	.datab(plif_memwbwsel_l_2),
	.datac(gnd),
	.datad(\Decoder0~32_combout ),
	.cin(gnd),
	.combout(\Decoder0~55_combout ),
	.cout());
// synopsys translate_off
defparam \Decoder0~55 .lut_mask = 16'h4400;
defparam \Decoder0~55 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X69_Y35_N21
dffeas \register[22][31] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\register~64_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~55_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\register[22][31]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \register[22][31] .is_wysiwyg = "true";
defparam \register[22][31] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X69_Y35_N20
cycloneive_lcell_comb \Mux32~2 (
// Equation(s):
// \Mux32~2_combout  = (Selector8 & (((\register[22][31]~q ) # (Selector7)))) # (!Selector8 & (\register[18][31]~q  & ((!Selector7))))

	.dataa(Selector8),
	.datab(\register[18][31]~q ),
	.datac(\register[22][31]~q ),
	.datad(Selector7),
	.cin(gnd),
	.combout(\Mux32~2_combout ),
	.cout());
// synopsys translate_off
defparam \Mux32~2 .lut_mask = 16'hAAE4;
defparam \Mux32~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X68_Y35_N2
cycloneive_lcell_comb \register[30][31]~feeder (
// Equation(s):
// \register[30][31]~feeder_combout  = \register~64_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(\register~64_combout ),
	.cin(gnd),
	.combout(\register[30][31]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \register[30][31]~feeder .lut_mask = 16'hFF00;
defparam \register[30][31]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y37_N12
cycloneive_lcell_comb \Decoder0~56 (
// Equation(s):
// \Decoder0~56_combout  = (\Decoder0~29_combout  & (plif_memwbwsel_l_4 & (plif_memwbwsel_l_2 & !plif_memwbwsel_l_0)))

	.dataa(\Decoder0~29_combout ),
	.datab(plif_memwbwsel_l_4),
	.datac(plif_memwbwsel_l_2),
	.datad(plif_memwbwsel_l_0),
	.cin(gnd),
	.combout(\Decoder0~56_combout ),
	.cout());
// synopsys translate_off
defparam \Decoder0~56 .lut_mask = 16'h0080;
defparam \Decoder0~56 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X68_Y35_N3
dffeas \register[30][31] (
	.clk(!CLK),
	.d(\register[30][31]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~56_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\register[30][31]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \register[30][31] .is_wysiwyg = "true";
defparam \register[30][31] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X68_Y35_N28
cycloneive_lcell_comb \Mux32~3 (
// Equation(s):
// \Mux32~3_combout  = (Selector7 & ((\Mux32~2_combout  & ((\register[30][31]~q ))) # (!\Mux32~2_combout  & (\register[26][31]~q )))) # (!Selector7 & (((\Mux32~2_combout ))))

	.dataa(Selector7),
	.datab(\register[26][31]~q ),
	.datac(\Mux32~2_combout ),
	.datad(\register[30][31]~q ),
	.cin(gnd),
	.combout(\Mux32~3_combout ),
	.cout());
// synopsys translate_off
defparam \Mux32~3 .lut_mask = 16'hF858;
defparam \Mux32~3 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X67_Y35_N16
cycloneive_lcell_comb \Mux32~6 (
// Equation(s):
// \Mux32~6_combout  = (Selector10 & (Selector91)) # (!Selector10 & ((Selector91 & ((\Mux32~3_combout ))) # (!Selector91 & (\Mux32~5_combout ))))

	.dataa(Selector10),
	.datab(Selector91),
	.datac(\Mux32~5_combout ),
	.datad(\Mux32~3_combout ),
	.cin(gnd),
	.combout(\Mux32~6_combout ),
	.cout());
// synopsys translate_off
defparam \Mux32~6 .lut_mask = 16'hDC98;
defparam \Mux32~6 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y37_N16
cycloneive_lcell_comb \Decoder0~41 (
// Equation(s):
// \Decoder0~41_combout  = (!plif_memwbwsel_l_3 & (!plif_memwbwsel_l_4 & (plif_memwbwsel_l_1 & plif_memwbregen_l)))

	.dataa(plif_memwbwsel_l_3),
	.datab(plif_memwbwsel_l_4),
	.datac(plif_memwbwsel_l_1),
	.datad(plif_memwbregen_l),
	.cin(gnd),
	.combout(\Decoder0~41_combout ),
	.cout());
// synopsys translate_off
defparam \Decoder0~41 .lut_mask = 16'h1000;
defparam \Decoder0~41 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X66_Y34_N22
cycloneive_lcell_comb \Decoder0~43 (
// Equation(s):
// \Decoder0~43_combout  = (plif_memwbwsel_l_2 & (plif_memwbwsel_l_0 & \Decoder0~41_combout ))

	.dataa(plif_memwbwsel_l_2),
	.datab(plif_memwbwsel_l_0),
	.datac(gnd),
	.datad(\Decoder0~41_combout ),
	.cin(gnd),
	.combout(\Decoder0~43_combout ),
	.cout());
// synopsys translate_off
defparam \Decoder0~43 .lut_mask = 16'h8800;
defparam \Decoder0~43 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X68_Y31_N27
dffeas \register[7][31] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\register~64_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~43_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\register[7][31]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \register[7][31] .is_wysiwyg = "true";
defparam \register[7][31] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X66_Y37_N2
cycloneive_lcell_comb \Decoder0~58 (
// Equation(s):
// \Decoder0~58_combout  = (\Decoder0~41_combout  & (!plif_memwbwsel_l_0 & plif_memwbwsel_l_2))

	.dataa(\Decoder0~41_combout ),
	.datab(plif_memwbwsel_l_0),
	.datac(gnd),
	.datad(plif_memwbwsel_l_2),
	.cin(gnd),
	.combout(\Decoder0~58_combout ),
	.cout());
// synopsys translate_off
defparam \Decoder0~58 .lut_mask = 16'h2200;
defparam \Decoder0~58 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X68_Y31_N9
dffeas \register[6][31] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\register~64_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~58_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\register[6][31]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \register[6][31] .is_wysiwyg = "true";
defparam \register[6][31] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X66_Y37_N8
cycloneive_lcell_comb \Decoder0~59 (
// Equation(s):
// \Decoder0~59_combout  = (!plif_memwbwsel_l_4 & (plif_memwbwsel_l_0 & (!plif_memwbwsel_l_3 & \Decoder0~21_combout )))

	.dataa(plif_memwbwsel_l_4),
	.datab(plif_memwbwsel_l_0),
	.datac(plif_memwbwsel_l_3),
	.datad(\Decoder0~21_combout ),
	.cin(gnd),
	.combout(\Decoder0~59_combout ),
	.cout());
// synopsys translate_off
defparam \Decoder0~59 .lut_mask = 16'h0400;
defparam \Decoder0~59 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X69_Y31_N25
dffeas \register[5][31] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\register~64_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~59_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\register[5][31]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \register[5][31] .is_wysiwyg = "true";
defparam \register[5][31] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X69_Y31_N24
cycloneive_lcell_comb \Mux32~10 (
// Equation(s):
// \Mux32~10_combout  = (Selector91 & (((Selector10)))) # (!Selector91 & ((Selector10 & ((\register[5][31]~q ))) # (!Selector10 & (\register[4][31]~q ))))

	.dataa(\register[4][31]~q ),
	.datab(Selector91),
	.datac(\register[5][31]~q ),
	.datad(Selector10),
	.cin(gnd),
	.combout(\Mux32~10_combout ),
	.cout());
// synopsys translate_off
defparam \Mux32~10 .lut_mask = 16'hFC22;
defparam \Mux32~10 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X68_Y31_N8
cycloneive_lcell_comb \Mux32~11 (
// Equation(s):
// \Mux32~11_combout  = (Selector91 & ((\Mux32~10_combout  & (\register[7][31]~q )) # (!\Mux32~10_combout  & ((\register[6][31]~q ))))) # (!Selector91 & (((\Mux32~10_combout ))))

	.dataa(\register[7][31]~q ),
	.datab(Selector91),
	.datac(\register[6][31]~q ),
	.datad(\Mux32~10_combout ),
	.cin(gnd),
	.combout(\Mux32~11_combout ),
	.cout());
// synopsys translate_off
defparam \Mux32~11 .lut_mask = 16'hBBC0;
defparam \Mux32~11 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y32_N24
cycloneive_lcell_comb \register[14][31]~feeder (
// Equation(s):
// \register[14][31]~feeder_combout  = \register~64_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(\register~64_combout ),
	.datad(gnd),
	.cin(gnd),
	.combout(\register[14][31]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \register[14][31]~feeder .lut_mask = 16'hF0F0;
defparam \register[14][31]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y37_N26
cycloneive_lcell_comb \Decoder0~61 (
// Equation(s):
// \Decoder0~61_combout  = (\Decoder0~29_combout  & (!plif_memwbwsel_l_4 & (plif_memwbwsel_l_2 & !plif_memwbwsel_l_0)))

	.dataa(\Decoder0~29_combout ),
	.datab(plif_memwbwsel_l_4),
	.datac(plif_memwbwsel_l_2),
	.datad(plif_memwbwsel_l_0),
	.cin(gnd),
	.combout(\Decoder0~61_combout ),
	.cout());
// synopsys translate_off
defparam \Decoder0~61 .lut_mask = 16'h0020;
defparam \Decoder0~61 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X62_Y32_N25
dffeas \register[14][31] (
	.clk(!CLK),
	.d(\register[14][31]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~61_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\register[14][31]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \register[14][31] .is_wysiwyg = "true";
defparam \register[14][31] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X59_Y37_N4
cycloneive_lcell_comb \Decoder0~51 (
// Equation(s):
// \Decoder0~51_combout  = (plif_memwbwsel_l_0 & (!plif_memwbwsel_l_1 & (!plif_memwbwsel_l_4 & plif_memwbwsel_l_2)))

	.dataa(plif_memwbwsel_l_0),
	.datab(plif_memwbwsel_l_1),
	.datac(plif_memwbwsel_l_4),
	.datad(plif_memwbwsel_l_2),
	.cin(gnd),
	.combout(\Decoder0~51_combout ),
	.cout());
// synopsys translate_off
defparam \Decoder0~51 .lut_mask = 16'h0200;
defparam \Decoder0~51 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y37_N2
cycloneive_lcell_comb \Decoder0~62 (
// Equation(s):
// \Decoder0~62_combout  = (plif_memwbwsel_l_3 & (\Decoder0~51_combout  & plif_memwbregen_l))

	.dataa(plif_memwbwsel_l_3),
	.datab(gnd),
	.datac(\Decoder0~51_combout ),
	.datad(plif_memwbregen_l),
	.cin(gnd),
	.combout(\Decoder0~62_combout ),
	.cout());
// synopsys translate_off
defparam \Decoder0~62 .lut_mask = 16'hA000;
defparam \Decoder0~62 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X62_Y30_N1
dffeas \register[13][31] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\register~64_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~62_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\register[13][31]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \register[13][31] .is_wysiwyg = "true";
defparam \register[13][31] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X62_Y30_N0
cycloneive_lcell_comb \Mux32~17 (
// Equation(s):
// \Mux32~17_combout  = (Selector91 & (((Selector10)))) # (!Selector91 & ((Selector10 & ((\register[13][31]~q ))) # (!Selector10 & (\register[12][31]~q ))))

	.dataa(\register[12][31]~q ),
	.datab(Selector91),
	.datac(\register[13][31]~q ),
	.datad(Selector10),
	.cin(gnd),
	.combout(\Mux32~17_combout ),
	.cout());
// synopsys translate_off
defparam \Mux32~17 .lut_mask = 16'hFC22;
defparam \Mux32~17 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y35_N2
cycloneive_lcell_comb \register[15][31]~feeder (
// Equation(s):
// \register[15][31]~feeder_combout  = \register~64_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(\register~64_combout ),
	.cin(gnd),
	.combout(\register[15][31]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \register[15][31]~feeder .lut_mask = 16'hFF00;
defparam \register[15][31]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y37_N14
cycloneive_lcell_comb \Decoder0~53 (
// Equation(s):
// \Decoder0~53_combout  = (plif_memwbwsel_l_2 & (plif_memwbwsel_l_0 & (!plif_memwbwsel_l_4 & \Decoder0~29_combout )))

	.dataa(plif_memwbwsel_l_2),
	.datab(plif_memwbwsel_l_0),
	.datac(plif_memwbwsel_l_4),
	.datad(\Decoder0~29_combout ),
	.cin(gnd),
	.combout(\Decoder0~53_combout ),
	.cout());
// synopsys translate_off
defparam \Decoder0~53 .lut_mask = 16'h0800;
defparam \Decoder0~53 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X61_Y35_N3
dffeas \register[15][31] (
	.clk(!CLK),
	.d(\register[15][31]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~53_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\register[15][31]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \register[15][31] .is_wysiwyg = "true";
defparam \register[15][31] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X61_Y35_N20
cycloneive_lcell_comb \Mux32~18 (
// Equation(s):
// \Mux32~18_combout  = (\Mux32~17_combout  & (((\register[15][31]~q ) # (!Selector91)))) # (!\Mux32~17_combout  & (\register[14][31]~q  & (Selector91)))

	.dataa(\register[14][31]~q ),
	.datab(\Mux32~17_combout ),
	.datac(Selector91),
	.datad(\register[15][31]~q ),
	.cin(gnd),
	.combout(\Mux32~18_combout ),
	.cout());
// synopsys translate_off
defparam \Mux32~18 .lut_mask = 16'hEC2C;
defparam \Mux32~18 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X66_Y37_N10
cycloneive_lcell_comb \Decoder0~50 (
// Equation(s):
// \Decoder0~50_combout  = (!plif_memwbwsel_l_0 & (\Decoder0~41_combout  & !plif_memwbwsel_l_2))

	.dataa(gnd),
	.datab(plif_memwbwsel_l_0),
	.datac(\Decoder0~41_combout ),
	.datad(plif_memwbwsel_l_2),
	.cin(gnd),
	.combout(\Decoder0~50_combout ),
	.cout());
// synopsys translate_off
defparam \Decoder0~50 .lut_mask = 16'h0030;
defparam \Decoder0~50 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X67_Y34_N5
dffeas \register[2][31] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\register~64_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~50_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\register[2][31]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \register[2][31] .is_wysiwyg = "true";
defparam \register[2][31] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X66_Y37_N4
cycloneive_lcell_comb \Decoder0~48 (
// Equation(s):
// \Decoder0~48_combout  = (plif_memwbwsel_l_0 & (\Decoder0~41_combout  & !plif_memwbwsel_l_2))

	.dataa(gnd),
	.datab(plif_memwbwsel_l_0),
	.datac(\Decoder0~41_combout ),
	.datad(plif_memwbwsel_l_2),
	.cin(gnd),
	.combout(\Decoder0~48_combout ),
	.cout());
// synopsys translate_off
defparam \Decoder0~48 .lut_mask = 16'h00C0;
defparam \Decoder0~48 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X65_Y33_N9
dffeas \register[3][31] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\register~64_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~48_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\register[3][31]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \register[3][31] .is_wysiwyg = "true";
defparam \register[3][31] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X59_Y37_N0
cycloneive_lcell_comb \Decoder0~42 (
// Equation(s):
// \Decoder0~42_combout  = (!plif_memwbwsel_l_4 & !plif_memwbwsel_l_3)

	.dataa(plif_memwbwsel_l_4),
	.datab(gnd),
	.datac(plif_memwbwsel_l_3),
	.datad(gnd),
	.cin(gnd),
	.combout(\Decoder0~42_combout ),
	.cout());
// synopsys translate_off
defparam \Decoder0~42 .lut_mask = 16'h0505;
defparam \Decoder0~42 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y37_N30
cycloneive_lcell_comb \Decoder0~49 (
// Equation(s):
// \Decoder0~49_combout  = (plif_memwbwsel_l_0 & (\Decoder0~42_combout  & (plif_memwbregen_l & Decoder0)))

	.dataa(plif_memwbwsel_l_0),
	.datab(\Decoder0~42_combout ),
	.datac(plif_memwbregen_l),
	.datad(Decoder0),
	.cin(gnd),
	.combout(\Decoder0~49_combout ),
	.cout());
// synopsys translate_off
defparam \Decoder0~49 .lut_mask = 16'h8000;
defparam \Decoder0~49 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X65_Y33_N7
dffeas \register[1][31] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\register~64_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~49_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\register[1][31]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \register[1][31] .is_wysiwyg = "true";
defparam \register[1][31] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X65_Y33_N6
cycloneive_lcell_comb \Mux32~14 (
// Equation(s):
// \Mux32~14_combout  = (Selector10 & ((Selector91 & (\register[3][31]~q )) # (!Selector91 & ((\register[1][31]~q )))))

	.dataa(Selector91),
	.datab(\register[3][31]~q ),
	.datac(\register[1][31]~q ),
	.datad(Selector10),
	.cin(gnd),
	.combout(\Mux32~14_combout ),
	.cout());
// synopsys translate_off
defparam \Mux32~14 .lut_mask = 16'hD800;
defparam \Mux32~14 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X67_Y34_N14
cycloneive_lcell_comb \Mux32~15 (
// Equation(s):
// \Mux32~15_combout  = (\Mux32~14_combout ) # ((!Selector10 & (\register[2][31]~q  & Selector91)))

	.dataa(Selector10),
	.datab(\register[2][31]~q ),
	.datac(\Mux32~14_combout ),
	.datad(Selector91),
	.cin(gnd),
	.combout(\Mux32~15_combout ),
	.cout());
// synopsys translate_off
defparam \Mux32~15 .lut_mask = 16'hF4F0;
defparam \Mux32~15 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y37_N24
cycloneive_lcell_comb \Decoder0~44 (
// Equation(s):
// \Decoder0~44_combout  = (plif_memwbwsel_l_0 & (Decoder0 & (!plif_memwbwsel_l_4 & \Decoder0~23_combout )))

	.dataa(plif_memwbwsel_l_0),
	.datab(Decoder0),
	.datac(plif_memwbwsel_l_4),
	.datad(\Decoder0~23_combout ),
	.cin(gnd),
	.combout(\Decoder0~44_combout ),
	.cout());
// synopsys translate_off
defparam \Decoder0~44 .lut_mask = 16'h0800;
defparam \Decoder0~44 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X66_Y38_N29
dffeas \register[9][31] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\register~64_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~44_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\register[9][31]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \register[9][31] .is_wysiwyg = "true";
defparam \register[9][31] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X61_Y37_N14
cycloneive_lcell_comb \Decoder0~46 (
// Equation(s):
// \Decoder0~46_combout  = (!plif_memwbwsel_l_0 & (Decoder0 & (!plif_memwbwsel_l_4 & \Decoder0~23_combout )))

	.dataa(plif_memwbwsel_l_0),
	.datab(Decoder0),
	.datac(plif_memwbwsel_l_4),
	.datad(\Decoder0~23_combout ),
	.cin(gnd),
	.combout(\Decoder0~46_combout ),
	.cout());
// synopsys translate_off
defparam \Decoder0~46 .lut_mask = 16'h0400;
defparam \Decoder0~46 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X62_Y41_N27
dffeas \register[8][31] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\register~64_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~46_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\register[8][31]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \register[8][31] .is_wysiwyg = "true";
defparam \register[8][31] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X66_Y37_N6
cycloneive_lcell_comb \Decoder0~45 (
// Equation(s):
// \Decoder0~45_combout  = (!plif_memwbwsel_l_4 & (!plif_memwbwsel_l_0 & (\Decoder0~29_combout  & !plif_memwbwsel_l_2)))

	.dataa(plif_memwbwsel_l_4),
	.datab(plif_memwbwsel_l_0),
	.datac(\Decoder0~29_combout ),
	.datad(plif_memwbwsel_l_2),
	.cin(gnd),
	.combout(\Decoder0~45_combout ),
	.cout());
// synopsys translate_off
defparam \Decoder0~45 .lut_mask = 16'h0010;
defparam \Decoder0~45 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X62_Y41_N17
dffeas \register[10][31] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\register~64_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~45_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\register[10][31]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \register[10][31] .is_wysiwyg = "true";
defparam \register[10][31] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X62_Y41_N26
cycloneive_lcell_comb \Mux32~12 (
// Equation(s):
// \Mux32~12_combout  = (Selector10 & (Selector91)) # (!Selector10 & ((Selector91 & ((\register[10][31]~q ))) # (!Selector91 & (\register[8][31]~q ))))

	.dataa(Selector10),
	.datab(Selector91),
	.datac(\register[8][31]~q ),
	.datad(\register[10][31]~q ),
	.cin(gnd),
	.combout(\Mux32~12_combout ),
	.cout());
// synopsys translate_off
defparam \Mux32~12 .lut_mask = 16'hDC98;
defparam \Mux32~12 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X67_Y34_N18
cycloneive_lcell_comb \Mux32~13 (
// Equation(s):
// \Mux32~13_combout  = (Selector10 & ((\Mux32~12_combout  & (\register[11][31]~q )) # (!\Mux32~12_combout  & ((\register[9][31]~q ))))) # (!Selector10 & (((\Mux32~12_combout ))))

	.dataa(\register[11][31]~q ),
	.datab(\register[9][31]~q ),
	.datac(Selector10),
	.datad(\Mux32~12_combout ),
	.cin(gnd),
	.combout(\Mux32~13_combout ),
	.cout());
// synopsys translate_off
defparam \Mux32~13 .lut_mask = 16'hAFC0;
defparam \Mux32~13 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X67_Y34_N0
cycloneive_lcell_comb \Mux32~16 (
// Equation(s):
// \Mux32~16_combout  = (Selector8 & (Selector7)) # (!Selector8 & ((Selector7 & ((\Mux32~13_combout ))) # (!Selector7 & (\Mux32~15_combout ))))

	.dataa(Selector8),
	.datab(Selector7),
	.datac(\Mux32~15_combout ),
	.datad(\Mux32~13_combout ),
	.cin(gnd),
	.combout(\Mux32~16_combout ),
	.cout());
// synopsys translate_off
defparam \Mux32~16 .lut_mask = 16'hDC98;
defparam \Mux32~16 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X63_Y37_N24
cycloneive_lcell_comb \register~65 (
// Equation(s):
// \register~65_combout  = (WideOr01 & ((\wdat[30]~2_combout ) # ((plif_memwbregsrc_l_1 & plif_memwbrtnaddr_l_30))))

	.dataa(plif_memwbregsrc_l_1),
	.datab(plif_memwbrtnaddr_l_30),
	.datac(WideOr0),
	.datad(wdat_30),
	.cin(gnd),
	.combout(\register~65_combout ),
	.cout());
// synopsys translate_off
defparam \register~65 .lut_mask = 16'hF080;
defparam \register~65 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X65_Y37_N30
cycloneive_lcell_comb \Decoder0~35 (
// Equation(s):
// \Decoder0~35_combout  = (!plif_memwbwsel_l_0 & (!plif_memwbwsel_l_3 & (\Decoder0~21_combout  & plif_memwbwsel_l_4)))

	.dataa(plif_memwbwsel_l_0),
	.datab(plif_memwbwsel_l_3),
	.datac(\Decoder0~21_combout ),
	.datad(plif_memwbwsel_l_4),
	.cin(gnd),
	.combout(\Decoder0~35_combout ),
	.cout());
// synopsys translate_off
defparam \Decoder0~35 .lut_mask = 16'h1000;
defparam \Decoder0~35 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X65_Y39_N23
dffeas \register[20][30] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\register~65_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~35_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\register[20][30]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \register[20][30] .is_wysiwyg = "true";
defparam \register[20][30] .power_up = "low";
// synopsys translate_on

// Location: FF_X65_Y35_N15
dffeas \register[16][30] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\register~65_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~36_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\register[16][30]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \register[16][30] .is_wysiwyg = "true";
defparam \register[16][30] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X65_Y35_N14
cycloneive_lcell_comb \Mux33~4 (
// Equation(s):
// \Mux33~4_combout  = (Selector8 & (((Selector7)))) # (!Selector8 & ((Selector7 & (\register[24][30]~q )) # (!Selector7 & ((\register[16][30]~q )))))

	.dataa(\register[24][30]~q ),
	.datab(Selector8),
	.datac(\register[16][30]~q ),
	.datad(Selector7),
	.cin(gnd),
	.combout(\Mux33~4_combout ),
	.cout());
// synopsys translate_off
defparam \Mux33~4 .lut_mask = 16'hEE30;
defparam \Mux33~4 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X67_Y39_N18
cycloneive_lcell_comb \Mux33~5 (
// Equation(s):
// \Mux33~5_combout  = (Selector8 & ((\Mux33~4_combout  & (\register[28][30]~q )) # (!\Mux33~4_combout  & ((\register[20][30]~q ))))) # (!Selector8 & (((\Mux33~4_combout ))))

	.dataa(\register[28][30]~q ),
	.datab(\register[20][30]~q ),
	.datac(Selector8),
	.datad(\Mux33~4_combout ),
	.cin(gnd),
	.combout(\Mux33~5_combout ),
	.cout());
// synopsys translate_off
defparam \Mux33~5 .lut_mask = 16'hAFC0;
defparam \Mux33~5 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X69_Y35_N23
dffeas \register[18][30] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\register~65_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~33_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\register[18][30]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \register[18][30] .is_wysiwyg = "true";
defparam \register[18][30] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X69_Y35_N22
cycloneive_lcell_comb \Mux33~2 (
// Equation(s):
// \Mux33~2_combout  = (Selector8 & (((Selector7)))) # (!Selector8 & ((Selector7 & (\register[26][30]~q )) # (!Selector7 & ((\register[18][30]~q )))))

	.dataa(\register[26][30]~q ),
	.datab(Selector8),
	.datac(\register[18][30]~q ),
	.datad(Selector7),
	.cin(gnd),
	.combout(\Mux33~2_combout ),
	.cout());
// synopsys translate_off
defparam \Mux33~2 .lut_mask = 16'hEE30;
defparam \Mux33~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X67_Y39_N12
cycloneive_lcell_comb \register[30][30]~feeder (
// Equation(s):
// \register[30][30]~feeder_combout  = \register~65_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(\register~65_combout ),
	.cin(gnd),
	.combout(\register[30][30]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \register[30][30]~feeder .lut_mask = 16'hFF00;
defparam \register[30][30]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X67_Y39_N13
dffeas \register[30][30] (
	.clk(!CLK),
	.d(\register[30][30]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~56_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\register[30][30]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \register[30][30] .is_wysiwyg = "true";
defparam \register[30][30] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X67_Y39_N22
cycloneive_lcell_comb \Mux33~3 (
// Equation(s):
// \Mux33~3_combout  = (\Mux33~2_combout  & (((\register[30][30]~q ) # (!Selector8)))) # (!\Mux33~2_combout  & (\register[22][30]~q  & (Selector8)))

	.dataa(\register[22][30]~q ),
	.datab(\Mux33~2_combout ),
	.datac(Selector8),
	.datad(\register[30][30]~q ),
	.cin(gnd),
	.combout(\Mux33~3_combout ),
	.cout());
// synopsys translate_off
defparam \Mux33~3 .lut_mask = 16'hEC2C;
defparam \Mux33~3 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y39_N6
cycloneive_lcell_comb \Mux33~6 (
// Equation(s):
// \Mux33~6_combout  = (Selector10 & (((Selector91)))) # (!Selector10 & ((Selector91 & ((\Mux33~3_combout ))) # (!Selector91 & (\Mux33~5_combout ))))

	.dataa(\Mux33~5_combout ),
	.datab(Selector10),
	.datac(Selector91),
	.datad(\Mux33~3_combout ),
	.cin(gnd),
	.combout(\Mux33~6_combout ),
	.cout());
// synopsys translate_off
defparam \Mux33~6 .lut_mask = 16'hF2C2;
defparam \Mux33~6 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X62_Y39_N7
dffeas \register[27][30] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\register~65_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~38_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\register[27][30]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \register[27][30] .is_wysiwyg = "true";
defparam \register[27][30] .power_up = "low";
// synopsys translate_on

// Location: FF_X62_Y39_N17
dffeas \register[31][30] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\register~65_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~40_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\register[31][30]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \register[31][30] .is_wysiwyg = "true";
defparam \register[31][30] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X62_Y38_N0
cycloneive_lcell_comb \register[23][30]~feeder (
// Equation(s):
// \register[23][30]~feeder_combout  = \register~65_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(\register~65_combout ),
	.cin(gnd),
	.combout(\register[23][30]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \register[23][30]~feeder .lut_mask = 16'hFF00;
defparam \register[23][30]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X62_Y38_N1
dffeas \register[23][30] (
	.clk(!CLK),
	.d(\register[23][30]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~37_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\register[23][30]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \register[23][30] .is_wysiwyg = "true";
defparam \register[23][30] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X62_Y38_N2
cycloneive_lcell_comb \register[19][30]~feeder (
// Equation(s):
// \register[19][30]~feeder_combout  = \register~65_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(\register~65_combout ),
	.cin(gnd),
	.combout(\register[19][30]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \register[19][30]~feeder .lut_mask = 16'hFF00;
defparam \register[19][30]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X62_Y38_N3
dffeas \register[19][30] (
	.clk(!CLK),
	.d(\register[19][30]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~39_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\register[19][30]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \register[19][30] .is_wysiwyg = "true";
defparam \register[19][30] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X62_Y38_N8
cycloneive_lcell_comb \Mux33~7 (
// Equation(s):
// \Mux33~7_combout  = (Selector7 & (((Selector8)))) # (!Selector7 & ((Selector8 & (\register[23][30]~q )) # (!Selector8 & ((\register[19][30]~q )))))

	.dataa(Selector7),
	.datab(\register[23][30]~q ),
	.datac(Selector8),
	.datad(\register[19][30]~q ),
	.cin(gnd),
	.combout(\Mux33~7_combout ),
	.cout());
// synopsys translate_off
defparam \Mux33~7 .lut_mask = 16'hE5E0;
defparam \Mux33~7 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y39_N8
cycloneive_lcell_comb \Mux33~8 (
// Equation(s):
// \Mux33~8_combout  = (\Mux33~7_combout  & (((\register[31][30]~q ) # (!Selector7)))) # (!\Mux33~7_combout  & (\register[27][30]~q  & ((Selector7))))

	.dataa(\register[27][30]~q ),
	.datab(\register[31][30]~q ),
	.datac(\Mux33~7_combout ),
	.datad(Selector7),
	.cin(gnd),
	.combout(\Mux33~8_combout ),
	.cout());
// synopsys translate_off
defparam \Mux33~8 .lut_mask = 16'hCAF0;
defparam \Mux33~8 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X63_Y37_N4
cycloneive_lcell_comb \register[25][30]~feeder (
// Equation(s):
// \register[25][30]~feeder_combout  = \register~65_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(\register~65_combout ),
	.cin(gnd),
	.combout(\register[25][30]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \register[25][30]~feeder .lut_mask = 16'hFF00;
defparam \register[25][30]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X63_Y37_N5
dffeas \register[25][30] (
	.clk(!CLK),
	.d(\register[25][30]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~24_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\register[25][30]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \register[25][30] .is_wysiwyg = "true";
defparam \register[25][30] .power_up = "low";
// synopsys translate_on

// Location: FF_X63_Y33_N21
dffeas \register[21][30] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\register~65_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~22_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\register[21][30]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \register[21][30] .is_wysiwyg = "true";
defparam \register[21][30] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X63_Y33_N20
cycloneive_lcell_comb \Mux33~0 (
// Equation(s):
// \Mux33~0_combout  = (Selector8 & (((\register[21][30]~q ) # (Selector7)))) # (!Selector8 & (\register[17][30]~q  & ((!Selector7))))

	.dataa(\register[17][30]~q ),
	.datab(Selector8),
	.datac(\register[21][30]~q ),
	.datad(Selector7),
	.cin(gnd),
	.combout(\Mux33~0_combout ),
	.cout());
// synopsys translate_off
defparam \Mux33~0 .lut_mask = 16'hCCE2;
defparam \Mux33~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X63_Y33_N3
dffeas \register[29][30] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\register~65_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~28_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\register[29][30]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \register[29][30] .is_wysiwyg = "true";
defparam \register[29][30] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X61_Y39_N4
cycloneive_lcell_comb \Mux33~1 (
// Equation(s):
// \Mux33~1_combout  = (Selector7 & ((\Mux33~0_combout  & ((\register[29][30]~q ))) # (!\Mux33~0_combout  & (\register[25][30]~q )))) # (!Selector7 & (((\Mux33~0_combout ))))

	.dataa(Selector7),
	.datab(\register[25][30]~q ),
	.datac(\Mux33~0_combout ),
	.datad(\register[29][30]~q ),
	.cin(gnd),
	.combout(\Mux33~1_combout ),
	.cout());
// synopsys translate_off
defparam \Mux33~1 .lut_mask = 16'hF858;
defparam \Mux33~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X62_Y32_N3
dffeas \register[14][30] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\register~65_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~61_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\register[14][30]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \register[14][30] .is_wysiwyg = "true";
defparam \register[14][30] .power_up = "low";
// synopsys translate_on

// Location: FF_X63_Y37_N27
dffeas \register[15][30] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\register~65_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~53_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\register[15][30]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \register[15][30] .is_wysiwyg = "true";
defparam \register[15][30] .power_up = "low";
// synopsys translate_on

// Location: FF_X62_Y30_N9
dffeas \register[13][30] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\register~65_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~62_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\register[13][30]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \register[13][30] .is_wysiwyg = "true";
defparam \register[13][30] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X62_Y37_N2
cycloneive_lcell_comb \Decoder0~31 (
// Equation(s):
// \Decoder0~31_combout  = (plif_memwbwsel_l_2 & !plif_memwbwsel_l_0)

	.dataa(gnd),
	.datab(gnd),
	.datac(plif_memwbwsel_l_2),
	.datad(plif_memwbwsel_l_0),
	.cin(gnd),
	.combout(\Decoder0~31_combout ),
	.cout());
// synopsys translate_off
defparam \Decoder0~31 .lut_mask = 16'h00F0;
defparam \Decoder0~31 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y37_N8
cycloneive_lcell_comb \Decoder0~52 (
// Equation(s):
// \Decoder0~52_combout  = (\Decoder0~23_combout  & (!plif_memwbwsel_l_4 & (!plif_memwbwsel_l_1 & \Decoder0~31_combout )))

	.dataa(\Decoder0~23_combout ),
	.datab(plif_memwbwsel_l_4),
	.datac(plif_memwbwsel_l_1),
	.datad(\Decoder0~31_combout ),
	.cin(gnd),
	.combout(\Decoder0~52_combout ),
	.cout());
// synopsys translate_off
defparam \Decoder0~52 .lut_mask = 16'h0200;
defparam \Decoder0~52 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X62_Y30_N11
dffeas \register[12][30] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\register~65_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~52_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\register[12][30]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \register[12][30] .is_wysiwyg = "true";
defparam \register[12][30] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X62_Y30_N10
cycloneive_lcell_comb \Mux33~17 (
// Equation(s):
// \Mux33~17_combout  = (Selector10 & ((\register[13][30]~q ) # ((Selector91)))) # (!Selector10 & (((\register[12][30]~q  & !Selector91))))

	.dataa(Selector10),
	.datab(\register[13][30]~q ),
	.datac(\register[12][30]~q ),
	.datad(Selector91),
	.cin(gnd),
	.combout(\Mux33~17_combout ),
	.cout());
// synopsys translate_off
defparam \Mux33~17 .lut_mask = 16'hAAD8;
defparam \Mux33~17 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X63_Y37_N26
cycloneive_lcell_comb \Mux33~18 (
// Equation(s):
// \Mux33~18_combout  = (Selector91 & ((\Mux33~17_combout  & ((\register[15][30]~q ))) # (!\Mux33~17_combout  & (\register[14][30]~q )))) # (!Selector91 & (((\Mux33~17_combout ))))

	.dataa(\register[14][30]~q ),
	.datab(Selector91),
	.datac(\register[15][30]~q ),
	.datad(\Mux33~17_combout ),
	.cin(gnd),
	.combout(\Mux33~18_combout ),
	.cout());
// synopsys translate_off
defparam \Mux33~18 .lut_mask = 16'hF388;
defparam \Mux33~18 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X62_Y41_N9
dffeas \register[10][30] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\register~65_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~45_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\register[10][30]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \register[10][30] .is_wysiwyg = "true";
defparam \register[10][30] .power_up = "low";
// synopsys translate_on

// Location: FF_X62_Y41_N19
dffeas \register[8][30] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\register~65_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~46_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\register[8][30]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \register[8][30] .is_wysiwyg = "true";
defparam \register[8][30] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X62_Y41_N18
cycloneive_lcell_comb \Mux33~10 (
// Equation(s):
// \Mux33~10_combout  = (Selector10 & (((Selector91)))) # (!Selector10 & ((Selector91 & (\register[10][30]~q )) # (!Selector91 & ((\register[8][30]~q )))))

	.dataa(Selector10),
	.datab(\register[10][30]~q ),
	.datac(\register[8][30]~q ),
	.datad(Selector91),
	.cin(gnd),
	.combout(\Mux33~10_combout ),
	.cout());
// synopsys translate_off
defparam \Mux33~10 .lut_mask = 16'hEE50;
defparam \Mux33~10 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y37_N22
cycloneive_lcell_comb \Decoder0~47 (
// Equation(s):
// \Decoder0~47_combout  = (!plif_memwbwsel_l_2 & (!plif_memwbwsel_l_4 & (plif_memwbwsel_l_0 & \Decoder0~29_combout )))

	.dataa(plif_memwbwsel_l_2),
	.datab(plif_memwbwsel_l_4),
	.datac(plif_memwbwsel_l_0),
	.datad(\Decoder0~29_combout ),
	.cin(gnd),
	.combout(\Decoder0~47_combout ),
	.cout());
// synopsys translate_off
defparam \Decoder0~47 .lut_mask = 16'h1000;
defparam \Decoder0~47 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X66_Y38_N25
dffeas \register[11][30] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\register~65_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~47_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\register[11][30]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \register[11][30] .is_wysiwyg = "true";
defparam \register[11][30] .power_up = "low";
// synopsys translate_on

// Location: FF_X66_Y38_N11
dffeas \register[9][30] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\register~65_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~44_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\register[9][30]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \register[9][30] .is_wysiwyg = "true";
defparam \register[9][30] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X66_Y38_N10
cycloneive_lcell_comb \Mux33~11 (
// Equation(s):
// \Mux33~11_combout  = (\Mux33~10_combout  & ((\register[11][30]~q ) # ((!Selector10)))) # (!\Mux33~10_combout  & (((\register[9][30]~q  & Selector10))))

	.dataa(\Mux33~10_combout ),
	.datab(\register[11][30]~q ),
	.datac(\register[9][30]~q ),
	.datad(Selector10),
	.cin(gnd),
	.combout(\Mux33~11_combout ),
	.cout());
// synopsys translate_off
defparam \Mux33~11 .lut_mask = 16'hD8AA;
defparam \Mux33~11 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X68_Y31_N21
dffeas \register[6][30] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\register~65_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~58_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\register[6][30]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \register[6][30] .is_wysiwyg = "true";
defparam \register[6][30] .power_up = "low";
// synopsys translate_on

// Location: FF_X68_Y31_N7
dffeas \register[7][30] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\register~65_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~43_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\register[7][30]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \register[7][30] .is_wysiwyg = "true";
defparam \register[7][30] .power_up = "low";
// synopsys translate_on

// Location: FF_X69_Y31_N5
dffeas \register[5][30] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\register~65_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~59_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\register[5][30]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \register[5][30] .is_wysiwyg = "true";
defparam \register[5][30] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X69_Y31_N4
cycloneive_lcell_comb \Mux33~12 (
// Equation(s):
// \Mux33~12_combout  = (Selector91 & (((Selector10)))) # (!Selector91 & ((Selector10 & ((\register[5][30]~q ))) # (!Selector10 & (\register[4][30]~q ))))

	.dataa(\register[4][30]~q ),
	.datab(Selector91),
	.datac(\register[5][30]~q ),
	.datad(Selector10),
	.cin(gnd),
	.combout(\Mux33~12_combout ),
	.cout());
// synopsys translate_off
defparam \Mux33~12 .lut_mask = 16'hFC22;
defparam \Mux33~12 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X68_Y31_N6
cycloneive_lcell_comb \Mux33~13 (
// Equation(s):
// \Mux33~13_combout  = (Selector91 & ((\Mux33~12_combout  & ((\register[7][30]~q ))) # (!\Mux33~12_combout  & (\register[6][30]~q )))) # (!Selector91 & (((\Mux33~12_combout ))))

	.dataa(Selector91),
	.datab(\register[6][30]~q ),
	.datac(\register[7][30]~q ),
	.datad(\Mux33~12_combout ),
	.cin(gnd),
	.combout(\Mux33~13_combout ),
	.cout());
// synopsys translate_off
defparam \Mux33~13 .lut_mask = 16'hF588;
defparam \Mux33~13 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X66_Y34_N13
dffeas \register[2][30] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\register~65_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~50_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\register[2][30]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \register[2][30] .is_wysiwyg = "true";
defparam \register[2][30] .power_up = "low";
// synopsys translate_on

// Location: FF_X65_Y33_N17
dffeas \register[3][30] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\register~65_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~48_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\register[3][30]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \register[3][30] .is_wysiwyg = "true";
defparam \register[3][30] .power_up = "low";
// synopsys translate_on

// Location: FF_X65_Y33_N27
dffeas \register[1][30] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\register~65_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~49_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\register[1][30]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \register[1][30] .is_wysiwyg = "true";
defparam \register[1][30] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X65_Y33_N26
cycloneive_lcell_comb \Mux33~14 (
// Equation(s):
// \Mux33~14_combout  = (Selector10 & ((Selector91 & (\register[3][30]~q )) # (!Selector91 & ((\register[1][30]~q )))))

	.dataa(Selector91),
	.datab(\register[3][30]~q ),
	.datac(\register[1][30]~q ),
	.datad(Selector10),
	.cin(gnd),
	.combout(\Mux33~14_combout ),
	.cout());
// synopsys translate_off
defparam \Mux33~14 .lut_mask = 16'hD800;
defparam \Mux33~14 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X65_Y32_N24
cycloneive_lcell_comb \Mux33~15 (
// Equation(s):
// \Mux33~15_combout  = (\Mux33~14_combout ) # ((!Selector10 & (\register[2][30]~q  & Selector91)))

	.dataa(Selector10),
	.datab(\register[2][30]~q ),
	.datac(\Mux33~14_combout ),
	.datad(Selector91),
	.cin(gnd),
	.combout(\Mux33~15_combout ),
	.cout());
// synopsys translate_off
defparam \Mux33~15 .lut_mask = 16'hF4F0;
defparam \Mux33~15 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X65_Y32_N22
cycloneive_lcell_comb \Mux33~16 (
// Equation(s):
// \Mux33~16_combout  = (Selector7 & (((Selector8)))) # (!Selector7 & ((Selector8 & (\Mux33~13_combout )) # (!Selector8 & ((\Mux33~15_combout )))))

	.dataa(\Mux33~13_combout ),
	.datab(Selector7),
	.datac(Selector8),
	.datad(\Mux33~15_combout ),
	.cin(gnd),
	.combout(\Mux33~16_combout ),
	.cout());
// synopsys translate_off
defparam \Mux33~16 .lut_mask = 16'hE3E0;
defparam \Mux33~16 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y35_N26
cycloneive_lcell_comb \register~66 (
// Equation(s):
// \register~66_combout  = (WideOr01 & ((\wdat[29]~4_combout ) # ((plif_memwbrtnaddr_l_29 & plif_memwbregsrc_l_1))))

	.dataa(plif_memwbrtnaddr_l_29),
	.datab(WideOr0),
	.datac(wdat_29),
	.datad(plif_memwbregsrc_l_1),
	.cin(gnd),
	.combout(\register~66_combout ),
	.cout());
// synopsys translate_off
defparam \register~66 .lut_mask = 16'hC8C0;
defparam \register~66 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X61_Y33_N13
dffeas \register[31][29] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\register~66_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~40_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\register[31][29]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \register[31][29] .is_wysiwyg = "true";
defparam \register[31][29] .power_up = "low";
// synopsys translate_on

// Location: FF_X60_Y35_N13
dffeas \register[23][29] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\register~66_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~37_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\register[23][29]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \register[23][29] .is_wysiwyg = "true";
defparam \register[23][29] .power_up = "low";
// synopsys translate_on

// Location: FF_X60_Y38_N9
dffeas \register[19][29] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\register~66_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~39_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\register[19][29]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \register[19][29] .is_wysiwyg = "true";
defparam \register[19][29] .power_up = "low";
// synopsys translate_on

// Location: FF_X63_Y35_N21
dffeas \register[27][29] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\register~66_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~38_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\register[27][29]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \register[27][29] .is_wysiwyg = "true";
defparam \register[27][29] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X63_Y35_N20
cycloneive_lcell_comb \Mux34~7 (
// Equation(s):
// \Mux34~7_combout  = (Selector7 & (((\register[27][29]~q ) # (Selector8)))) # (!Selector7 & (\register[19][29]~q  & ((!Selector8))))

	.dataa(Selector7),
	.datab(\register[19][29]~q ),
	.datac(\register[27][29]~q ),
	.datad(Selector8),
	.cin(gnd),
	.combout(\Mux34~7_combout ),
	.cout());
// synopsys translate_off
defparam \Mux34~7 .lut_mask = 16'hAAE4;
defparam \Mux34~7 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y35_N12
cycloneive_lcell_comb \Mux34~8 (
// Equation(s):
// \Mux34~8_combout  = (Selector8 & ((\Mux34~7_combout  & (\register[31][29]~q )) # (!\Mux34~7_combout  & ((\register[23][29]~q ))))) # (!Selector8 & (((\Mux34~7_combout ))))

	.dataa(\register[31][29]~q ),
	.datab(Selector8),
	.datac(\register[23][29]~q ),
	.datad(\Mux34~7_combout ),
	.cin(gnd),
	.combout(\Mux34~8_combout ),
	.cout());
// synopsys translate_off
defparam \Mux34~8 .lut_mask = 16'hBBC0;
defparam \Mux34~8 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y31_N22
cycloneive_lcell_comb \register[29][29]~feeder (
// Equation(s):
// \register[29][29]~feeder_combout  = \register~66_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(\register~66_combout ),
	.cin(gnd),
	.combout(\register[29][29]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \register[29][29]~feeder .lut_mask = 16'hFF00;
defparam \register[29][29]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X61_Y31_N23
dffeas \register[29][29] (
	.clk(!CLK),
	.d(\register[29][29]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~28_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\register[29][29]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \register[29][29] .is_wysiwyg = "true";
defparam \register[29][29] .power_up = "low";
// synopsys translate_on

// Location: FF_X61_Y35_N27
dffeas \register[21][29] (
	.clk(!CLK),
	.d(\register~66_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~22_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\register[21][29]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \register[21][29] .is_wysiwyg = "true";
defparam \register[21][29] .power_up = "low";
// synopsys translate_on

// Location: FF_X61_Y37_N11
dffeas \register[25][29] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\register~66_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~24_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\register[25][29]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \register[25][29] .is_wysiwyg = "true";
defparam \register[25][29] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X58_Y37_N12
cycloneive_lcell_comb \Decoder0~26 (
// Equation(s):
// \Decoder0~26_combout  = (plif_memwbwsel_l_0 & \Decoder0~25_combout )

	.dataa(plif_memwbwsel_l_0),
	.datab(gnd),
	.datac(gnd),
	.datad(\Decoder0~25_combout ),
	.cin(gnd),
	.combout(\Decoder0~26_combout ),
	.cout());
// synopsys translate_off
defparam \Decoder0~26 .lut_mask = 16'hAA00;
defparam \Decoder0~26 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X62_Y35_N5
dffeas \register[17][29] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\register~66_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~26_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\register[17][29]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \register[17][29] .is_wysiwyg = "true";
defparam \register[17][29] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X61_Y37_N10
cycloneive_lcell_comb \Mux34~0 (
// Equation(s):
// \Mux34~0_combout  = (Selector7 & ((Selector8) # ((\register[25][29]~q )))) # (!Selector7 & (!Selector8 & ((\register[17][29]~q ))))

	.dataa(Selector7),
	.datab(Selector8),
	.datac(\register[25][29]~q ),
	.datad(\register[17][29]~q ),
	.cin(gnd),
	.combout(\Mux34~0_combout ),
	.cout());
// synopsys translate_off
defparam \Mux34~0 .lut_mask = 16'hB9A8;
defparam \Mux34~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y32_N12
cycloneive_lcell_comb \Mux34~1 (
// Equation(s):
// \Mux34~1_combout  = (Selector8 & ((\Mux34~0_combout  & (\register[29][29]~q )) # (!\Mux34~0_combout  & ((\register[21][29]~q ))))) # (!Selector8 & (((\Mux34~0_combout ))))

	.dataa(Selector8),
	.datab(\register[29][29]~q ),
	.datac(\register[21][29]~q ),
	.datad(\Mux34~0_combout ),
	.cin(gnd),
	.combout(\Mux34~1_combout ),
	.cout());
// synopsys translate_off
defparam \Mux34~1 .lut_mask = 16'hDDA0;
defparam \Mux34~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X69_Y35_N9
dffeas \register[22][29] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\register~66_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~55_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\register[22][29]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \register[22][29] .is_wysiwyg = "true";
defparam \register[22][29] .power_up = "low";
// synopsys translate_on

// Location: FF_X69_Y35_N7
dffeas \register[18][29] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\register~66_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~33_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\register[18][29]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \register[18][29] .is_wysiwyg = "true";
defparam \register[18][29] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X69_Y35_N8
cycloneive_lcell_comb \Mux34~2 (
// Equation(s):
// \Mux34~2_combout  = (Selector7 & (Selector8)) # (!Selector7 & ((Selector8 & (\register[22][29]~q )) # (!Selector8 & ((\register[18][29]~q )))))

	.dataa(Selector7),
	.datab(Selector8),
	.datac(\register[22][29]~q ),
	.datad(\register[18][29]~q ),
	.cin(gnd),
	.combout(\Mux34~2_combout ),
	.cout());
// synopsys translate_off
defparam \Mux34~2 .lut_mask = 16'hD9C8;
defparam \Mux34~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X68_Y35_N17
dffeas \register[26][29] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\register~66_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~54_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\register[26][29]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \register[26][29] .is_wysiwyg = "true";
defparam \register[26][29] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X68_Y35_N16
cycloneive_lcell_comb \Mux34~3 (
// Equation(s):
// \Mux34~3_combout  = (\Mux34~2_combout  & ((\register[30][29]~q ) # ((!Selector7)))) # (!\Mux34~2_combout  & (((\register[26][29]~q  & Selector7))))

	.dataa(\register[30][29]~q ),
	.datab(\Mux34~2_combout ),
	.datac(\register[26][29]~q ),
	.datad(Selector7),
	.cin(gnd),
	.combout(\Mux34~3_combout ),
	.cout());
// synopsys translate_off
defparam \Mux34~3 .lut_mask = 16'hB8CC;
defparam \Mux34~3 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X66_Y35_N21
dffeas \register[28][29] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\register~66_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~57_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\register[28][29]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \register[28][29] .is_wysiwyg = "true";
defparam \register[28][29] .power_up = "low";
// synopsys translate_on

// Location: FF_X65_Y35_N19
dffeas \register[16][29] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\register~66_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~36_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\register[16][29]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \register[16][29] .is_wysiwyg = "true";
defparam \register[16][29] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X65_Y39_N28
cycloneive_lcell_comb \register[20][29]~feeder (
// Equation(s):
// \register[20][29]~feeder_combout  = \register~66_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(\register~66_combout ),
	.cin(gnd),
	.combout(\register[20][29]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \register[20][29]~feeder .lut_mask = 16'hFF00;
defparam \register[20][29]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X65_Y39_N29
dffeas \register[20][29] (
	.clk(!CLK),
	.d(\register[20][29]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~35_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\register[20][29]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \register[20][29] .is_wysiwyg = "true";
defparam \register[20][29] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X65_Y35_N18
cycloneive_lcell_comb \Mux34~4 (
// Equation(s):
// \Mux34~4_combout  = (Selector7 & (Selector8)) # (!Selector7 & ((Selector8 & ((\register[20][29]~q ))) # (!Selector8 & (\register[16][29]~q ))))

	.dataa(Selector7),
	.datab(Selector8),
	.datac(\register[16][29]~q ),
	.datad(\register[20][29]~q ),
	.cin(gnd),
	.combout(\Mux34~4_combout ),
	.cout());
// synopsys translate_off
defparam \Mux34~4 .lut_mask = 16'hDC98;
defparam \Mux34~4 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y32_N2
cycloneive_lcell_comb \Mux34~5 (
// Equation(s):
// \Mux34~5_combout  = (\Mux34~4_combout  & (((\register[28][29]~q ) # (!Selector7)))) # (!\Mux34~4_combout  & (\register[24][29]~q  & ((Selector7))))

	.dataa(\register[24][29]~q ),
	.datab(\register[28][29]~q ),
	.datac(\Mux34~4_combout ),
	.datad(Selector7),
	.cin(gnd),
	.combout(\Mux34~5_combout ),
	.cout());
// synopsys translate_off
defparam \Mux34~5 .lut_mask = 16'hCAF0;
defparam \Mux34~5 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y32_N28
cycloneive_lcell_comb \Mux34~6 (
// Equation(s):
// \Mux34~6_combout  = (Selector10 & (((Selector91)))) # (!Selector10 & ((Selector91 & (\Mux34~3_combout )) # (!Selector91 & ((\Mux34~5_combout )))))

	.dataa(Selector10),
	.datab(\Mux34~3_combout ),
	.datac(Selector91),
	.datad(\Mux34~5_combout ),
	.cin(gnd),
	.combout(\Mux34~6_combout ),
	.cout());
// synopsys translate_off
defparam \Mux34~6 .lut_mask = 16'hE5E0;
defparam \Mux34~6 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X60_Y36_N9
dffeas \register[14][29] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\register~66_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~61_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\register[14][29]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \register[14][29] .is_wysiwyg = "true";
defparam \register[14][29] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X61_Y35_N8
cycloneive_lcell_comb \register[15][29]~feeder (
// Equation(s):
// \register[15][29]~feeder_combout  = \register~66_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(\register~66_combout ),
	.datad(gnd),
	.cin(gnd),
	.combout(\register[15][29]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \register[15][29]~feeder .lut_mask = 16'hF0F0;
defparam \register[15][29]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X61_Y35_N9
dffeas \register[15][29] (
	.clk(!CLK),
	.d(\register[15][29]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~53_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\register[15][29]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \register[15][29] .is_wysiwyg = "true";
defparam \register[15][29] .power_up = "low";
// synopsys translate_on

// Location: FF_X60_Y36_N31
dffeas \register[12][29] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\register~66_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~52_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\register[12][29]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \register[12][29] .is_wysiwyg = "true";
defparam \register[12][29] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X59_Y36_N20
cycloneive_lcell_comb \register[13][29]~feeder (
// Equation(s):
// \register[13][29]~feeder_combout  = \register~66_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(\register~66_combout ),
	.datad(gnd),
	.cin(gnd),
	.combout(\register[13][29]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \register[13][29]~feeder .lut_mask = 16'hF0F0;
defparam \register[13][29]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X59_Y36_N21
dffeas \register[13][29] (
	.clk(!CLK),
	.d(\register[13][29]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~62_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\register[13][29]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \register[13][29] .is_wysiwyg = "true";
defparam \register[13][29] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X60_Y36_N30
cycloneive_lcell_comb \Mux34~17 (
// Equation(s):
// \Mux34~17_combout  = (Selector91 & (Selector10)) # (!Selector91 & ((Selector10 & ((\register[13][29]~q ))) # (!Selector10 & (\register[12][29]~q ))))

	.dataa(Selector91),
	.datab(Selector10),
	.datac(\register[12][29]~q ),
	.datad(\register[13][29]~q ),
	.cin(gnd),
	.combout(\Mux34~17_combout ),
	.cout());
// synopsys translate_off
defparam \Mux34~17 .lut_mask = 16'hDC98;
defparam \Mux34~17 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y35_N6
cycloneive_lcell_comb \Mux34~18 (
// Equation(s):
// \Mux34~18_combout  = (\Mux34~17_combout  & (((\register[15][29]~q ) # (!Selector91)))) # (!\Mux34~17_combout  & (\register[14][29]~q  & ((Selector91))))

	.dataa(\register[14][29]~q ),
	.datab(\register[15][29]~q ),
	.datac(\Mux34~17_combout ),
	.datad(Selector91),
	.cin(gnd),
	.combout(\Mux34~18_combout ),
	.cout());
// synopsys translate_off
defparam \Mux34~18 .lut_mask = 16'hCAF0;
defparam \Mux34~18 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X66_Y31_N27
dffeas \register[7][29] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\register~66_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~43_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\register[7][29]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \register[7][29] .is_wysiwyg = "true";
defparam \register[7][29] .power_up = "low";
// synopsys translate_on

// Location: FF_X66_Y31_N5
dffeas \register[6][29] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\register~66_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~58_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\register[6][29]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \register[6][29] .is_wysiwyg = "true";
defparam \register[6][29] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X66_Y37_N22
cycloneive_lcell_comb \Decoder0~60 (
// Equation(s):
// \Decoder0~60_combout  = (!plif_memwbwsel_l_4 & (!plif_memwbwsel_l_0 & (!plif_memwbwsel_l_3 & \Decoder0~21_combout )))

	.dataa(plif_memwbwsel_l_4),
	.datab(plif_memwbwsel_l_0),
	.datac(plif_memwbwsel_l_3),
	.datad(\Decoder0~21_combout ),
	.cin(gnd),
	.combout(\Decoder0~60_combout ),
	.cout());
// synopsys translate_off
defparam \Decoder0~60 .lut_mask = 16'h0100;
defparam \Decoder0~60 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X69_Y31_N15
dffeas \register[4][29] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\register~66_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~60_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\register[4][29]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \register[4][29] .is_wysiwyg = "true";
defparam \register[4][29] .power_up = "low";
// synopsys translate_on

// Location: FF_X69_Y31_N13
dffeas \register[5][29] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\register~66_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~59_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\register[5][29]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \register[5][29] .is_wysiwyg = "true";
defparam \register[5][29] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X69_Y31_N14
cycloneive_lcell_comb \Mux34~10 (
// Equation(s):
// \Mux34~10_combout  = (Selector10 & ((Selector91) # ((\register[5][29]~q )))) # (!Selector10 & (!Selector91 & (\register[4][29]~q )))

	.dataa(Selector10),
	.datab(Selector91),
	.datac(\register[4][29]~q ),
	.datad(\register[5][29]~q ),
	.cin(gnd),
	.combout(\Mux34~10_combout ),
	.cout());
// synopsys translate_off
defparam \Mux34~10 .lut_mask = 16'hBA98;
defparam \Mux34~10 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X66_Y31_N4
cycloneive_lcell_comb \Mux34~11 (
// Equation(s):
// \Mux34~11_combout  = (Selector91 & ((\Mux34~10_combout  & (\register[7][29]~q )) # (!\Mux34~10_combout  & ((\register[6][29]~q ))))) # (!Selector91 & (((\Mux34~10_combout ))))

	.dataa(\register[7][29]~q ),
	.datab(Selector91),
	.datac(\register[6][29]~q ),
	.datad(\Mux34~10_combout ),
	.cin(gnd),
	.combout(\Mux34~11_combout ),
	.cout());
// synopsys translate_off
defparam \Mux34~11 .lut_mask = 16'hBBC0;
defparam \Mux34~11 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X66_Y32_N0
cycloneive_lcell_comb \register[2][29]~feeder (
// Equation(s):
// \register[2][29]~feeder_combout  = \register~66_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(\register~66_combout ),
	.cin(gnd),
	.combout(\register[2][29]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \register[2][29]~feeder .lut_mask = 16'hFF00;
defparam \register[2][29]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X66_Y32_N1
dffeas \register[2][29] (
	.clk(!CLK),
	.d(\register[2][29]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~50_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\register[2][29]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \register[2][29] .is_wysiwyg = "true";
defparam \register[2][29] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X66_Y32_N22
cycloneive_lcell_comb \Mux34~15 (
// Equation(s):
// \Mux34~15_combout  = (Selector10 & (\Mux34~14_combout )) # (!Selector10 & (((\register[2][29]~q  & Selector91))))

	.dataa(\Mux34~14_combout ),
	.datab(\register[2][29]~q ),
	.datac(Selector91),
	.datad(Selector10),
	.cin(gnd),
	.combout(\Mux34~15_combout ),
	.cout());
// synopsys translate_off
defparam \Mux34~15 .lut_mask = 16'hAAC0;
defparam \Mux34~15 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X65_Y40_N1
dffeas \register[9][29] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\register~66_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~44_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\register[9][29]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \register[9][29] .is_wysiwyg = "true";
defparam \register[9][29] .power_up = "low";
// synopsys translate_on

// Location: FF_X65_Y40_N27
dffeas \register[11][29] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\register~66_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~47_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\register[11][29]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \register[11][29] .is_wysiwyg = "true";
defparam \register[11][29] .power_up = "low";
// synopsys translate_on

// Location: FF_X62_Y41_N21
dffeas \register[10][29] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\register~66_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~45_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\register[10][29]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \register[10][29] .is_wysiwyg = "true";
defparam \register[10][29] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X62_Y41_N20
cycloneive_lcell_comb \Mux34~12 (
// Equation(s):
// \Mux34~12_combout  = (Selector91 & (((\register[10][29]~q ) # (Selector10)))) # (!Selector91 & (\register[8][29]~q  & ((!Selector10))))

	.dataa(\register[8][29]~q ),
	.datab(Selector91),
	.datac(\register[10][29]~q ),
	.datad(Selector10),
	.cin(gnd),
	.combout(\Mux34~12_combout ),
	.cout());
// synopsys translate_off
defparam \Mux34~12 .lut_mask = 16'hCCE2;
defparam \Mux34~12 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X65_Y40_N26
cycloneive_lcell_comb \Mux34~13 (
// Equation(s):
// \Mux34~13_combout  = (Selector10 & ((\Mux34~12_combout  & ((\register[11][29]~q ))) # (!\Mux34~12_combout  & (\register[9][29]~q )))) # (!Selector10 & (((\Mux34~12_combout ))))

	.dataa(Selector10),
	.datab(\register[9][29]~q ),
	.datac(\register[11][29]~q ),
	.datad(\Mux34~12_combout ),
	.cin(gnd),
	.combout(\Mux34~13_combout ),
	.cout());
// synopsys translate_off
defparam \Mux34~13 .lut_mask = 16'hF588;
defparam \Mux34~13 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y32_N24
cycloneive_lcell_comb \Mux34~16 (
// Equation(s):
// \Mux34~16_combout  = (Selector8 & (Selector7)) # (!Selector8 & ((Selector7 & ((\Mux34~13_combout ))) # (!Selector7 & (\Mux34~15_combout ))))

	.dataa(Selector8),
	.datab(Selector7),
	.datac(\Mux34~15_combout ),
	.datad(\Mux34~13_combout ),
	.cin(gnd),
	.combout(\Mux34~16_combout ),
	.cout());
// synopsys translate_off
defparam \Mux34~16 .lut_mask = 16'hDC98;
defparam \Mux34~16 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X63_Y37_N12
cycloneive_lcell_comb \register~67 (
// Equation(s):
// \register~67_combout  = (WideOr01 & ((\wdat[28]~6_combout ) # ((plif_memwbregsrc_l_1 & plif_memwbrtnaddr_l_28))))

	.dataa(plif_memwbregsrc_l_1),
	.datab(plif_memwbrtnaddr_l_28),
	.datac(WideOr0),
	.datad(wdat_28),
	.cin(gnd),
	.combout(\register~67_combout ),
	.cout());
// synopsys translate_off
defparam \register~67 .lut_mask = 16'hF080;
defparam \register~67 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X67_Y35_N10
cycloneive_lcell_comb \register[27][28]~feeder (
// Equation(s):
// \register[27][28]~feeder_combout  = \register~67_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(\register~67_combout ),
	.cin(gnd),
	.combout(\register[27][28]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \register[27][28]~feeder .lut_mask = 16'hFF00;
defparam \register[27][28]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X67_Y35_N11
dffeas \register[27][28] (
	.clk(!CLK),
	.d(\register[27][28]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~38_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\register[27][28]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \register[27][28] .is_wysiwyg = "true";
defparam \register[27][28] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X62_Y35_N20
cycloneive_lcell_comb \register[31][28]~feeder (
// Equation(s):
// \register[31][28]~feeder_combout  = \register~67_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(\register~67_combout ),
	.cin(gnd),
	.combout(\register[31][28]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \register[31][28]~feeder .lut_mask = 16'hFF00;
defparam \register[31][28]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X62_Y35_N21
dffeas \register[31][28] (
	.clk(!CLK),
	.d(\register[31][28]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~40_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\register[31][28]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \register[31][28] .is_wysiwyg = "true";
defparam \register[31][28] .power_up = "low";
// synopsys translate_on

// Location: FF_X60_Y35_N29
dffeas \register[19][28] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\register~67_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~39_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\register[19][28]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \register[19][28] .is_wysiwyg = "true";
defparam \register[19][28] .power_up = "low";
// synopsys translate_on

// Location: FF_X60_Y35_N7
dffeas \register[23][28] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\register~67_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~37_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\register[23][28]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \register[23][28] .is_wysiwyg = "true";
defparam \register[23][28] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X60_Y35_N6
cycloneive_lcell_comb \Mux35~7 (
// Equation(s):
// \Mux35~7_combout  = (Selector7 & (((Selector8)))) # (!Selector7 & ((Selector8 & ((\register[23][28]~q ))) # (!Selector8 & (\register[19][28]~q ))))

	.dataa(Selector7),
	.datab(\register[19][28]~q ),
	.datac(\register[23][28]~q ),
	.datad(Selector8),
	.cin(gnd),
	.combout(\Mux35~7_combout ),
	.cout());
// synopsys translate_off
defparam \Mux35~7 .lut_mask = 16'hFA44;
defparam \Mux35~7 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X67_Y35_N20
cycloneive_lcell_comb \Mux35~8 (
// Equation(s):
// \Mux35~8_combout  = (Selector7 & ((\Mux35~7_combout  & ((\register[31][28]~q ))) # (!\Mux35~7_combout  & (\register[27][28]~q )))) # (!Selector7 & (((\Mux35~7_combout ))))

	.dataa(\register[27][28]~q ),
	.datab(\register[31][28]~q ),
	.datac(Selector7),
	.datad(\Mux35~7_combout ),
	.cin(gnd),
	.combout(\Mux35~8_combout ),
	.cout());
// synopsys translate_off
defparam \Mux35~8 .lut_mask = 16'hCFA0;
defparam \Mux35~8 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X63_Y35_N14
cycloneive_lcell_comb \register[21][28]~feeder (
// Equation(s):
// \register[21][28]~feeder_combout  = \register~67_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(\register~67_combout ),
	.cin(gnd),
	.combout(\register[21][28]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \register[21][28]~feeder .lut_mask = 16'hFF00;
defparam \register[21][28]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X63_Y35_N15
dffeas \register[21][28] (
	.clk(!CLK),
	.d(\register[21][28]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~22_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\register[21][28]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \register[21][28] .is_wysiwyg = "true";
defparam \register[21][28] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X63_Y35_N28
cycloneive_lcell_comb \Mux35~0 (
// Equation(s):
// \Mux35~0_combout  = (Selector7 & (((Selector8)))) # (!Selector7 & ((Selector8 & ((\register[21][28]~q ))) # (!Selector8 & (\register[17][28]~q ))))

	.dataa(\register[17][28]~q ),
	.datab(\register[21][28]~q ),
	.datac(Selector7),
	.datad(Selector8),
	.cin(gnd),
	.combout(\Mux35~0_combout ),
	.cout());
// synopsys translate_off
defparam \Mux35~0 .lut_mask = 16'hFC0A;
defparam \Mux35~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X63_Y39_N6
cycloneive_lcell_comb \register[29][28]~feeder (
// Equation(s):
// \register[29][28]~feeder_combout  = \register~67_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(\register~67_combout ),
	.cin(gnd),
	.combout(\register[29][28]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \register[29][28]~feeder .lut_mask = 16'hFF00;
defparam \register[29][28]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X63_Y39_N7
dffeas \register[29][28] (
	.clk(!CLK),
	.d(\register[29][28]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~28_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\register[29][28]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \register[29][28] .is_wysiwyg = "true";
defparam \register[29][28] .power_up = "low";
// synopsys translate_on

// Location: FF_X63_Y37_N13
dffeas \register[25][28] (
	.clk(!CLK),
	.d(\register~67_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~24_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\register[25][28]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \register[25][28] .is_wysiwyg = "true";
defparam \register[25][28] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X67_Y35_N8
cycloneive_lcell_comb \Mux35~1 (
// Equation(s):
// \Mux35~1_combout  = (Selector7 & ((\Mux35~0_combout  & (\register[29][28]~q )) # (!\Mux35~0_combout  & ((\register[25][28]~q ))))) # (!Selector7 & (\Mux35~0_combout ))

	.dataa(Selector7),
	.datab(\Mux35~0_combout ),
	.datac(\register[29][28]~q ),
	.datad(\register[25][28]~q ),
	.cin(gnd),
	.combout(\Mux35~1_combout ),
	.cout());
// synopsys translate_off
defparam \Mux35~1 .lut_mask = 16'hE6C4;
defparam \Mux35~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X65_Y39_N11
dffeas \register[20][28] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\register~67_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~35_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\register[20][28]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \register[20][28] .is_wysiwyg = "true";
defparam \register[20][28] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X67_Y39_N24
cycloneive_lcell_comb \register[28][28]~feeder (
// Equation(s):
// \register[28][28]~feeder_combout  = \register~67_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(\register~67_combout ),
	.datad(gnd),
	.cin(gnd),
	.combout(\register[28][28]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \register[28][28]~feeder .lut_mask = 16'hF0F0;
defparam \register[28][28]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X67_Y39_N25
dffeas \register[28][28] (
	.clk(!CLK),
	.d(\register[28][28]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~57_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\register[28][28]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \register[28][28] .is_wysiwyg = "true";
defparam \register[28][28] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X67_Y35_N6
cycloneive_lcell_comb \Mux35~5 (
// Equation(s):
// \Mux35~5_combout  = (\Mux35~4_combout  & (((\register[28][28]~q ) # (!Selector8)))) # (!\Mux35~4_combout  & (\register[20][28]~q  & (Selector8)))

	.dataa(\Mux35~4_combout ),
	.datab(\register[20][28]~q ),
	.datac(Selector8),
	.datad(\register[28][28]~q ),
	.cin(gnd),
	.combout(\Mux35~5_combout ),
	.cout());
// synopsys translate_off
defparam \Mux35~5 .lut_mask = 16'hEA4A;
defparam \Mux35~5 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X69_Y39_N3
dffeas \register[18][28] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\register~67_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~33_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\register[18][28]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \register[18][28] .is_wysiwyg = "true";
defparam \register[18][28] .power_up = "low";
// synopsys translate_on

// Location: FF_X69_Y39_N13
dffeas \register[26][28] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\register~67_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~54_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\register[26][28]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \register[26][28] .is_wysiwyg = "true";
defparam \register[26][28] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X69_Y39_N12
cycloneive_lcell_comb \Mux35~2 (
// Equation(s):
// \Mux35~2_combout  = (Selector8 & (((Selector7)))) # (!Selector8 & ((Selector7 & ((\register[26][28]~q ))) # (!Selector7 & (\register[18][28]~q ))))

	.dataa(Selector8),
	.datab(\register[18][28]~q ),
	.datac(\register[26][28]~q ),
	.datad(Selector7),
	.cin(gnd),
	.combout(\Mux35~2_combout ),
	.cout());
// synopsys translate_off
defparam \Mux35~2 .lut_mask = 16'hFA44;
defparam \Mux35~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X69_Y35_N28
cycloneive_lcell_comb \register[22][28]~feeder (
// Equation(s):
// \register[22][28]~feeder_combout  = \register~67_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(\register~67_combout ),
	.cin(gnd),
	.combout(\register[22][28]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \register[22][28]~feeder .lut_mask = 16'hFF00;
defparam \register[22][28]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X69_Y35_N29
dffeas \register[22][28] (
	.clk(!CLK),
	.d(\register[22][28]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~55_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\register[22][28]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \register[22][28] .is_wysiwyg = "true";
defparam \register[22][28] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X67_Y39_N6
cycloneive_lcell_comb \Mux35~3 (
// Equation(s):
// \Mux35~3_combout  = (\Mux35~2_combout  & ((\register[30][28]~q ) # ((!Selector8)))) # (!\Mux35~2_combout  & (((Selector8 & \register[22][28]~q ))))

	.dataa(\register[30][28]~q ),
	.datab(\Mux35~2_combout ),
	.datac(Selector8),
	.datad(\register[22][28]~q ),
	.cin(gnd),
	.combout(\Mux35~3_combout ),
	.cout());
// synopsys translate_off
defparam \Mux35~3 .lut_mask = 16'hBC8C;
defparam \Mux35~3 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X67_Y35_N28
cycloneive_lcell_comb \Mux35~6 (
// Equation(s):
// \Mux35~6_combout  = (Selector10 & (((Selector91)))) # (!Selector10 & ((Selector91 & ((\Mux35~3_combout ))) # (!Selector91 & (\Mux35~5_combout ))))

	.dataa(\Mux35~5_combout ),
	.datab(Selector10),
	.datac(Selector91),
	.datad(\Mux35~3_combout ),
	.cin(gnd),
	.combout(\Mux35~6_combout ),
	.cout());
// synopsys translate_off
defparam \Mux35~6 .lut_mask = 16'hF2C2;
defparam \Mux35~6 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X63_Y37_N22
cycloneive_lcell_comb \register[15][28]~feeder (
// Equation(s):
// \register[15][28]~feeder_combout  = \register~67_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(\register~67_combout ),
	.cin(gnd),
	.combout(\register[15][28]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \register[15][28]~feeder .lut_mask = 16'hFF00;
defparam \register[15][28]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X63_Y37_N23
dffeas \register[15][28] (
	.clk(!CLK),
	.d(\register[15][28]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~53_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\register[15][28]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \register[15][28] .is_wysiwyg = "true";
defparam \register[15][28] .power_up = "low";
// synopsys translate_on

// Location: FF_X60_Y36_N1
dffeas \register[14][28] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\register~67_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~61_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\register[14][28]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \register[14][28] .is_wysiwyg = "true";
defparam \register[14][28] .power_up = "low";
// synopsys translate_on

// Location: FF_X60_Y36_N19
dffeas \register[12][28] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\register~67_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~52_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\register[12][28]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \register[12][28] .is_wysiwyg = "true";
defparam \register[12][28] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X60_Y36_N18
cycloneive_lcell_comb \Mux35~17 (
// Equation(s):
// \Mux35~17_combout  = (Selector10 & ((\register[13][28]~q ) # ((Selector91)))) # (!Selector10 & (((\register[12][28]~q  & !Selector91))))

	.dataa(\register[13][28]~q ),
	.datab(Selector10),
	.datac(\register[12][28]~q ),
	.datad(Selector91),
	.cin(gnd),
	.combout(\Mux35~17_combout ),
	.cout());
// synopsys translate_off
defparam \Mux35~17 .lut_mask = 16'hCCB8;
defparam \Mux35~17 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y36_N0
cycloneive_lcell_comb \Mux35~18 (
// Equation(s):
// \Mux35~18_combout  = (Selector91 & ((\Mux35~17_combout  & (\register[15][28]~q )) # (!\Mux35~17_combout  & ((\register[14][28]~q ))))) # (!Selector91 & (((\Mux35~17_combout ))))

	.dataa(Selector91),
	.datab(\register[15][28]~q ),
	.datac(\register[14][28]~q ),
	.datad(\Mux35~17_combout ),
	.cin(gnd),
	.combout(\Mux35~18_combout ),
	.cout());
// synopsys translate_off
defparam \Mux35~18 .lut_mask = 16'hDDA0;
defparam \Mux35~18 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X66_Y32_N8
cycloneive_lcell_comb \register[2][28]~feeder (
// Equation(s):
// \register[2][28]~feeder_combout  = \register~67_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(\register~67_combout ),
	.datad(gnd),
	.cin(gnd),
	.combout(\register[2][28]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \register[2][28]~feeder .lut_mask = 16'hF0F0;
defparam \register[2][28]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X66_Y32_N9
dffeas \register[2][28] (
	.clk(!CLK),
	.d(\register[2][28]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~50_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\register[2][28]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \register[2][28] .is_wysiwyg = "true";
defparam \register[2][28] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X66_Y32_N2
cycloneive_lcell_comb \Mux35~15 (
// Equation(s):
// \Mux35~15_combout  = (\Mux35~14_combout ) # ((\register[2][28]~q  & (Selector91 & !Selector10)))

	.dataa(\Mux35~14_combout ),
	.datab(\register[2][28]~q ),
	.datac(Selector91),
	.datad(Selector10),
	.cin(gnd),
	.combout(\Mux35~15_combout ),
	.cout());
// synopsys translate_off
defparam \Mux35~15 .lut_mask = 16'hAAEA;
defparam \Mux35~15 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X66_Y32_N28
cycloneive_lcell_comb \register[7][28]~feeder (
// Equation(s):
// \register[7][28]~feeder_combout  = \register~67_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(\register~67_combout ),
	.datad(gnd),
	.cin(gnd),
	.combout(\register[7][28]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \register[7][28]~feeder .lut_mask = 16'hF0F0;
defparam \register[7][28]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X66_Y32_N29
dffeas \register[7][28] (
	.clk(!CLK),
	.d(\register[7][28]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~43_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\register[7][28]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \register[7][28] .is_wysiwyg = "true";
defparam \register[7][28] .power_up = "low";
// synopsys translate_on

// Location: FF_X69_Y31_N21
dffeas \register[5][28] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\register~67_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~59_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\register[5][28]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \register[5][28] .is_wysiwyg = "true";
defparam \register[5][28] .power_up = "low";
// synopsys translate_on

// Location: FF_X69_Y31_N19
dffeas \register[4][28] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\register~67_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~60_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\register[4][28]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \register[4][28] .is_wysiwyg = "true";
defparam \register[4][28] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X69_Y31_N18
cycloneive_lcell_comb \Mux35~12 (
// Equation(s):
// \Mux35~12_combout  = (Selector10 & ((\register[5][28]~q ) # ((Selector91)))) # (!Selector10 & (((\register[4][28]~q  & !Selector91))))

	.dataa(Selector10),
	.datab(\register[5][28]~q ),
	.datac(\register[4][28]~q ),
	.datad(Selector91),
	.cin(gnd),
	.combout(\Mux35~12_combout ),
	.cout());
// synopsys translate_off
defparam \Mux35~12 .lut_mask = 16'hAAD8;
defparam \Mux35~12 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X66_Y32_N14
cycloneive_lcell_comb \Mux35~13 (
// Equation(s):
// \Mux35~13_combout  = (Selector91 & ((\Mux35~12_combout  & ((\register[7][28]~q ))) # (!\Mux35~12_combout  & (\register[6][28]~q )))) # (!Selector91 & (((\Mux35~12_combout ))))

	.dataa(\register[6][28]~q ),
	.datab(\register[7][28]~q ),
	.datac(Selector91),
	.datad(\Mux35~12_combout ),
	.cin(gnd),
	.combout(\Mux35~13_combout ),
	.cout());
// synopsys translate_off
defparam \Mux35~13 .lut_mask = 16'hCFA0;
defparam \Mux35~13 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X67_Y35_N4
cycloneive_lcell_comb \Mux35~16 (
// Equation(s):
// \Mux35~16_combout  = (Selector8 & ((Selector7) # ((\Mux35~13_combout )))) # (!Selector8 & (!Selector7 & (\Mux35~15_combout )))

	.dataa(Selector8),
	.datab(Selector7),
	.datac(\Mux35~15_combout ),
	.datad(\Mux35~13_combout ),
	.cin(gnd),
	.combout(\Mux35~16_combout ),
	.cout());
// synopsys translate_off
defparam \Mux35~16 .lut_mask = 16'hBA98;
defparam \Mux35~16 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X65_Y40_N19
dffeas \register[11][28] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\register~67_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~47_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\register[11][28]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \register[11][28] .is_wysiwyg = "true";
defparam \register[11][28] .power_up = "low";
// synopsys translate_on

// Location: FF_X65_Y40_N9
dffeas \register[9][28] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\register~67_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~44_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\register[9][28]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \register[9][28] .is_wysiwyg = "true";
defparam \register[9][28] .power_up = "low";
// synopsys translate_on

// Location: FF_X62_Y41_N3
dffeas \register[8][28] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\register~67_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~46_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\register[8][28]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \register[8][28] .is_wysiwyg = "true";
defparam \register[8][28] .power_up = "low";
// synopsys translate_on

// Location: FF_X62_Y41_N5
dffeas \register[10][28] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\register~67_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~45_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\register[10][28]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \register[10][28] .is_wysiwyg = "true";
defparam \register[10][28] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X62_Y41_N4
cycloneive_lcell_comb \Mux35~10 (
// Equation(s):
// \Mux35~10_combout  = (Selector10 & (((Selector91)))) # (!Selector10 & ((Selector91 & ((\register[10][28]~q ))) # (!Selector91 & (\register[8][28]~q ))))

	.dataa(Selector10),
	.datab(\register[8][28]~q ),
	.datac(\register[10][28]~q ),
	.datad(Selector91),
	.cin(gnd),
	.combout(\Mux35~10_combout ),
	.cout());
// synopsys translate_off
defparam \Mux35~10 .lut_mask = 16'hFA44;
defparam \Mux35~10 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X65_Y40_N8
cycloneive_lcell_comb \Mux35~11 (
// Equation(s):
// \Mux35~11_combout  = (Selector10 & ((\Mux35~10_combout  & (\register[11][28]~q )) # (!\Mux35~10_combout  & ((\register[9][28]~q ))))) # (!Selector10 & (((\Mux35~10_combout ))))

	.dataa(Selector10),
	.datab(\register[11][28]~q ),
	.datac(\register[9][28]~q ),
	.datad(\Mux35~10_combout ),
	.cin(gnd),
	.combout(\Mux35~11_combout ),
	.cout());
// synopsys translate_off
defparam \Mux35~11 .lut_mask = 16'hDDA0;
defparam \Mux35~11 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y35_N0
cycloneive_lcell_comb \register~68 (
// Equation(s):
// \register~68_combout  = (WideOr01 & ((\wdat[27]~8_combout ) # ((plif_memwbrtnaddr_l_27 & plif_memwbregsrc_l_1))))

	.dataa(plif_memwbrtnaddr_l_27),
	.datab(plif_memwbregsrc_l_1),
	.datac(WideOr0),
	.datad(wdat_27),
	.cin(gnd),
	.combout(\register~68_combout ),
	.cout());
// synopsys translate_off
defparam \register~68 .lut_mask = 16'hF080;
defparam \register~68 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y39_N18
cycloneive_lcell_comb \register[23][27]~feeder (
// Equation(s):
// \register[23][27]~feeder_combout  = \register~68_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(\register~68_combout ),
	.datad(gnd),
	.cin(gnd),
	.combout(\register[23][27]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \register[23][27]~feeder .lut_mask = 16'hF0F0;
defparam \register[23][27]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X61_Y39_N19
dffeas \register[23][27] (
	.clk(!CLK),
	.d(\register[23][27]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~37_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\register[23][27]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \register[23][27] .is_wysiwyg = "true";
defparam \register[23][27] .power_up = "low";
// synopsys translate_on

// Location: FF_X62_Y39_N1
dffeas \register[31][27] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\register~68_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~40_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\register[31][27]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \register[31][27] .is_wysiwyg = "true";
defparam \register[31][27] .power_up = "low";
// synopsys translate_on

// Location: FF_X62_Y39_N19
dffeas \register[27][27] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\register~68_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~38_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\register[27][27]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \register[27][27] .is_wysiwyg = "true";
defparam \register[27][27] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X62_Y39_N18
cycloneive_lcell_comb \Mux36~7 (
// Equation(s):
// \Mux36~7_combout  = (Selector8 & (((Selector7)))) # (!Selector8 & ((Selector7 & ((\register[27][27]~q ))) # (!Selector7 & (\register[19][27]~q ))))

	.dataa(\register[19][27]~q ),
	.datab(Selector8),
	.datac(\register[27][27]~q ),
	.datad(Selector7),
	.cin(gnd),
	.combout(\Mux36~7_combout ),
	.cout());
// synopsys translate_off
defparam \Mux36~7 .lut_mask = 16'hFC22;
defparam \Mux36~7 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y39_N12
cycloneive_lcell_comb \Mux36~8 (
// Equation(s):
// \Mux36~8_combout  = (Selector8 & ((\Mux36~7_combout  & ((\register[31][27]~q ))) # (!\Mux36~7_combout  & (\register[23][27]~q )))) # (!Selector8 & (((\Mux36~7_combout ))))

	.dataa(Selector8),
	.datab(\register[23][27]~q ),
	.datac(\register[31][27]~q ),
	.datad(\Mux36~7_combout ),
	.cin(gnd),
	.combout(\Mux36~8_combout ),
	.cout());
// synopsys translate_off
defparam \Mux36~8 .lut_mask = 16'hF588;
defparam \Mux36~8 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X63_Y39_N16
cycloneive_lcell_comb \register[29][27]~feeder (
// Equation(s):
// \register[29][27]~feeder_combout  = \register~68_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(\register~68_combout ),
	.cin(gnd),
	.combout(\register[29][27]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \register[29][27]~feeder .lut_mask = 16'hFF00;
defparam \register[29][27]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X63_Y39_N17
dffeas \register[29][27] (
	.clk(!CLK),
	.d(\register[29][27]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~28_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\register[29][27]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \register[29][27] .is_wysiwyg = "true";
defparam \register[29][27] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X62_Y35_N6
cycloneive_lcell_comb \register[17][27]~feeder (
// Equation(s):
// \register[17][27]~feeder_combout  = \register~68_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(\register~68_combout ),
	.cin(gnd),
	.combout(\register[17][27]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \register[17][27]~feeder .lut_mask = 16'hFF00;
defparam \register[17][27]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X62_Y35_N7
dffeas \register[17][27] (
	.clk(!CLK),
	.d(\register[17][27]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~26_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\register[17][27]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \register[17][27] .is_wysiwyg = "true";
defparam \register[17][27] .power_up = "low";
// synopsys translate_on

// Location: FF_X61_Y37_N5
dffeas \register[25][27] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\register~68_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~24_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\register[25][27]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \register[25][27] .is_wysiwyg = "true";
defparam \register[25][27] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X61_Y37_N4
cycloneive_lcell_comb \Mux36~0 (
// Equation(s):
// \Mux36~0_combout  = (Selector8 & (((Selector7)))) # (!Selector8 & ((Selector7 & ((\register[25][27]~q ))) # (!Selector7 & (\register[17][27]~q ))))

	.dataa(Selector8),
	.datab(\register[17][27]~q ),
	.datac(\register[25][27]~q ),
	.datad(Selector7),
	.cin(gnd),
	.combout(\Mux36~0_combout ),
	.cout());
// synopsys translate_off
defparam \Mux36~0 .lut_mask = 16'hFA44;
defparam \Mux36~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X61_Y35_N1
dffeas \register[21][27] (
	.clk(!CLK),
	.d(\register~68_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~22_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\register[21][27]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \register[21][27] .is_wysiwyg = "true";
defparam \register[21][27] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X61_Y39_N22
cycloneive_lcell_comb \Mux36~1 (
// Equation(s):
// \Mux36~1_combout  = (Selector8 & ((\Mux36~0_combout  & (\register[29][27]~q )) # (!\Mux36~0_combout  & ((\register[21][27]~q ))))) # (!Selector8 & (((\Mux36~0_combout ))))

	.dataa(Selector8),
	.datab(\register[29][27]~q ),
	.datac(\Mux36~0_combout ),
	.datad(\register[21][27]~q ),
	.cin(gnd),
	.combout(\Mux36~1_combout ),
	.cout());
// synopsys translate_off
defparam \Mux36~1 .lut_mask = 16'hDAD0;
defparam \Mux36~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X65_Y39_N25
dffeas \register[16][27] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\register~68_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~36_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\register[16][27]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \register[16][27] .is_wysiwyg = "true";
defparam \register[16][27] .power_up = "low";
// synopsys translate_on

// Location: FF_X65_Y39_N27
dffeas \register[20][27] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\register~68_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~35_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\register[20][27]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \register[20][27] .is_wysiwyg = "true";
defparam \register[20][27] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X65_Y39_N26
cycloneive_lcell_comb \Mux36~4 (
// Equation(s):
// \Mux36~4_combout  = (Selector7 & (((Selector8)))) # (!Selector7 & ((Selector8 & ((\register[20][27]~q ))) # (!Selector8 & (\register[16][27]~q ))))

	.dataa(Selector7),
	.datab(\register[16][27]~q ),
	.datac(\register[20][27]~q ),
	.datad(Selector8),
	.cin(gnd),
	.combout(\Mux36~4_combout ),
	.cout());
// synopsys translate_off
defparam \Mux36~4 .lut_mask = 16'hFA44;
defparam \Mux36~4 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X61_Y37_N23
dffeas \register[24][27] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\register~68_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~34_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\register[24][27]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \register[24][27] .is_wysiwyg = "true";
defparam \register[24][27] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X66_Y39_N28
cycloneive_lcell_comb \register[28][27]~feeder (
// Equation(s):
// \register[28][27]~feeder_combout  = \register~68_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(\register~68_combout ),
	.cin(gnd),
	.combout(\register[28][27]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \register[28][27]~feeder .lut_mask = 16'hFF00;
defparam \register[28][27]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X66_Y39_N29
dffeas \register[28][27] (
	.clk(!CLK),
	.d(\register[28][27]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~57_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\register[28][27]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \register[28][27] .is_wysiwyg = "true";
defparam \register[28][27] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X61_Y37_N22
cycloneive_lcell_comb \Mux36~5 (
// Equation(s):
// \Mux36~5_combout  = (Selector7 & ((\Mux36~4_combout  & ((\register[28][27]~q ))) # (!\Mux36~4_combout  & (\register[24][27]~q )))) # (!Selector7 & (\Mux36~4_combout ))

	.dataa(Selector7),
	.datab(\Mux36~4_combout ),
	.datac(\register[24][27]~q ),
	.datad(\register[28][27]~q ),
	.cin(gnd),
	.combout(\Mux36~5_combout ),
	.cout());
// synopsys translate_off
defparam \Mux36~5 .lut_mask = 16'hEC64;
defparam \Mux36~5 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X68_Y35_N19
dffeas \register[30][27] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\register~68_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~56_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\register[30][27]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \register[30][27] .is_wysiwyg = "true";
defparam \register[30][27] .power_up = "low";
// synopsys translate_on

// Location: FF_X67_Y37_N5
dffeas \register[22][27] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\register~68_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~55_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\register[22][27]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \register[22][27] .is_wysiwyg = "true";
defparam \register[22][27] .power_up = "low";
// synopsys translate_on

// Location: FF_X67_Y37_N15
dffeas \register[18][27] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\register~68_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~33_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\register[18][27]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \register[18][27] .is_wysiwyg = "true";
defparam \register[18][27] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X67_Y37_N14
cycloneive_lcell_comb \Mux36~2 (
// Equation(s):
// \Mux36~2_combout  = (Selector8 & ((\register[22][27]~q ) # ((Selector7)))) # (!Selector8 & (((\register[18][27]~q  & !Selector7))))

	.dataa(Selector8),
	.datab(\register[22][27]~q ),
	.datac(\register[18][27]~q ),
	.datad(Selector7),
	.cin(gnd),
	.combout(\Mux36~2_combout ),
	.cout());
// synopsys translate_off
defparam \Mux36~2 .lut_mask = 16'hAAD8;
defparam \Mux36~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X68_Y35_N1
dffeas \register[26][27] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\register~68_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~54_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\register[26][27]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \register[26][27] .is_wysiwyg = "true";
defparam \register[26][27] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X68_Y35_N24
cycloneive_lcell_comb \Mux36~3 (
// Equation(s):
// \Mux36~3_combout  = (Selector7 & ((\Mux36~2_combout  & (\register[30][27]~q )) # (!\Mux36~2_combout  & ((\register[26][27]~q ))))) # (!Selector7 & (((\Mux36~2_combout ))))

	.dataa(Selector7),
	.datab(\register[30][27]~q ),
	.datac(\Mux36~2_combout ),
	.datad(\register[26][27]~q ),
	.cin(gnd),
	.combout(\Mux36~3_combout ),
	.cout());
// synopsys translate_off
defparam \Mux36~3 .lut_mask = 16'hDAD0;
defparam \Mux36~3 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y39_N28
cycloneive_lcell_comb \Mux36~6 (
// Equation(s):
// \Mux36~6_combout  = (Selector10 & (Selector91)) # (!Selector10 & ((Selector91 & ((\Mux36~3_combout ))) # (!Selector91 & (\Mux36~5_combout ))))

	.dataa(Selector10),
	.datab(Selector91),
	.datac(\Mux36~5_combout ),
	.datad(\Mux36~3_combout ),
	.cin(gnd),
	.combout(\Mux36~6_combout ),
	.cout());
// synopsys translate_off
defparam \Mux36~6 .lut_mask = 16'hDC98;
defparam \Mux36~6 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X69_Y31_N9
dffeas \register[5][27] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\register~68_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~59_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\register[5][27]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \register[5][27] .is_wysiwyg = "true";
defparam \register[5][27] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X69_Y31_N8
cycloneive_lcell_comb \Mux36~10 (
// Equation(s):
// \Mux36~10_combout  = (Selector91 & (((Selector10)))) # (!Selector91 & ((Selector10 & ((\register[5][27]~q ))) # (!Selector10 & (\register[4][27]~q ))))

	.dataa(\register[4][27]~q ),
	.datab(Selector91),
	.datac(\register[5][27]~q ),
	.datad(Selector10),
	.cin(gnd),
	.combout(\Mux36~10_combout ),
	.cout());
// synopsys translate_off
defparam \Mux36~10 .lut_mask = 16'hFC22;
defparam \Mux36~10 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X68_Y31_N29
dffeas \register[6][27] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\register~68_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~58_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\register[6][27]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \register[6][27] .is_wysiwyg = "true";
defparam \register[6][27] .power_up = "low";
// synopsys translate_on

// Location: FF_X68_Y31_N3
dffeas \register[7][27] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\register~68_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~43_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\register[7][27]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \register[7][27] .is_wysiwyg = "true";
defparam \register[7][27] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X68_Y31_N28
cycloneive_lcell_comb \Mux36~11 (
// Equation(s):
// \Mux36~11_combout  = (Selector91 & ((\Mux36~10_combout  & ((\register[7][27]~q ))) # (!\Mux36~10_combout  & (\register[6][27]~q )))) # (!Selector91 & (\Mux36~10_combout ))

	.dataa(Selector91),
	.datab(\Mux36~10_combout ),
	.datac(\register[6][27]~q ),
	.datad(\register[7][27]~q ),
	.cin(gnd),
	.combout(\Mux36~11_combout ),
	.cout());
// synopsys translate_off
defparam \Mux36~11 .lut_mask = 16'hEC64;
defparam \Mux36~11 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y35_N18
cycloneive_lcell_comb \register[15][27]~feeder (
// Equation(s):
// \register[15][27]~feeder_combout  = \register~68_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(\register~68_combout ),
	.cin(gnd),
	.combout(\register[15][27]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \register[15][27]~feeder .lut_mask = 16'hFF00;
defparam \register[15][27]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X61_Y35_N19
dffeas \register[15][27] (
	.clk(!CLK),
	.d(\register[15][27]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~53_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\register[15][27]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \register[15][27] .is_wysiwyg = "true";
defparam \register[15][27] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X62_Y32_N8
cycloneive_lcell_comb \register[14][27]~feeder (
// Equation(s):
// \register[14][27]~feeder_combout  = \register~68_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(\register~68_combout ),
	.cin(gnd),
	.combout(\register[14][27]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \register[14][27]~feeder .lut_mask = 16'hFF00;
defparam \register[14][27]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X62_Y32_N9
dffeas \register[14][27] (
	.clk(!CLK),
	.d(\register[14][27]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~61_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\register[14][27]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \register[14][27] .is_wysiwyg = "true";
defparam \register[14][27] .power_up = "low";
// synopsys translate_on

// Location: FF_X62_Y30_N13
dffeas \register[13][27] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\register~68_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~62_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\register[13][27]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \register[13][27] .is_wysiwyg = "true";
defparam \register[13][27] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X62_Y30_N12
cycloneive_lcell_comb \Mux36~17 (
// Equation(s):
// \Mux36~17_combout  = (Selector91 & (((Selector10)))) # (!Selector91 & ((Selector10 & ((\register[13][27]~q ))) # (!Selector10 & (\register[12][27]~q ))))

	.dataa(\register[12][27]~q ),
	.datab(Selector91),
	.datac(\register[13][27]~q ),
	.datad(Selector10),
	.cin(gnd),
	.combout(\Mux36~17_combout ),
	.cout());
// synopsys translate_off
defparam \Mux36~17 .lut_mask = 16'hFC22;
defparam \Mux36~17 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y35_N16
cycloneive_lcell_comb \Mux36~18 (
// Equation(s):
// \Mux36~18_combout  = (\Mux36~17_combout  & ((\register[15][27]~q ) # ((!Selector91)))) # (!\Mux36~17_combout  & (((\register[14][27]~q  & Selector91))))

	.dataa(\register[15][27]~q ),
	.datab(\register[14][27]~q ),
	.datac(\Mux36~17_combout ),
	.datad(Selector91),
	.cin(gnd),
	.combout(\Mux36~18_combout ),
	.cout());
// synopsys translate_off
defparam \Mux36~18 .lut_mask = 16'hACF0;
defparam \Mux36~18 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X69_Y33_N27
dffeas \register[1][27] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\register~68_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~49_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\register[1][27]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \register[1][27] .is_wysiwyg = "true";
defparam \register[1][27] .power_up = "low";
// synopsys translate_on

// Location: FF_X69_Y33_N1
dffeas \register[3][27] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\register~68_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~48_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\register[3][27]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \register[3][27] .is_wysiwyg = "true";
defparam \register[3][27] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X69_Y33_N26
cycloneive_lcell_comb \Mux36~14 (
// Equation(s):
// \Mux36~14_combout  = (Selector9 & ((plif_ifidinstr_l_17 & ((\register[3][27]~q ))) # (!plif_ifidinstr_l_17 & (\register[1][27]~q )))) # (!Selector9 & (((\register[1][27]~q ))))

	.dataa(Selector9),
	.datab(plif_ifidinstr_l_17),
	.datac(\register[1][27]~q ),
	.datad(\register[3][27]~q ),
	.cin(gnd),
	.combout(\Mux36~14_combout ),
	.cout());
// synopsys translate_off
defparam \Mux36~14 .lut_mask = 16'hF870;
defparam \Mux36~14 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y39_N24
cycloneive_lcell_comb \Mux36~15 (
// Equation(s):
// \Mux36~15_combout  = (Selector10 & (((\Mux36~14_combout )))) # (!Selector10 & (\register[2][27]~q  & (Selector91)))

	.dataa(\register[2][27]~q ),
	.datab(Selector10),
	.datac(Selector91),
	.datad(\Mux36~14_combout ),
	.cin(gnd),
	.combout(\Mux36~15_combout ),
	.cout());
// synopsys translate_off
defparam \Mux36~15 .lut_mask = 16'hEC20;
defparam \Mux36~15 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X66_Y38_N23
dffeas \register[9][27] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\register~68_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~44_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\register[9][27]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \register[9][27] .is_wysiwyg = "true";
defparam \register[9][27] .power_up = "low";
// synopsys translate_on

// Location: FF_X67_Y34_N23
dffeas \register[11][27] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\register~68_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~47_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\register[11][27]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \register[11][27] .is_wysiwyg = "true";
defparam \register[11][27] .power_up = "low";
// synopsys translate_on

// Location: FF_X62_Y41_N1
dffeas \register[10][27] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\register~68_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~45_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\register[10][27]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \register[10][27] .is_wysiwyg = "true";
defparam \register[10][27] .power_up = "low";
// synopsys translate_on

// Location: FF_X62_Y41_N11
dffeas \register[8][27] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\register~68_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~46_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\register[8][27]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \register[8][27] .is_wysiwyg = "true";
defparam \register[8][27] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X62_Y41_N0
cycloneive_lcell_comb \Mux36~12 (
// Equation(s):
// \Mux36~12_combout  = (Selector10 & (Selector91)) # (!Selector10 & ((Selector91 & (\register[10][27]~q )) # (!Selector91 & ((\register[8][27]~q )))))

	.dataa(Selector10),
	.datab(Selector91),
	.datac(\register[10][27]~q ),
	.datad(\register[8][27]~q ),
	.cin(gnd),
	.combout(\Mux36~12_combout ),
	.cout());
// synopsys translate_off
defparam \Mux36~12 .lut_mask = 16'hD9C8;
defparam \Mux36~12 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X67_Y34_N22
cycloneive_lcell_comb \Mux36~13 (
// Equation(s):
// \Mux36~13_combout  = (Selector10 & ((\Mux36~12_combout  & ((\register[11][27]~q ))) # (!\Mux36~12_combout  & (\register[9][27]~q )))) # (!Selector10 & (((\Mux36~12_combout ))))

	.dataa(Selector10),
	.datab(\register[9][27]~q ),
	.datac(\register[11][27]~q ),
	.datad(\Mux36~12_combout ),
	.cin(gnd),
	.combout(\Mux36~13_combout ),
	.cout());
// synopsys translate_off
defparam \Mux36~13 .lut_mask = 16'hF588;
defparam \Mux36~13 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y39_N10
cycloneive_lcell_comb \Mux36~16 (
// Equation(s):
// \Mux36~16_combout  = (Selector7 & (((Selector8) # (\Mux36~13_combout )))) # (!Selector7 & (\Mux36~15_combout  & (!Selector8)))

	.dataa(Selector7),
	.datab(\Mux36~15_combout ),
	.datac(Selector8),
	.datad(\Mux36~13_combout ),
	.cin(gnd),
	.combout(\Mux36~16_combout ),
	.cout());
// synopsys translate_off
defparam \Mux36~16 .lut_mask = 16'hAEA4;
defparam \Mux36~16 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X63_Y37_N10
cycloneive_lcell_comb \register~69 (
// Equation(s):
// \register~69_combout  = (WideOr01 & ((\wdat[26]~10_combout ) # ((plif_memwbregsrc_l_1 & plif_memwbrtnaddr_l_26))))

	.dataa(plif_memwbregsrc_l_1),
	.datab(plif_memwbrtnaddr_l_26),
	.datac(WideOr0),
	.datad(wdat_26),
	.cin(gnd),
	.combout(\register~69_combout ),
	.cout());
// synopsys translate_off
defparam \register~69 .lut_mask = 16'hF080;
defparam \register~69 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X60_Y37_N25
dffeas \register[17][26] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\register~69_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~26_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\register[17][26]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \register[17][26] .is_wysiwyg = "true";
defparam \register[17][26] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X63_Y35_N18
cycloneive_lcell_comb \register[21][26]~feeder (
// Equation(s):
// \register[21][26]~feeder_combout  = \register~69_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(\register~69_combout ),
	.datad(gnd),
	.cin(gnd),
	.combout(\register[21][26]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \register[21][26]~feeder .lut_mask = 16'hF0F0;
defparam \register[21][26]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X63_Y35_N19
dffeas \register[21][26] (
	.clk(!CLK),
	.d(\register[21][26]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~22_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\register[21][26]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \register[21][26] .is_wysiwyg = "true";
defparam \register[21][26] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X63_Y35_N4
cycloneive_lcell_comb \Mux37~0 (
// Equation(s):
// \Mux37~0_combout  = (Selector7 & (Selector8)) # (!Selector7 & ((Selector8 & ((\register[21][26]~q ))) # (!Selector8 & (\register[17][26]~q ))))

	.dataa(Selector7),
	.datab(Selector8),
	.datac(\register[17][26]~q ),
	.datad(\register[21][26]~q ),
	.cin(gnd),
	.combout(\Mux37~0_combout ),
	.cout());
// synopsys translate_off
defparam \Mux37~0 .lut_mask = 16'hDC98;
defparam \Mux37~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X61_Y32_N21
dffeas \register[29][26] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\register~69_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~28_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\register[29][26]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \register[29][26] .is_wysiwyg = "true";
defparam \register[29][26] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X63_Y37_N16
cycloneive_lcell_comb \register[25][26]~feeder (
// Equation(s):
// \register[25][26]~feeder_combout  = \register~69_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(\register~69_combout ),
	.cin(gnd),
	.combout(\register[25][26]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \register[25][26]~feeder .lut_mask = 16'hFF00;
defparam \register[25][26]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X63_Y37_N17
dffeas \register[25][26] (
	.clk(!CLK),
	.d(\register[25][26]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~24_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\register[25][26]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \register[25][26] .is_wysiwyg = "true";
defparam \register[25][26] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X61_Y32_N20
cycloneive_lcell_comb \Mux37~1 (
// Equation(s):
// \Mux37~1_combout  = (\Mux37~0_combout  & (((\register[29][26]~q )) # (!Selector7))) # (!\Mux37~0_combout  & (Selector7 & ((\register[25][26]~q ))))

	.dataa(\Mux37~0_combout ),
	.datab(Selector7),
	.datac(\register[29][26]~q ),
	.datad(\register[25][26]~q ),
	.cin(gnd),
	.combout(\Mux37~1_combout ),
	.cout());
// synopsys translate_off
defparam \Mux37~1 .lut_mask = 16'hE6A2;
defparam \Mux37~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X60_Y35_N5
dffeas \register[19][26] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\register~69_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~39_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\register[19][26]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \register[19][26] .is_wysiwyg = "true";
defparam \register[19][26] .power_up = "low";
// synopsys translate_on

// Location: FF_X60_Y35_N15
dffeas \register[23][26] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\register~69_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~37_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\register[23][26]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \register[23][26] .is_wysiwyg = "true";
defparam \register[23][26] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X60_Y35_N14
cycloneive_lcell_comb \Mux37~7 (
// Equation(s):
// \Mux37~7_combout  = (Selector7 & (((Selector8)))) # (!Selector7 & ((Selector8 & ((\register[23][26]~q ))) # (!Selector8 & (\register[19][26]~q ))))

	.dataa(Selector7),
	.datab(\register[19][26]~q ),
	.datac(\register[23][26]~q ),
	.datad(Selector8),
	.cin(gnd),
	.combout(\Mux37~7_combout ),
	.cout());
// synopsys translate_off
defparam \Mux37~7 .lut_mask = 16'hFA44;
defparam \Mux37~7 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X63_Y35_N2
cycloneive_lcell_comb \register[27][26]~feeder (
// Equation(s):
// \register[27][26]~feeder_combout  = \register~69_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(\register~69_combout ),
	.datad(gnd),
	.cin(gnd),
	.combout(\register[27][26]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \register[27][26]~feeder .lut_mask = 16'hF0F0;
defparam \register[27][26]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X63_Y35_N3
dffeas \register[27][26] (
	.clk(!CLK),
	.d(\register[27][26]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~38_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\register[27][26]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \register[27][26] .is_wysiwyg = "true";
defparam \register[27][26] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X63_Y32_N2
cycloneive_lcell_comb \register[31][26]~feeder (
// Equation(s):
// \register[31][26]~feeder_combout  = \register~69_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(\register~69_combout ),
	.cin(gnd),
	.combout(\register[31][26]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \register[31][26]~feeder .lut_mask = 16'hFF00;
defparam \register[31][26]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X63_Y32_N3
dffeas \register[31][26] (
	.clk(!CLK),
	.d(\register[31][26]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~40_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\register[31][26]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \register[31][26] .is_wysiwyg = "true";
defparam \register[31][26] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X63_Y35_N8
cycloneive_lcell_comb \Mux37~8 (
// Equation(s):
// \Mux37~8_combout  = (\Mux37~7_combout  & (((\register[31][26]~q ) # (!Selector7)))) # (!\Mux37~7_combout  & (\register[27][26]~q  & (Selector7)))

	.dataa(\Mux37~7_combout ),
	.datab(\register[27][26]~q ),
	.datac(Selector7),
	.datad(\register[31][26]~q ),
	.cin(gnd),
	.combout(\Mux37~8_combout ),
	.cout());
// synopsys translate_off
defparam \Mux37~8 .lut_mask = 16'hEA4A;
defparam \Mux37~8 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X68_Y34_N16
cycloneive_lcell_comb \register[30][26]~feeder (
// Equation(s):
// \register[30][26]~feeder_combout  = \register~69_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(\register~69_combout ),
	.cin(gnd),
	.combout(\register[30][26]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \register[30][26]~feeder .lut_mask = 16'hFF00;
defparam \register[30][26]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X68_Y34_N17
dffeas \register[30][26] (
	.clk(!CLK),
	.d(\register[30][26]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~56_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\register[30][26]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \register[30][26] .is_wysiwyg = "true";
defparam \register[30][26] .power_up = "low";
// synopsys translate_on

// Location: FF_X69_Y35_N15
dffeas \register[22][26] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\register~69_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~55_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\register[22][26]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \register[22][26] .is_wysiwyg = "true";
defparam \register[22][26] .power_up = "low";
// synopsys translate_on

// Location: FF_X69_Y35_N17
dffeas \register[18][26] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\register~69_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~33_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\register[18][26]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \register[18][26] .is_wysiwyg = "true";
defparam \register[18][26] .power_up = "low";
// synopsys translate_on

// Location: FF_X69_Y39_N25
dffeas \register[26][26] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\register~69_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~54_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\register[26][26]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \register[26][26] .is_wysiwyg = "true";
defparam \register[26][26] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X69_Y39_N24
cycloneive_lcell_comb \Mux37~2 (
// Equation(s):
// \Mux37~2_combout  = (Selector8 & (((Selector7)))) # (!Selector8 & ((Selector7 & ((\register[26][26]~q ))) # (!Selector7 & (\register[18][26]~q ))))

	.dataa(Selector8),
	.datab(\register[18][26]~q ),
	.datac(\register[26][26]~q ),
	.datad(Selector7),
	.cin(gnd),
	.combout(\Mux37~2_combout ),
	.cout());
// synopsys translate_off
defparam \Mux37~2 .lut_mask = 16'hFA44;
defparam \Mux37~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X69_Y35_N14
cycloneive_lcell_comb \Mux37~3 (
// Equation(s):
// \Mux37~3_combout  = (Selector8 & ((\Mux37~2_combout  & (\register[30][26]~q )) # (!\Mux37~2_combout  & ((\register[22][26]~q ))))) # (!Selector8 & (((\Mux37~2_combout ))))

	.dataa(Selector8),
	.datab(\register[30][26]~q ),
	.datac(\register[22][26]~q ),
	.datad(\Mux37~2_combout ),
	.cin(gnd),
	.combout(\Mux37~3_combout ),
	.cout());
// synopsys translate_off
defparam \Mux37~3 .lut_mask = 16'hDDA0;
defparam \Mux37~3 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X66_Y35_N10
cycloneive_lcell_comb \register[28][26]~feeder (
// Equation(s):
// \register[28][26]~feeder_combout  = \register~69_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(\register~69_combout ),
	.datad(gnd),
	.cin(gnd),
	.combout(\register[28][26]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \register[28][26]~feeder .lut_mask = 16'hF0F0;
defparam \register[28][26]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X66_Y35_N11
dffeas \register[28][26] (
	.clk(!CLK),
	.d(\register[28][26]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~57_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\register[28][26]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \register[28][26] .is_wysiwyg = "true";
defparam \register[28][26] .power_up = "low";
// synopsys translate_on

// Location: FF_X66_Y36_N17
dffeas \register[20][26] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\register~69_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~35_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\register[20][26]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \register[20][26] .is_wysiwyg = "true";
defparam \register[20][26] .power_up = "low";
// synopsys translate_on

// Location: FF_X65_Y35_N3
dffeas \register[24][26] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\register~69_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~34_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\register[24][26]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \register[24][26] .is_wysiwyg = "true";
defparam \register[24][26] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X65_Y35_N2
cycloneive_lcell_comb \Mux37~4 (
// Equation(s):
// \Mux37~4_combout  = (Selector8 & (((Selector7)))) # (!Selector8 & ((Selector7 & ((\register[24][26]~q ))) # (!Selector7 & (\register[16][26]~q ))))

	.dataa(\register[16][26]~q ),
	.datab(Selector8),
	.datac(\register[24][26]~q ),
	.datad(Selector7),
	.cin(gnd),
	.combout(\Mux37~4_combout ),
	.cout());
// synopsys translate_off
defparam \Mux37~4 .lut_mask = 16'hFC22;
defparam \Mux37~4 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X66_Y36_N16
cycloneive_lcell_comb \Mux37~5 (
// Equation(s):
// \Mux37~5_combout  = (Selector8 & ((\Mux37~4_combout  & (\register[28][26]~q )) # (!\Mux37~4_combout  & ((\register[20][26]~q ))))) # (!Selector8 & (((\Mux37~4_combout ))))

	.dataa(Selector8),
	.datab(\register[28][26]~q ),
	.datac(\register[20][26]~q ),
	.datad(\Mux37~4_combout ),
	.cin(gnd),
	.combout(\Mux37~5_combout ),
	.cout());
// synopsys translate_off
defparam \Mux37~5 .lut_mask = 16'hDDA0;
defparam \Mux37~5 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y32_N10
cycloneive_lcell_comb \Mux37~6 (
// Equation(s):
// \Mux37~6_combout  = (Selector10 & (Selector91)) # (!Selector10 & ((Selector91 & (\Mux37~3_combout )) # (!Selector91 & ((\Mux37~5_combout )))))

	.dataa(Selector10),
	.datab(Selector91),
	.datac(\Mux37~3_combout ),
	.datad(\Mux37~5_combout ),
	.cin(gnd),
	.combout(\Mux37~6_combout ),
	.cout());
// synopsys translate_off
defparam \Mux37~6 .lut_mask = 16'hD9C8;
defparam \Mux37~6 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X66_Y34_N10
cycloneive_lcell_comb \register[11][26]~feeder (
// Equation(s):
// \register[11][26]~feeder_combout  = \register~69_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(\register~69_combout ),
	.cin(gnd),
	.combout(\register[11][26]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \register[11][26]~feeder .lut_mask = 16'hFF00;
defparam \register[11][26]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X66_Y34_N11
dffeas \register[11][26] (
	.clk(!CLK),
	.d(\register[11][26]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~47_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\register[11][26]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \register[11][26] .is_wysiwyg = "true";
defparam \register[11][26] .power_up = "low";
// synopsys translate_on

// Location: FF_X63_Y34_N1
dffeas \register[9][26] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\register~69_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~44_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\register[9][26]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \register[9][26] .is_wysiwyg = "true";
defparam \register[9][26] .power_up = "low";
// synopsys translate_on

// Location: FF_X66_Y40_N13
dffeas \register[10][26] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\register~69_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~45_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\register[10][26]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \register[10][26] .is_wysiwyg = "true";
defparam \register[10][26] .power_up = "low";
// synopsys translate_on

// Location: FF_X66_Y40_N3
dffeas \register[8][26] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\register~69_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~46_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\register[8][26]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \register[8][26] .is_wysiwyg = "true";
defparam \register[8][26] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X66_Y40_N12
cycloneive_lcell_comb \Mux37~10 (
// Equation(s):
// \Mux37~10_combout  = (Selector91 & ((Selector10) # ((\register[10][26]~q )))) # (!Selector91 & (!Selector10 & ((\register[8][26]~q ))))

	.dataa(Selector91),
	.datab(Selector10),
	.datac(\register[10][26]~q ),
	.datad(\register[8][26]~q ),
	.cin(gnd),
	.combout(\Mux37~10_combout ),
	.cout());
// synopsys translate_off
defparam \Mux37~10 .lut_mask = 16'hB9A8;
defparam \Mux37~10 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X63_Y34_N30
cycloneive_lcell_comb \Mux37~11 (
// Equation(s):
// \Mux37~11_combout  = (Selector10 & ((\Mux37~10_combout  & (\register[11][26]~q )) # (!\Mux37~10_combout  & ((\register[9][26]~q ))))) # (!Selector10 & (((\Mux37~10_combout ))))

	.dataa(\register[11][26]~q ),
	.datab(\register[9][26]~q ),
	.datac(Selector10),
	.datad(\Mux37~10_combout ),
	.cin(gnd),
	.combout(\Mux37~11_combout ),
	.cout());
// synopsys translate_off
defparam \Mux37~11 .lut_mask = 16'hAFC0;
defparam \Mux37~11 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X69_Y33_N15
dffeas \register[1][26] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\register~69_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~49_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\register[1][26]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \register[1][26] .is_wysiwyg = "true";
defparam \register[1][26] .power_up = "low";
// synopsys translate_on

// Location: FF_X69_Y33_N21
dffeas \register[3][26] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\register~69_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~48_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\register[3][26]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \register[3][26] .is_wysiwyg = "true";
defparam \register[3][26] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X69_Y33_N14
cycloneive_lcell_comb \Mux37~14 (
// Equation(s):
// \Mux37~14_combout  = (Selector9 & ((plif_ifidinstr_l_17 & ((\register[3][26]~q ))) # (!plif_ifidinstr_l_17 & (\register[1][26]~q )))) # (!Selector9 & (((\register[1][26]~q ))))

	.dataa(Selector9),
	.datab(plif_ifidinstr_l_17),
	.datac(\register[1][26]~q ),
	.datad(\register[3][26]~q ),
	.cin(gnd),
	.combout(\Mux37~14_combout ),
	.cout());
// synopsys translate_off
defparam \Mux37~14 .lut_mask = 16'hF870;
defparam \Mux37~14 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y32_N30
cycloneive_lcell_comb \Mux37~15 (
// Equation(s):
// \Mux37~15_combout  = (Selector10 & (((\Mux37~14_combout )))) # (!Selector10 & (\register[2][26]~q  & (Selector91)))

	.dataa(\register[2][26]~q ),
	.datab(Selector10),
	.datac(Selector91),
	.datad(\Mux37~14_combout ),
	.cin(gnd),
	.combout(\Mux37~15_combout ),
	.cout());
// synopsys translate_off
defparam \Mux37~15 .lut_mask = 16'hEC20;
defparam \Mux37~15 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X69_Y31_N29
dffeas \register[5][26] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\register~69_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~59_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\register[5][26]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \register[5][26] .is_wysiwyg = "true";
defparam \register[5][26] .power_up = "low";
// synopsys translate_on

// Location: FF_X69_Y31_N27
dffeas \register[4][26] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\register~69_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~60_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\register[4][26]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \register[4][26] .is_wysiwyg = "true";
defparam \register[4][26] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X69_Y31_N26
cycloneive_lcell_comb \Mux37~12 (
// Equation(s):
// \Mux37~12_combout  = (Selector10 & ((\register[5][26]~q ) # ((Selector91)))) # (!Selector10 & (((\register[4][26]~q  & !Selector91))))

	.dataa(Selector10),
	.datab(\register[5][26]~q ),
	.datac(\register[4][26]~q ),
	.datad(Selector91),
	.cin(gnd),
	.combout(\Mux37~12_combout ),
	.cout());
// synopsys translate_off
defparam \Mux37~12 .lut_mask = 16'hAAD8;
defparam \Mux37~12 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X68_Y31_N15
dffeas \register[7][26] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\register~69_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~43_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\register[7][26]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \register[7][26] .is_wysiwyg = "true";
defparam \register[7][26] .power_up = "low";
// synopsys translate_on

// Location: FF_X68_Y31_N1
dffeas \register[6][26] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\register~69_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~58_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\register[6][26]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \register[6][26] .is_wysiwyg = "true";
defparam \register[6][26] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X68_Y31_N14
cycloneive_lcell_comb \Mux37~13 (
// Equation(s):
// \Mux37~13_combout  = (Selector91 & ((\Mux37~12_combout  & (\register[7][26]~q )) # (!\Mux37~12_combout  & ((\register[6][26]~q ))))) # (!Selector91 & (\Mux37~12_combout ))

	.dataa(Selector91),
	.datab(\Mux37~12_combout ),
	.datac(\register[7][26]~q ),
	.datad(\register[6][26]~q ),
	.cin(gnd),
	.combout(\Mux37~13_combout ),
	.cout());
// synopsys translate_off
defparam \Mux37~13 .lut_mask = 16'hE6C4;
defparam \Mux37~13 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y32_N4
cycloneive_lcell_comb \Mux37~16 (
// Equation(s):
// \Mux37~16_combout  = (Selector8 & ((Selector7) # ((\Mux37~13_combout )))) # (!Selector8 & (!Selector7 & (\Mux37~15_combout )))

	.dataa(Selector8),
	.datab(Selector7),
	.datac(\Mux37~15_combout ),
	.datad(\Mux37~13_combout ),
	.cin(gnd),
	.combout(\Mux37~16_combout ),
	.cout());
// synopsys translate_off
defparam \Mux37~16 .lut_mask = 16'hBA98;
defparam \Mux37~16 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y32_N10
cycloneive_lcell_comb \register[14][26]~feeder (
// Equation(s):
// \register[14][26]~feeder_combout  = \register~69_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(\register~69_combout ),
	.cin(gnd),
	.combout(\register[14][26]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \register[14][26]~feeder .lut_mask = 16'hFF00;
defparam \register[14][26]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X62_Y32_N11
dffeas \register[14][26] (
	.clk(!CLK),
	.d(\register[14][26]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~61_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\register[14][26]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \register[14][26] .is_wysiwyg = "true";
defparam \register[14][26] .power_up = "low";
// synopsys translate_on

// Location: FF_X63_Y37_N11
dffeas \register[15][26] (
	.clk(!CLK),
	.d(\register~69_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~53_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\register[15][26]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \register[15][26] .is_wysiwyg = "true";
defparam \register[15][26] .power_up = "low";
// synopsys translate_on

// Location: FF_X62_Y30_N29
dffeas \register[13][26] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\register~69_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~62_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\register[13][26]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \register[13][26] .is_wysiwyg = "true";
defparam \register[13][26] .power_up = "low";
// synopsys translate_on

// Location: FF_X62_Y30_N19
dffeas \register[12][26] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\register~69_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~52_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\register[12][26]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \register[12][26] .is_wysiwyg = "true";
defparam \register[12][26] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X62_Y30_N28
cycloneive_lcell_comb \Mux37~17 (
// Equation(s):
// \Mux37~17_combout  = (Selector10 & ((Selector91) # ((\register[13][26]~q )))) # (!Selector10 & (!Selector91 & ((\register[12][26]~q ))))

	.dataa(Selector10),
	.datab(Selector91),
	.datac(\register[13][26]~q ),
	.datad(\register[12][26]~q ),
	.cin(gnd),
	.combout(\Mux37~17_combout ),
	.cout());
// synopsys translate_off
defparam \Mux37~17 .lut_mask = 16'hB9A8;
defparam \Mux37~17 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X63_Y37_N20
cycloneive_lcell_comb \Mux37~18 (
// Equation(s):
// \Mux37~18_combout  = (\Mux37~17_combout  & (((\register[15][26]~q ) # (!Selector91)))) # (!\Mux37~17_combout  & (\register[14][26]~q  & ((Selector91))))

	.dataa(\register[14][26]~q ),
	.datab(\register[15][26]~q ),
	.datac(\Mux37~17_combout ),
	.datad(Selector91),
	.cin(gnd),
	.combout(\Mux37~18_combout ),
	.cout());
// synopsys translate_off
defparam \Mux37~18 .lut_mask = 16'hCAF0;
defparam \Mux37~18 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y35_N30
cycloneive_lcell_comb \register~70 (
// Equation(s):
// \register~70_combout  = (WideOr01 & ((\wdat[25]~12_combout ) # ((plif_memwbregsrc_l_1 & plif_memwbrtnaddr_l_25))))

	.dataa(WideOr0),
	.datab(plif_memwbregsrc_l_1),
	.datac(plif_memwbrtnaddr_l_25),
	.datad(wdat_25),
	.cin(gnd),
	.combout(\register~70_combout ),
	.cout());
// synopsys translate_off
defparam \register~70 .lut_mask = 16'hAA80;
defparam \register~70 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y31_N24
cycloneive_lcell_comb \register[29][25]~feeder (
// Equation(s):
// \register[29][25]~feeder_combout  = \register~70_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(\register~70_combout ),
	.datad(gnd),
	.cin(gnd),
	.combout(\register[29][25]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \register[29][25]~feeder .lut_mask = 16'hF0F0;
defparam \register[29][25]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X61_Y31_N25
dffeas \register[29][25] (
	.clk(!CLK),
	.d(\register[29][25]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~28_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\register[29][25]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \register[29][25] .is_wysiwyg = "true";
defparam \register[29][25] .power_up = "low";
// synopsys translate_on

// Location: FF_X61_Y35_N31
dffeas \register[21][25] (
	.clk(!CLK),
	.d(\register~70_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~22_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\register[21][25]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \register[21][25] .is_wysiwyg = "true";
defparam \register[21][25] .power_up = "low";
// synopsys translate_on

// Location: FF_X61_Y37_N21
dffeas \register[25][25] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\register~70_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~24_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\register[25][25]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \register[25][25] .is_wysiwyg = "true";
defparam \register[25][25] .power_up = "low";
// synopsys translate_on

// Location: FF_X62_Y35_N13
dffeas \register[17][25] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\register~70_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~26_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\register[17][25]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \register[17][25] .is_wysiwyg = "true";
defparam \register[17][25] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X61_Y37_N20
cycloneive_lcell_comb \Mux38~0 (
// Equation(s):
// \Mux38~0_combout  = (Selector7 & ((Selector8) # ((\register[25][25]~q )))) # (!Selector7 & (!Selector8 & ((\register[17][25]~q ))))

	.dataa(Selector7),
	.datab(Selector8),
	.datac(\register[25][25]~q ),
	.datad(\register[17][25]~q ),
	.cin(gnd),
	.combout(\Mux38~0_combout ),
	.cout());
// synopsys translate_off
defparam \Mux38~0 .lut_mask = 16'hB9A8;
defparam \Mux38~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X65_Y32_N28
cycloneive_lcell_comb \Mux38~1 (
// Equation(s):
// \Mux38~1_combout  = (Selector8 & ((\Mux38~0_combout  & (\register[29][25]~q )) # (!\Mux38~0_combout  & ((\register[21][25]~q ))))) # (!Selector8 & (((\Mux38~0_combout ))))

	.dataa(\register[29][25]~q ),
	.datab(\register[21][25]~q ),
	.datac(Selector8),
	.datad(\Mux38~0_combout ),
	.cin(gnd),
	.combout(\Mux38~1_combout ),
	.cout());
// synopsys translate_off
defparam \Mux38~1 .lut_mask = 16'hAFC0;
defparam \Mux38~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X65_Y32_N10
cycloneive_lcell_comb \register[23][25]~feeder (
// Equation(s):
// \register[23][25]~feeder_combout  = \register~70_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(\register~70_combout ),
	.cin(gnd),
	.combout(\register[23][25]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \register[23][25]~feeder .lut_mask = 16'hFF00;
defparam \register[23][25]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X65_Y32_N11
dffeas \register[23][25] (
	.clk(!CLK),
	.d(\register[23][25]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~37_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\register[23][25]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \register[23][25] .is_wysiwyg = "true";
defparam \register[23][25] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X65_Y31_N0
cycloneive_lcell_comb \register[31][25]~feeder (
// Equation(s):
// \register[31][25]~feeder_combout  = \register~70_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(\register~70_combout ),
	.datad(gnd),
	.cin(gnd),
	.combout(\register[31][25]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \register[31][25]~feeder .lut_mask = 16'hF0F0;
defparam \register[31][25]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X65_Y31_N1
dffeas \register[31][25] (
	.clk(!CLK),
	.d(\register[31][25]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~40_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\register[31][25]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \register[31][25] .is_wysiwyg = "true";
defparam \register[31][25] .power_up = "low";
// synopsys translate_on

// Location: FF_X60_Y38_N15
dffeas \register[19][25] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\register~70_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~39_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\register[19][25]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \register[19][25] .is_wysiwyg = "true";
defparam \register[19][25] .power_up = "low";
// synopsys translate_on

// Location: FF_X60_Y38_N17
dffeas \register[27][25] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\register~70_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~38_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\register[27][25]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \register[27][25] .is_wysiwyg = "true";
defparam \register[27][25] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X60_Y38_N16
cycloneive_lcell_comb \Mux38~7 (
// Equation(s):
// \Mux38~7_combout  = (Selector7 & (((\register[27][25]~q ) # (Selector8)))) # (!Selector7 & (\register[19][25]~q  & ((!Selector8))))

	.dataa(Selector7),
	.datab(\register[19][25]~q ),
	.datac(\register[27][25]~q ),
	.datad(Selector8),
	.cin(gnd),
	.combout(\Mux38~7_combout ),
	.cout());
// synopsys translate_off
defparam \Mux38~7 .lut_mask = 16'hAAE4;
defparam \Mux38~7 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X65_Y32_N8
cycloneive_lcell_comb \Mux38~8 (
// Equation(s):
// \Mux38~8_combout  = (Selector8 & ((\Mux38~7_combout  & ((\register[31][25]~q ))) # (!\Mux38~7_combout  & (\register[23][25]~q )))) # (!Selector8 & (((\Mux38~7_combout ))))

	.dataa(\register[23][25]~q ),
	.datab(\register[31][25]~q ),
	.datac(Selector8),
	.datad(\Mux38~7_combout ),
	.cin(gnd),
	.combout(\Mux38~8_combout ),
	.cout());
// synopsys translate_off
defparam \Mux38~8 .lut_mask = 16'hCFA0;
defparam \Mux38~8 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X66_Y39_N17
dffeas \register[28][25] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\register~70_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~57_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\register[28][25]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \register[28][25] .is_wysiwyg = "true";
defparam \register[28][25] .power_up = "low";
// synopsys translate_on

// Location: FF_X69_Y38_N29
dffeas \register[20][25] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\register~70_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~35_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\register[20][25]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \register[20][25] .is_wysiwyg = "true";
defparam \register[20][25] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X69_Y38_N28
cycloneive_lcell_comb \Mux38~4 (
// Equation(s):
// \Mux38~4_combout  = (Selector8 & (((\register[20][25]~q ) # (Selector7)))) # (!Selector8 & (\register[16][25]~q  & ((!Selector7))))

	.dataa(\register[16][25]~q ),
	.datab(Selector8),
	.datac(\register[20][25]~q ),
	.datad(Selector7),
	.cin(gnd),
	.combout(\Mux38~4_combout ),
	.cout());
// synopsys translate_off
defparam \Mux38~4 .lut_mask = 16'hCCE2;
defparam \Mux38~4 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X65_Y32_N18
cycloneive_lcell_comb \Mux38~5 (
// Equation(s):
// \Mux38~5_combout  = (Selector7 & ((\Mux38~4_combout  & ((\register[28][25]~q ))) # (!\Mux38~4_combout  & (\register[24][25]~q )))) # (!Selector7 & (((\Mux38~4_combout ))))

	.dataa(\register[24][25]~q ),
	.datab(Selector7),
	.datac(\register[28][25]~q ),
	.datad(\Mux38~4_combout ),
	.cin(gnd),
	.combout(\Mux38~5_combout ),
	.cout());
// synopsys translate_off
defparam \Mux38~5 .lut_mask = 16'hF388;
defparam \Mux38~5 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X68_Y35_N8
cycloneive_lcell_comb \register[30][25]~feeder (
// Equation(s):
// \register[30][25]~feeder_combout  = \register~70_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(\register~70_combout ),
	.cin(gnd),
	.combout(\register[30][25]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \register[30][25]~feeder .lut_mask = 16'hFF00;
defparam \register[30][25]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X68_Y35_N9
dffeas \register[30][25] (
	.clk(!CLK),
	.d(\register[30][25]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~56_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\register[30][25]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \register[30][25] .is_wysiwyg = "true";
defparam \register[30][25] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X68_Y35_N22
cycloneive_lcell_comb \register[26][25]~feeder (
// Equation(s):
// \register[26][25]~feeder_combout  = \register~70_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(\register~70_combout ),
	.cin(gnd),
	.combout(\register[26][25]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \register[26][25]~feeder .lut_mask = 16'hFF00;
defparam \register[26][25]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X68_Y35_N23
dffeas \register[26][25] (
	.clk(!CLK),
	.d(\register[26][25]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~54_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\register[26][25]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \register[26][25] .is_wysiwyg = "true";
defparam \register[26][25] .power_up = "low";
// synopsys translate_on

// Location: FF_X68_Y39_N17
dffeas \register[22][25] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\register~70_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~55_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\register[22][25]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \register[22][25] .is_wysiwyg = "true";
defparam \register[22][25] .power_up = "low";
// synopsys translate_on

// Location: FF_X69_Y35_N27
dffeas \register[18][25] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\register~70_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~33_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\register[18][25]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \register[18][25] .is_wysiwyg = "true";
defparam \register[18][25] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X68_Y39_N16
cycloneive_lcell_comb \Mux38~2 (
// Equation(s):
// \Mux38~2_combout  = (Selector7 & (Selector8)) # (!Selector7 & ((Selector8 & (\register[22][25]~q )) # (!Selector8 & ((\register[18][25]~q )))))

	.dataa(Selector7),
	.datab(Selector8),
	.datac(\register[22][25]~q ),
	.datad(\register[18][25]~q ),
	.cin(gnd),
	.combout(\Mux38~2_combout ),
	.cout());
// synopsys translate_off
defparam \Mux38~2 .lut_mask = 16'hD9C8;
defparam \Mux38~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X68_Y35_N26
cycloneive_lcell_comb \Mux38~3 (
// Equation(s):
// \Mux38~3_combout  = (Selector7 & ((\Mux38~2_combout  & (\register[30][25]~q )) # (!\Mux38~2_combout  & ((\register[26][25]~q ))))) # (!Selector7 & (((\Mux38~2_combout ))))

	.dataa(Selector7),
	.datab(\register[30][25]~q ),
	.datac(\register[26][25]~q ),
	.datad(\Mux38~2_combout ),
	.cin(gnd),
	.combout(\Mux38~3_combout ),
	.cout());
// synopsys translate_off
defparam \Mux38~3 .lut_mask = 16'hDDA0;
defparam \Mux38~3 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X65_Y32_N12
cycloneive_lcell_comb \Mux38~6 (
// Equation(s):
// \Mux38~6_combout  = (Selector10 & (((Selector91)))) # (!Selector10 & ((Selector91 & ((\Mux38~3_combout ))) # (!Selector91 & (\Mux38~5_combout ))))

	.dataa(Selector10),
	.datab(\Mux38~5_combout ),
	.datac(\Mux38~3_combout ),
	.datad(Selector91),
	.cin(gnd),
	.combout(\Mux38~6_combout ),
	.cout());
// synopsys translate_off
defparam \Mux38~6 .lut_mask = 16'hFA44;
defparam \Mux38~6 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X60_Y36_N27
dffeas \register[12][25] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\register~70_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~52_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\register[12][25]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \register[12][25] .is_wysiwyg = "true";
defparam \register[12][25] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X60_Y36_N26
cycloneive_lcell_comb \Mux38~17 (
// Equation(s):
// \Mux38~17_combout  = (Selector10 & ((\register[13][25]~q ) # ((Selector91)))) # (!Selector10 & (((\register[12][25]~q  & !Selector91))))

	.dataa(\register[13][25]~q ),
	.datab(Selector10),
	.datac(\register[12][25]~q ),
	.datad(Selector91),
	.cin(gnd),
	.combout(\Mux38~17_combout ),
	.cout());
// synopsys translate_off
defparam \Mux38~17 .lut_mask = 16'hCCB8;
defparam \Mux38~17 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X60_Y36_N13
dffeas \register[14][25] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\register~70_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~61_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\register[14][25]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \register[14][25] .is_wysiwyg = "true";
defparam \register[14][25] .power_up = "low";
// synopsys translate_on

// Location: FF_X61_Y35_N25
dffeas \register[15][25] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\register~70_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~53_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\register[15][25]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \register[15][25] .is_wysiwyg = "true";
defparam \register[15][25] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X60_Y36_N12
cycloneive_lcell_comb \Mux38~18 (
// Equation(s):
// \Mux38~18_combout  = (\Mux38~17_combout  & (((\register[15][25]~q )) # (!Selector91))) # (!\Mux38~17_combout  & (Selector91 & (\register[14][25]~q )))

	.dataa(\Mux38~17_combout ),
	.datab(Selector91),
	.datac(\register[14][25]~q ),
	.datad(\register[15][25]~q ),
	.cin(gnd),
	.combout(\Mux38~18_combout ),
	.cout());
// synopsys translate_off
defparam \Mux38~18 .lut_mask = 16'hEA62;
defparam \Mux38~18 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X67_Y31_N21
dffeas \register[5][25] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\register~70_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~59_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\register[5][25]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \register[5][25] .is_wysiwyg = "true";
defparam \register[5][25] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X67_Y31_N20
cycloneive_lcell_comb \Mux38~10 (
// Equation(s):
// \Mux38~10_combout  = (Selector91 & (((Selector10)))) # (!Selector91 & ((Selector10 & ((\register[5][25]~q ))) # (!Selector10 & (\register[4][25]~q ))))

	.dataa(\register[4][25]~q ),
	.datab(Selector91),
	.datac(\register[5][25]~q ),
	.datad(Selector10),
	.cin(gnd),
	.combout(\Mux38~10_combout ),
	.cout());
// synopsys translate_off
defparam \Mux38~10 .lut_mask = 16'hFC22;
defparam \Mux38~10 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X66_Y31_N23
dffeas \register[6][25] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\register~70_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~58_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\register[6][25]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \register[6][25] .is_wysiwyg = "true";
defparam \register[6][25] .power_up = "low";
// synopsys translate_on

// Location: FF_X66_Y31_N13
dffeas \register[7][25] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\register~70_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~43_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\register[7][25]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \register[7][25] .is_wysiwyg = "true";
defparam \register[7][25] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X66_Y31_N22
cycloneive_lcell_comb \Mux38~11 (
// Equation(s):
// \Mux38~11_combout  = (\Mux38~10_combout  & (((\register[7][25]~q )) # (!Selector91))) # (!\Mux38~10_combout  & (Selector91 & (\register[6][25]~q )))

	.dataa(\Mux38~10_combout ),
	.datab(Selector91),
	.datac(\register[6][25]~q ),
	.datad(\register[7][25]~q ),
	.cin(gnd),
	.combout(\Mux38~11_combout ),
	.cout());
// synopsys translate_off
defparam \Mux38~11 .lut_mask = 16'hEA62;
defparam \Mux38~11 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X66_Y32_N17
dffeas \register[2][25] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\register~70_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~50_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\register[2][25]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \register[2][25] .is_wysiwyg = "true";
defparam \register[2][25] .power_up = "low";
// synopsys translate_on

// Location: FF_X65_Y36_N29
dffeas \register[3][25] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\register~70_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~48_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\register[3][25]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \register[3][25] .is_wysiwyg = "true";
defparam \register[3][25] .power_up = "low";
// synopsys translate_on

// Location: FF_X65_Y36_N31
dffeas \register[1][25] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\register~70_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~49_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\register[1][25]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \register[1][25] .is_wysiwyg = "true";
defparam \register[1][25] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X65_Y36_N30
cycloneive_lcell_comb \Mux38~14 (
// Equation(s):
// \Mux38~14_combout  = (Selector10 & ((Selector91 & (\register[3][25]~q )) # (!Selector91 & ((\register[1][25]~q )))))

	.dataa(Selector10),
	.datab(\register[3][25]~q ),
	.datac(\register[1][25]~q ),
	.datad(Selector91),
	.cin(gnd),
	.combout(\Mux38~14_combout ),
	.cout());
// synopsys translate_off
defparam \Mux38~14 .lut_mask = 16'h88A0;
defparam \Mux38~14 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X66_Y32_N16
cycloneive_lcell_comb \Mux38~15 (
// Equation(s):
// \Mux38~15_combout  = (\Mux38~14_combout ) # ((!Selector10 & (Selector91 & \register[2][25]~q )))

	.dataa(Selector10),
	.datab(Selector91),
	.datac(\register[2][25]~q ),
	.datad(\Mux38~14_combout ),
	.cin(gnd),
	.combout(\Mux38~15_combout ),
	.cout());
// synopsys translate_off
defparam \Mux38~15 .lut_mask = 16'hFF40;
defparam \Mux38~15 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X65_Y40_N29
dffeas \register[9][25] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\register~70_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~44_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\register[9][25]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \register[9][25] .is_wysiwyg = "true";
defparam \register[9][25] .power_up = "low";
// synopsys translate_on

// Location: FF_X65_Y40_N11
dffeas \register[11][25] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\register~70_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~47_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\register[11][25]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \register[11][25] .is_wysiwyg = "true";
defparam \register[11][25] .power_up = "low";
// synopsys translate_on

// Location: FF_X66_Y40_N7
dffeas \register[8][25] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\register~70_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~46_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\register[8][25]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \register[8][25] .is_wysiwyg = "true";
defparam \register[8][25] .power_up = "low";
// synopsys translate_on

// Location: FF_X66_Y40_N29
dffeas \register[10][25] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\register~70_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~45_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\register[10][25]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \register[10][25] .is_wysiwyg = "true";
defparam \register[10][25] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X66_Y40_N6
cycloneive_lcell_comb \Mux38~12 (
// Equation(s):
// \Mux38~12_combout  = (Selector91 & ((Selector10) # ((\register[10][25]~q )))) # (!Selector91 & (!Selector10 & (\register[8][25]~q )))

	.dataa(Selector91),
	.datab(Selector10),
	.datac(\register[8][25]~q ),
	.datad(\register[10][25]~q ),
	.cin(gnd),
	.combout(\Mux38~12_combout ),
	.cout());
// synopsys translate_off
defparam \Mux38~12 .lut_mask = 16'hBA98;
defparam \Mux38~12 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X65_Y40_N10
cycloneive_lcell_comb \Mux38~13 (
// Equation(s):
// \Mux38~13_combout  = (Selector10 & ((\Mux38~12_combout  & ((\register[11][25]~q ))) # (!\Mux38~12_combout  & (\register[9][25]~q )))) # (!Selector10 & (((\Mux38~12_combout ))))

	.dataa(Selector10),
	.datab(\register[9][25]~q ),
	.datac(\register[11][25]~q ),
	.datad(\Mux38~12_combout ),
	.cin(gnd),
	.combout(\Mux38~13_combout ),
	.cout());
// synopsys translate_off
defparam \Mux38~13 .lut_mask = 16'hF588;
defparam \Mux38~13 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X65_Y32_N16
cycloneive_lcell_comb \Mux38~16 (
// Equation(s):
// \Mux38~16_combout  = (Selector7 & (((Selector8) # (\Mux38~13_combout )))) # (!Selector7 & (\Mux38~15_combout  & (!Selector8)))

	.dataa(\Mux38~15_combout ),
	.datab(Selector7),
	.datac(Selector8),
	.datad(\Mux38~13_combout ),
	.cin(gnd),
	.combout(\Mux38~16_combout ),
	.cout());
// synopsys translate_off
defparam \Mux38~16 .lut_mask = 16'hCEC2;
defparam \Mux38~16 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X67_Y37_N28
cycloneive_lcell_comb \register~71 (
// Equation(s):
// \register~71_combout  = (WideOr01 & ((\wdat[24]~14_combout ) # ((plif_memwbregsrc_l_1 & plif_memwbrtnaddr_l_24))))

	.dataa(WideOr0),
	.datab(plif_memwbregsrc_l_1),
	.datac(plif_memwbrtnaddr_l_24),
	.datad(wdat_24),
	.cin(gnd),
	.combout(\register~71_combout ),
	.cout());
// synopsys translate_off
defparam \register~71 .lut_mask = 16'hAA80;
defparam \register~71 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y36_N4
cycloneive_lcell_comb \register[25][24]~feeder (
// Equation(s):
// \register[25][24]~feeder_combout  = \register~71_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(\register~71_combout ),
	.datad(gnd),
	.cin(gnd),
	.combout(\register[25][24]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \register[25][24]~feeder .lut_mask = 16'hF0F0;
defparam \register[25][24]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X62_Y36_N5
dffeas \register[25][24] (
	.clk(!CLK),
	.d(\register[25][24]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~24_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\register[25][24]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \register[25][24] .is_wysiwyg = "true";
defparam \register[25][24] .power_up = "low";
// synopsys translate_on

// Location: FF_X61_Y31_N7
dffeas \register[29][24] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\register~71_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~28_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\register[29][24]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \register[29][24] .is_wysiwyg = "true";
defparam \register[29][24] .power_up = "low";
// synopsys translate_on

// Location: FF_X62_Y34_N9
dffeas \register[17][24] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\register~71_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~26_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\register[17][24]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \register[17][24] .is_wysiwyg = "true";
defparam \register[17][24] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X62_Y34_N2
cycloneive_lcell_comb \Mux39~0 (
// Equation(s):
// \Mux39~0_combout  = (Selector8 & ((\register[21][24]~q ) # ((Selector7)))) # (!Selector8 & (((\register[17][24]~q  & !Selector7))))

	.dataa(\register[21][24]~q ),
	.datab(Selector8),
	.datac(\register[17][24]~q ),
	.datad(Selector7),
	.cin(gnd),
	.combout(\Mux39~0_combout ),
	.cout());
// synopsys translate_off
defparam \Mux39~0 .lut_mask = 16'hCCB8;
defparam \Mux39~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y31_N6
cycloneive_lcell_comb \Mux39~1 (
// Equation(s):
// \Mux39~1_combout  = (Selector7 & ((\Mux39~0_combout  & ((\register[29][24]~q ))) # (!\Mux39~0_combout  & (\register[25][24]~q )))) # (!Selector7 & (((\Mux39~0_combout ))))

	.dataa(Selector7),
	.datab(\register[25][24]~q ),
	.datac(\register[29][24]~q ),
	.datad(\Mux39~0_combout ),
	.cin(gnd),
	.combout(\Mux39~1_combout ),
	.cout());
// synopsys translate_off
defparam \Mux39~1 .lut_mask = 16'hF588;
defparam \Mux39~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X65_Y34_N31
dffeas \register[16][24] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\register~71_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~36_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\register[16][24]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \register[16][24] .is_wysiwyg = "true";
defparam \register[16][24] .power_up = "low";
// synopsys translate_on

// Location: FF_X66_Y37_N29
dffeas \register[24][24] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\register~71_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~34_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\register[24][24]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \register[24][24] .is_wysiwyg = "true";
defparam \register[24][24] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X65_Y34_N30
cycloneive_lcell_comb \Mux39~4 (
// Equation(s):
// \Mux39~4_combout  = (Selector7 & ((Selector8) # ((\register[24][24]~q )))) # (!Selector7 & (!Selector8 & (\register[16][24]~q )))

	.dataa(Selector7),
	.datab(Selector8),
	.datac(\register[16][24]~q ),
	.datad(\register[24][24]~q ),
	.cin(gnd),
	.combout(\Mux39~4_combout ),
	.cout());
// synopsys translate_off
defparam \Mux39~4 .lut_mask = 16'hBA98;
defparam \Mux39~4 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X65_Y34_N13
dffeas \register[20][24] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\register~71_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~35_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\register[20][24]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \register[20][24] .is_wysiwyg = "true";
defparam \register[20][24] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X65_Y34_N28
cycloneive_lcell_comb \Mux39~5 (
// Equation(s):
// \Mux39~5_combout  = (Selector8 & ((\Mux39~4_combout  & (\register[28][24]~q )) # (!\Mux39~4_combout  & ((\register[20][24]~q ))))) # (!Selector8 & (((\Mux39~4_combout ))))

	.dataa(\register[28][24]~q ),
	.datab(Selector8),
	.datac(\Mux39~4_combout ),
	.datad(\register[20][24]~q ),
	.cin(gnd),
	.combout(\Mux39~5_combout ),
	.cout());
// synopsys translate_off
defparam \Mux39~5 .lut_mask = 16'hBCB0;
defparam \Mux39~5 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X67_Y37_N29
dffeas \register[22][24] (
	.clk(!CLK),
	.d(\register~71_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~55_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\register[22][24]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \register[22][24] .is_wysiwyg = "true";
defparam \register[22][24] .power_up = "low";
// synopsys translate_on

// Location: FF_X68_Y37_N15
dffeas \register[30][24] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\register~71_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~56_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\register[30][24]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \register[30][24] .is_wysiwyg = "true";
defparam \register[30][24] .power_up = "low";
// synopsys translate_on

// Location: FF_X68_Y37_N25
dffeas \register[26][24] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\register~71_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~54_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\register[26][24]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \register[26][24] .is_wysiwyg = "true";
defparam \register[26][24] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X68_Y37_N24
cycloneive_lcell_comb \Mux39~2 (
// Equation(s):
// \Mux39~2_combout  = (Selector8 & (((Selector7)))) # (!Selector8 & ((Selector7 & ((\register[26][24]~q ))) # (!Selector7 & (\register[18][24]~q ))))

	.dataa(\register[18][24]~q ),
	.datab(Selector8),
	.datac(\register[26][24]~q ),
	.datad(Selector7),
	.cin(gnd),
	.combout(\Mux39~2_combout ),
	.cout());
// synopsys translate_off
defparam \Mux39~2 .lut_mask = 16'hFC22;
defparam \Mux39~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X67_Y37_N12
cycloneive_lcell_comb \Mux39~3 (
// Equation(s):
// \Mux39~3_combout  = (Selector8 & ((\Mux39~2_combout  & ((\register[30][24]~q ))) # (!\Mux39~2_combout  & (\register[22][24]~q )))) # (!Selector8 & (((\Mux39~2_combout ))))

	.dataa(Selector8),
	.datab(\register[22][24]~q ),
	.datac(\register[30][24]~q ),
	.datad(\Mux39~2_combout ),
	.cin(gnd),
	.combout(\Mux39~3_combout ),
	.cout());
// synopsys translate_off
defparam \Mux39~3 .lut_mask = 16'hF588;
defparam \Mux39~3 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X65_Y34_N14
cycloneive_lcell_comb \Mux39~6 (
// Equation(s):
// \Mux39~6_combout  = (Selector91 & (((Selector10) # (\Mux39~3_combout )))) # (!Selector91 & (\Mux39~5_combout  & (!Selector10)))

	.dataa(Selector91),
	.datab(\Mux39~5_combout ),
	.datac(Selector10),
	.datad(\Mux39~3_combout ),
	.cin(gnd),
	.combout(\Mux39~6_combout ),
	.cout());
// synopsys translate_off
defparam \Mux39~6 .lut_mask = 16'hAEA4;
defparam \Mux39~6 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X60_Y35_N31
dffeas \register[23][24] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\register~71_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~37_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\register[23][24]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \register[23][24] .is_wysiwyg = "true";
defparam \register[23][24] .power_up = "low";
// synopsys translate_on

// Location: FF_X60_Y35_N25
dffeas \register[19][24] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\register~71_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~39_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\register[19][24]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \register[19][24] .is_wysiwyg = "true";
defparam \register[19][24] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X60_Y35_N30
cycloneive_lcell_comb \Mux39~7 (
// Equation(s):
// \Mux39~7_combout  = (Selector7 & (Selector8)) # (!Selector7 & ((Selector8 & (\register[23][24]~q )) # (!Selector8 & ((\register[19][24]~q )))))

	.dataa(Selector7),
	.datab(Selector8),
	.datac(\register[23][24]~q ),
	.datad(\register[19][24]~q ),
	.cin(gnd),
	.combout(\Mux39~7_combout ),
	.cout());
// synopsys translate_off
defparam \Mux39~7 .lut_mask = 16'hD9C8;
defparam \Mux39~7 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X63_Y35_N30
cycloneive_lcell_comb \register[27][24]~feeder (
// Equation(s):
// \register[27][24]~feeder_combout  = \register~71_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(\register~71_combout ),
	.datad(gnd),
	.cin(gnd),
	.combout(\register[27][24]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \register[27][24]~feeder .lut_mask = 16'hF0F0;
defparam \register[27][24]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X63_Y35_N31
dffeas \register[27][24] (
	.clk(!CLK),
	.d(\register[27][24]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~38_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\register[27][24]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \register[27][24] .is_wysiwyg = "true";
defparam \register[27][24] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X62_Y34_N20
cycloneive_lcell_comb \register[31][24]~feeder (
// Equation(s):
// \register[31][24]~feeder_combout  = \register~71_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(\register~71_combout ),
	.datad(gnd),
	.cin(gnd),
	.combout(\register[31][24]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \register[31][24]~feeder .lut_mask = 16'hF0F0;
defparam \register[31][24]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X62_Y34_N21
dffeas \register[31][24] (
	.clk(!CLK),
	.d(\register[31][24]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~40_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\register[31][24]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \register[31][24] .is_wysiwyg = "true";
defparam \register[31][24] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X62_Y34_N30
cycloneive_lcell_comb \Mux39~8 (
// Equation(s):
// \Mux39~8_combout  = (Selector7 & ((\Mux39~7_combout  & ((\register[31][24]~q ))) # (!\Mux39~7_combout  & (\register[27][24]~q )))) # (!Selector7 & (\Mux39~7_combout ))

	.dataa(Selector7),
	.datab(\Mux39~7_combout ),
	.datac(\register[27][24]~q ),
	.datad(\register[31][24]~q ),
	.cin(gnd),
	.combout(\Mux39~8_combout ),
	.cout());
// synopsys translate_off
defparam \Mux39~8 .lut_mask = 16'hEC64;
defparam \Mux39~8 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X66_Y34_N4
cycloneive_lcell_comb \register[2][24]~feeder (
// Equation(s):
// \register[2][24]~feeder_combout  = \register~71_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(\register~71_combout ),
	.cin(gnd),
	.combout(\register[2][24]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \register[2][24]~feeder .lut_mask = 16'hFF00;
defparam \register[2][24]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X66_Y34_N5
dffeas \register[2][24] (
	.clk(!CLK),
	.d(\register[2][24]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~50_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\register[2][24]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \register[2][24] .is_wysiwyg = "true";
defparam \register[2][24] .power_up = "low";
// synopsys translate_on

// Location: FF_X69_Y33_N23
dffeas \register[1][24] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\register~71_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~49_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\register[1][24]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \register[1][24] .is_wysiwyg = "true";
defparam \register[1][24] .power_up = "low";
// synopsys translate_on

// Location: FF_X69_Y33_N25
dffeas \register[3][24] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\register~71_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~48_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\register[3][24]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \register[3][24] .is_wysiwyg = "true";
defparam \register[3][24] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X69_Y33_N22
cycloneive_lcell_comb \Mux39~14 (
// Equation(s):
// \Mux39~14_combout  = (Selector9 & ((plif_ifidinstr_l_17 & ((\register[3][24]~q ))) # (!plif_ifidinstr_l_17 & (\register[1][24]~q )))) # (!Selector9 & (((\register[1][24]~q ))))

	.dataa(Selector9),
	.datab(plif_ifidinstr_l_17),
	.datac(\register[1][24]~q ),
	.datad(\register[3][24]~q ),
	.cin(gnd),
	.combout(\Mux39~14_combout ),
	.cout());
// synopsys translate_off
defparam \Mux39~14 .lut_mask = 16'hF870;
defparam \Mux39~14 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X65_Y32_N4
cycloneive_lcell_comb \Mux39~15 (
// Equation(s):
// \Mux39~15_combout  = (Selector10 & (((\Mux39~14_combout )))) # (!Selector10 & (\register[2][24]~q  & ((Selector91))))

	.dataa(Selector10),
	.datab(\register[2][24]~q ),
	.datac(\Mux39~14_combout ),
	.datad(Selector91),
	.cin(gnd),
	.combout(\Mux39~15_combout ),
	.cout());
// synopsys translate_off
defparam \Mux39~15 .lut_mask = 16'hE4A0;
defparam \Mux39~15 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X68_Y31_N23
dffeas \register[7][24] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\register~71_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~43_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\register[7][24]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \register[7][24] .is_wysiwyg = "true";
defparam \register[7][24] .power_up = "low";
// synopsys translate_on

// Location: FF_X68_Y31_N17
dffeas \register[6][24] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\register~71_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~58_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\register[6][24]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \register[6][24] .is_wysiwyg = "true";
defparam \register[6][24] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X68_Y31_N22
cycloneive_lcell_comb \Mux39~13 (
// Equation(s):
// \Mux39~13_combout  = (\Mux39~12_combout  & (((\register[7][24]~q )) # (!Selector91))) # (!\Mux39~12_combout  & (Selector91 & ((\register[6][24]~q ))))

	.dataa(\Mux39~12_combout ),
	.datab(Selector91),
	.datac(\register[7][24]~q ),
	.datad(\register[6][24]~q ),
	.cin(gnd),
	.combout(\Mux39~13_combout ),
	.cout());
// synopsys translate_off
defparam \Mux39~13 .lut_mask = 16'hE6A2;
defparam \Mux39~13 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X65_Y32_N26
cycloneive_lcell_comb \Mux39~16 (
// Equation(s):
// \Mux39~16_combout  = (Selector8 & ((Selector7) # ((\Mux39~13_combout )))) # (!Selector8 & (!Selector7 & (\Mux39~15_combout )))

	.dataa(Selector8),
	.datab(Selector7),
	.datac(\Mux39~15_combout ),
	.datad(\Mux39~13_combout ),
	.cin(gnd),
	.combout(\Mux39~16_combout ),
	.cout());
// synopsys translate_off
defparam \Mux39~16 .lut_mask = 16'hBA98;
defparam \Mux39~16 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y36_N26
cycloneive_lcell_comb \register[15][24]~feeder (
// Equation(s):
// \register[15][24]~feeder_combout  = \register~71_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(\register~71_combout ),
	.datad(gnd),
	.cin(gnd),
	.combout(\register[15][24]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \register[15][24]~feeder .lut_mask = 16'hF0F0;
defparam \register[15][24]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X62_Y36_N27
dffeas \register[15][24] (
	.clk(!CLK),
	.d(\register[15][24]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~53_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\register[15][24]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \register[15][24] .is_wysiwyg = "true";
defparam \register[15][24] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X62_Y32_N4
cycloneive_lcell_comb \register[14][24]~feeder (
// Equation(s):
// \register[14][24]~feeder_combout  = \register~71_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(\register~71_combout ),
	.datad(gnd),
	.cin(gnd),
	.combout(\register[14][24]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \register[14][24]~feeder .lut_mask = 16'hF0F0;
defparam \register[14][24]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X62_Y32_N5
dffeas \register[14][24] (
	.clk(!CLK),
	.d(\register[14][24]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~61_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\register[14][24]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \register[14][24] .is_wysiwyg = "true";
defparam \register[14][24] .power_up = "low";
// synopsys translate_on

// Location: FF_X62_Y30_N7
dffeas \register[12][24] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\register~71_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~52_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\register[12][24]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \register[12][24] .is_wysiwyg = "true";
defparam \register[12][24] .power_up = "low";
// synopsys translate_on

// Location: FF_X62_Y30_N25
dffeas \register[13][24] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\register~71_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~62_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\register[13][24]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \register[13][24] .is_wysiwyg = "true";
defparam \register[13][24] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X62_Y30_N6
cycloneive_lcell_comb \Mux39~17 (
// Equation(s):
// \Mux39~17_combout  = (Selector10 & ((Selector91) # ((\register[13][24]~q )))) # (!Selector10 & (!Selector91 & (\register[12][24]~q )))

	.dataa(Selector10),
	.datab(Selector91),
	.datac(\register[12][24]~q ),
	.datad(\register[13][24]~q ),
	.cin(gnd),
	.combout(\Mux39~17_combout ),
	.cout());
// synopsys translate_off
defparam \Mux39~17 .lut_mask = 16'hBA98;
defparam \Mux39~17 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y32_N26
cycloneive_lcell_comb \Mux39~18 (
// Equation(s):
// \Mux39~18_combout  = (Selector91 & ((\Mux39~17_combout  & (\register[15][24]~q )) # (!\Mux39~17_combout  & ((\register[14][24]~q ))))) # (!Selector91 & (((\Mux39~17_combout ))))

	.dataa(\register[15][24]~q ),
	.datab(Selector91),
	.datac(\register[14][24]~q ),
	.datad(\Mux39~17_combout ),
	.cin(gnd),
	.combout(\Mux39~18_combout ),
	.cout());
// synopsys translate_off
defparam \Mux39~18 .lut_mask = 16'hBBC0;
defparam \Mux39~18 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X66_Y34_N2
cycloneive_lcell_comb \register[11][24]~feeder (
// Equation(s):
// \register[11][24]~feeder_combout  = \register~71_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(\register~71_combout ),
	.cin(gnd),
	.combout(\register[11][24]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \register[11][24]~feeder .lut_mask = 16'hFF00;
defparam \register[11][24]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X66_Y34_N3
dffeas \register[11][24] (
	.clk(!CLK),
	.d(\register[11][24]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~47_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\register[11][24]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \register[11][24] .is_wysiwyg = "true";
defparam \register[11][24] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X63_Y34_N4
cycloneive_lcell_comb \register[9][24]~feeder (
// Equation(s):
// \register[9][24]~feeder_combout  = \register~71_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(\register~71_combout ),
	.cin(gnd),
	.combout(\register[9][24]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \register[9][24]~feeder .lut_mask = 16'hFF00;
defparam \register[9][24]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X63_Y34_N5
dffeas \register[9][24] (
	.clk(!CLK),
	.d(\register[9][24]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~44_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\register[9][24]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \register[9][24] .is_wysiwyg = "true";
defparam \register[9][24] .power_up = "low";
// synopsys translate_on

// Location: FF_X67_Y38_N3
dffeas \register[8][24] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\register~71_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~46_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\register[8][24]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \register[8][24] .is_wysiwyg = "true";
defparam \register[8][24] .power_up = "low";
// synopsys translate_on

// Location: FF_X67_Y38_N13
dffeas \register[10][24] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\register~71_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~45_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\register[10][24]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \register[10][24] .is_wysiwyg = "true";
defparam \register[10][24] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X67_Y38_N12
cycloneive_lcell_comb \Mux39~10 (
// Equation(s):
// \Mux39~10_combout  = (Selector10 & (((Selector91)))) # (!Selector10 & ((Selector91 & ((\register[10][24]~q ))) # (!Selector91 & (\register[8][24]~q ))))

	.dataa(Selector10),
	.datab(\register[8][24]~q ),
	.datac(\register[10][24]~q ),
	.datad(Selector91),
	.cin(gnd),
	.combout(\Mux39~10_combout ),
	.cout());
// synopsys translate_off
defparam \Mux39~10 .lut_mask = 16'hFA44;
defparam \Mux39~10 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X63_Y34_N22
cycloneive_lcell_comb \Mux39~11 (
// Equation(s):
// \Mux39~11_combout  = (Selector10 & ((\Mux39~10_combout  & (\register[11][24]~q )) # (!\Mux39~10_combout  & ((\register[9][24]~q ))))) # (!Selector10 & (((\Mux39~10_combout ))))

	.dataa(\register[11][24]~q ),
	.datab(\register[9][24]~q ),
	.datac(Selector10),
	.datad(\Mux39~10_combout ),
	.cin(gnd),
	.combout(\Mux39~11_combout ),
	.cout());
// synopsys translate_off
defparam \Mux39~11 .lut_mask = 16'hAFC0;
defparam \Mux39~11 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y36_N30
cycloneive_lcell_comb \register~72 (
// Equation(s):
// \register~72_combout  = (WideOr01 & ((\wdat[23]~16_combout ) # ((plif_memwbrtnaddr_l_23 & plif_memwbregsrc_l_1))))

	.dataa(plif_memwbrtnaddr_l_23),
	.datab(wdat_23),
	.datac(plif_memwbregsrc_l_1),
	.datad(WideOr0),
	.cin(gnd),
	.combout(\register~72_combout ),
	.cout());
// synopsys translate_off
defparam \register~72 .lut_mask = 16'hEC00;
defparam \register~72 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y34_N18
cycloneive_lcell_comb \register[31][23]~feeder (
// Equation(s):
// \register[31][23]~feeder_combout  = \register~72_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(\register~72_combout ),
	.cin(gnd),
	.combout(\register[31][23]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \register[31][23]~feeder .lut_mask = 16'hFF00;
defparam \register[31][23]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X62_Y34_N19
dffeas \register[31][23] (
	.clk(!CLK),
	.d(\register[31][23]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~40_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\register[31][23]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \register[31][23] .is_wysiwyg = "true";
defparam \register[31][23] .power_up = "low";
// synopsys translate_on

// Location: FF_X62_Y31_N25
dffeas \register[23][23] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\register~72_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~37_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\register[23][23]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \register[23][23] .is_wysiwyg = "true";
defparam \register[23][23] .power_up = "low";
// synopsys translate_on

// Location: FF_X62_Y31_N3
dffeas \register[19][23] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\register~72_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~39_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\register[19][23]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \register[19][23] .is_wysiwyg = "true";
defparam \register[19][23] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X63_Y31_N16
cycloneive_lcell_comb \register[27][23]~feeder (
// Equation(s):
// \register[27][23]~feeder_combout  = \register~72_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(\register~72_combout ),
	.cin(gnd),
	.combout(\register[27][23]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \register[27][23]~feeder .lut_mask = 16'hFF00;
defparam \register[27][23]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X63_Y31_N17
dffeas \register[27][23] (
	.clk(!CLK),
	.d(\register[27][23]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~38_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\register[27][23]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \register[27][23] .is_wysiwyg = "true";
defparam \register[27][23] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X62_Y31_N2
cycloneive_lcell_comb \Mux40~7 (
// Equation(s):
// \Mux40~7_combout  = (Selector8 & (Selector7)) # (!Selector8 & ((Selector7 & ((\register[27][23]~q ))) # (!Selector7 & (\register[19][23]~q ))))

	.dataa(Selector8),
	.datab(Selector7),
	.datac(\register[19][23]~q ),
	.datad(\register[27][23]~q ),
	.cin(gnd),
	.combout(\Mux40~7_combout ),
	.cout());
// synopsys translate_off
defparam \Mux40~7 .lut_mask = 16'hDC98;
defparam \Mux40~7 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X63_Y31_N22
cycloneive_lcell_comb \Mux40~8 (
// Equation(s):
// \Mux40~8_combout  = (Selector8 & ((\Mux40~7_combout  & (\register[31][23]~q )) # (!\Mux40~7_combout  & ((\register[23][23]~q ))))) # (!Selector8 & (((\Mux40~7_combout ))))

	.dataa(\register[31][23]~q ),
	.datab(Selector8),
	.datac(\register[23][23]~q ),
	.datad(\Mux40~7_combout ),
	.cin(gnd),
	.combout(\Mux40~8_combout ),
	.cout());
// synopsys translate_off
defparam \Mux40~8 .lut_mask = 16'hBBC0;
defparam \Mux40~8 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X67_Y30_N10
cycloneive_lcell_comb \register[29][23]~feeder (
// Equation(s):
// \register[29][23]~feeder_combout  = \register~72_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(\register~72_combout ),
	.datad(gnd),
	.cin(gnd),
	.combout(\register[29][23]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \register[29][23]~feeder .lut_mask = 16'hF0F0;
defparam \register[29][23]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X67_Y30_N11
dffeas \register[29][23] (
	.clk(!CLK),
	.d(\register[29][23]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~28_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\register[29][23]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \register[29][23] .is_wysiwyg = "true";
defparam \register[29][23] .power_up = "low";
// synopsys translate_on

// Location: FF_X62_Y33_N29
dffeas \register[21][23] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\register~72_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~22_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\register[21][23]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \register[21][23] .is_wysiwyg = "true";
defparam \register[21][23] .power_up = "low";
// synopsys translate_on

// Location: FF_X62_Y36_N25
dffeas \register[25][23] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\register~72_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~24_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\register[25][23]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \register[25][23] .is_wysiwyg = "true";
defparam \register[25][23] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X62_Y36_N24
cycloneive_lcell_comb \Mux40~0 (
// Equation(s):
// \Mux40~0_combout  = (Selector7 & (((\register[25][23]~q ) # (Selector8)))) # (!Selector7 & (\register[17][23]~q  & ((!Selector8))))

	.dataa(\register[17][23]~q ),
	.datab(Selector7),
	.datac(\register[25][23]~q ),
	.datad(Selector8),
	.cin(gnd),
	.combout(\Mux40~0_combout ),
	.cout());
// synopsys translate_off
defparam \Mux40~0 .lut_mask = 16'hCCE2;
defparam \Mux40~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X67_Y30_N8
cycloneive_lcell_comb \Mux40~1 (
// Equation(s):
// \Mux40~1_combout  = (Selector8 & ((\Mux40~0_combout  & (\register[29][23]~q )) # (!\Mux40~0_combout  & ((\register[21][23]~q ))))) # (!Selector8 & (((\Mux40~0_combout ))))

	.dataa(\register[29][23]~q ),
	.datab(\register[21][23]~q ),
	.datac(Selector8),
	.datad(\Mux40~0_combout ),
	.cin(gnd),
	.combout(\Mux40~1_combout ),
	.cout());
// synopsys translate_off
defparam \Mux40~1 .lut_mask = 16'hAFC0;
defparam \Mux40~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X68_Y34_N14
cycloneive_lcell_comb \register[28][23]~feeder (
// Equation(s):
// \register[28][23]~feeder_combout  = \register~72_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(\register~72_combout ),
	.datad(gnd),
	.cin(gnd),
	.combout(\register[28][23]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \register[28][23]~feeder .lut_mask = 16'hF0F0;
defparam \register[28][23]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X68_Y34_N15
dffeas \register[28][23] (
	.clk(!CLK),
	.d(\register[28][23]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~57_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\register[28][23]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \register[28][23] .is_wysiwyg = "true";
defparam \register[28][23] .power_up = "low";
// synopsys translate_on

// Location: FF_X70_Y38_N29
dffeas \register[24][23] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\register~72_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~34_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\register[24][23]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \register[24][23] .is_wysiwyg = "true";
defparam \register[24][23] .power_up = "low";
// synopsys translate_on

// Location: FF_X69_Y38_N21
dffeas \register[20][23] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\register~72_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~35_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\register[20][23]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \register[20][23] .is_wysiwyg = "true";
defparam \register[20][23] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X69_Y38_N20
cycloneive_lcell_comb \Mux40~4 (
// Equation(s):
// \Mux40~4_combout  = (Selector8 & (((\register[20][23]~q ) # (Selector7)))) # (!Selector8 & (\register[16][23]~q  & ((!Selector7))))

	.dataa(\register[16][23]~q ),
	.datab(Selector8),
	.datac(\register[20][23]~q ),
	.datad(Selector7),
	.cin(gnd),
	.combout(\Mux40~4_combout ),
	.cout());
// synopsys translate_off
defparam \Mux40~4 .lut_mask = 16'hCCE2;
defparam \Mux40~4 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X68_Y34_N28
cycloneive_lcell_comb \Mux40~5 (
// Equation(s):
// \Mux40~5_combout  = (Selector7 & ((\Mux40~4_combout  & (\register[28][23]~q )) # (!\Mux40~4_combout  & ((\register[24][23]~q ))))) # (!Selector7 & (((\Mux40~4_combout ))))

	.dataa(Selector7),
	.datab(\register[28][23]~q ),
	.datac(\register[24][23]~q ),
	.datad(\Mux40~4_combout ),
	.cin(gnd),
	.combout(\Mux40~5_combout ),
	.cout());
// synopsys translate_off
defparam \Mux40~5 .lut_mask = 16'hDDA0;
defparam \Mux40~5 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X68_Y39_N15
dffeas \register[22][23] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\register~72_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~55_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\register[22][23]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \register[22][23] .is_wysiwyg = "true";
defparam \register[22][23] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X68_Y39_N14
cycloneive_lcell_comb \Mux40~2 (
// Equation(s):
// \Mux40~2_combout  = (Selector8 & (((\register[22][23]~q ) # (Selector7)))) # (!Selector8 & (\register[18][23]~q  & ((!Selector7))))

	.dataa(\register[18][23]~q ),
	.datab(Selector8),
	.datac(\register[22][23]~q ),
	.datad(Selector7),
	.cin(gnd),
	.combout(\Mux40~2_combout ),
	.cout());
// synopsys translate_off
defparam \Mux40~2 .lut_mask = 16'hCCE2;
defparam \Mux40~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X68_Y39_N1
dffeas \register[30][23] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\register~72_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~56_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\register[30][23]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \register[30][23] .is_wysiwyg = "true";
defparam \register[30][23] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X68_Y39_N0
cycloneive_lcell_comb \Mux40~3 (
// Equation(s):
// \Mux40~3_combout  = (\Mux40~2_combout  & (((\register[30][23]~q ) # (!Selector7)))) # (!\Mux40~2_combout  & (\register[26][23]~q  & ((Selector7))))

	.dataa(\register[26][23]~q ),
	.datab(\Mux40~2_combout ),
	.datac(\register[30][23]~q ),
	.datad(Selector7),
	.cin(gnd),
	.combout(\Mux40~3_combout ),
	.cout());
// synopsys translate_off
defparam \Mux40~3 .lut_mask = 16'hE2CC;
defparam \Mux40~3 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X67_Y30_N6
cycloneive_lcell_comb \Mux40~6 (
// Equation(s):
// \Mux40~6_combout  = (Selector10 & (Selector91)) # (!Selector10 & ((Selector91 & ((\Mux40~3_combout ))) # (!Selector91 & (\Mux40~5_combout ))))

	.dataa(Selector10),
	.datab(Selector91),
	.datac(\Mux40~5_combout ),
	.datad(\Mux40~3_combout ),
	.cin(gnd),
	.combout(\Mux40~6_combout ),
	.cout());
// synopsys translate_off
defparam \Mux40~6 .lut_mask = 16'hDC98;
defparam \Mux40~6 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X66_Y32_N31
dffeas \register[2][23] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\register~72_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~50_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\register[2][23]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \register[2][23] .is_wysiwyg = "true";
defparam \register[2][23] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X66_Y32_N30
cycloneive_lcell_comb \Mux40~15 (
// Equation(s):
// \Mux40~15_combout  = (Selector10 & (\Mux40~14_combout )) # (!Selector10 & (((Selector91 & \register[2][23]~q ))))

	.dataa(\Mux40~14_combout ),
	.datab(Selector91),
	.datac(\register[2][23]~q ),
	.datad(Selector10),
	.cin(gnd),
	.combout(\Mux40~15_combout ),
	.cout());
// synopsys translate_off
defparam \Mux40~15 .lut_mask = 16'hAAC0;
defparam \Mux40~15 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X65_Y40_N24
cycloneive_lcell_comb \register[9][23]~feeder (
// Equation(s):
// \register[9][23]~feeder_combout  = \register~72_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(\register~72_combout ),
	.datad(gnd),
	.cin(gnd),
	.combout(\register[9][23]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \register[9][23]~feeder .lut_mask = 16'hF0F0;
defparam \register[9][23]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X65_Y40_N25
dffeas \register[9][23] (
	.clk(!CLK),
	.d(\register[9][23]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~44_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\register[9][23]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \register[9][23] .is_wysiwyg = "true";
defparam \register[9][23] .power_up = "low";
// synopsys translate_on

// Location: FF_X65_Y40_N7
dffeas \register[11][23] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\register~72_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~47_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\register[11][23]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \register[11][23] .is_wysiwyg = "true";
defparam \register[11][23] .power_up = "low";
// synopsys translate_on

// Location: FF_X66_Y40_N23
dffeas \register[8][23] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\register~72_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~46_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\register[8][23]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \register[8][23] .is_wysiwyg = "true";
defparam \register[8][23] .power_up = "low";
// synopsys translate_on

// Location: FF_X66_Y40_N25
dffeas \register[10][23] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\register~72_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~45_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\register[10][23]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \register[10][23] .is_wysiwyg = "true";
defparam \register[10][23] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X66_Y40_N22
cycloneive_lcell_comb \Mux40~12 (
// Equation(s):
// \Mux40~12_combout  = (Selector91 & ((Selector10) # ((\register[10][23]~q )))) # (!Selector91 & (!Selector10 & (\register[8][23]~q )))

	.dataa(Selector91),
	.datab(Selector10),
	.datac(\register[8][23]~q ),
	.datad(\register[10][23]~q ),
	.cin(gnd),
	.combout(\Mux40~12_combout ),
	.cout());
// synopsys translate_off
defparam \Mux40~12 .lut_mask = 16'hBA98;
defparam \Mux40~12 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X65_Y40_N6
cycloneive_lcell_comb \Mux40~13 (
// Equation(s):
// \Mux40~13_combout  = (Selector10 & ((\Mux40~12_combout  & ((\register[11][23]~q ))) # (!\Mux40~12_combout  & (\register[9][23]~q )))) # (!Selector10 & (((\Mux40~12_combout ))))

	.dataa(Selector10),
	.datab(\register[9][23]~q ),
	.datac(\register[11][23]~q ),
	.datad(\Mux40~12_combout ),
	.cin(gnd),
	.combout(\Mux40~13_combout ),
	.cout());
// synopsys translate_off
defparam \Mux40~13 .lut_mask = 16'hF588;
defparam \Mux40~13 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X67_Y30_N18
cycloneive_lcell_comb \Mux40~16 (
// Equation(s):
// \Mux40~16_combout  = (Selector8 & (Selector7)) # (!Selector8 & ((Selector7 & ((\Mux40~13_combout ))) # (!Selector7 & (\Mux40~15_combout ))))

	.dataa(Selector8),
	.datab(Selector7),
	.datac(\Mux40~15_combout ),
	.datad(\Mux40~13_combout ),
	.cin(gnd),
	.combout(\Mux40~16_combout ),
	.cout());
// synopsys translate_off
defparam \Mux40~16 .lut_mask = 16'hDC98;
defparam \Mux40~16 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y36_N0
cycloneive_lcell_comb \register[15][23]~feeder (
// Equation(s):
// \register[15][23]~feeder_combout  = \register~72_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(\register~72_combout ),
	.datad(gnd),
	.cin(gnd),
	.combout(\register[15][23]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \register[15][23]~feeder .lut_mask = 16'hF0F0;
defparam \register[15][23]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X61_Y36_N1
dffeas \register[15][23] (
	.clk(!CLK),
	.d(\register[15][23]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~53_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\register[15][23]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \register[15][23] .is_wysiwyg = "true";
defparam \register[15][23] .power_up = "low";
// synopsys translate_on

// Location: FF_X63_Y30_N5
dffeas \register[13][23] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\register~72_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~62_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\register[13][23]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \register[13][23] .is_wysiwyg = "true";
defparam \register[13][23] .power_up = "low";
// synopsys translate_on

// Location: FF_X63_Y30_N23
dffeas \register[12][23] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\register~72_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~52_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\register[12][23]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \register[12][23] .is_wysiwyg = "true";
defparam \register[12][23] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X63_Y30_N22
cycloneive_lcell_comb \Mux40~17 (
// Equation(s):
// \Mux40~17_combout  = (Selector91 & (((Selector10)))) # (!Selector91 & ((Selector10 & (\register[13][23]~q )) # (!Selector10 & ((\register[12][23]~q )))))

	.dataa(Selector91),
	.datab(\register[13][23]~q ),
	.datac(\register[12][23]~q ),
	.datad(Selector10),
	.cin(gnd),
	.combout(\Mux40~17_combout ),
	.cout());
// synopsys translate_off
defparam \Mux40~17 .lut_mask = 16'hEE50;
defparam \Mux40~17 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y32_N28
cycloneive_lcell_comb \register[14][23]~feeder (
// Equation(s):
// \register[14][23]~feeder_combout  = \register~72_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(\register~72_combout ),
	.cin(gnd),
	.combout(\register[14][23]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \register[14][23]~feeder .lut_mask = 16'hFF00;
defparam \register[14][23]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X62_Y32_N29
dffeas \register[14][23] (
	.clk(!CLK),
	.d(\register[14][23]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~61_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\register[14][23]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \register[14][23] .is_wysiwyg = "true";
defparam \register[14][23] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X62_Y32_N22
cycloneive_lcell_comb \Mux40~18 (
// Equation(s):
// \Mux40~18_combout  = (Selector91 & ((\Mux40~17_combout  & (\register[15][23]~q )) # (!\Mux40~17_combout  & ((\register[14][23]~q ))))) # (!Selector91 & (((\Mux40~17_combout ))))

	.dataa(Selector91),
	.datab(\register[15][23]~q ),
	.datac(\Mux40~17_combout ),
	.datad(\register[14][23]~q ),
	.cin(gnd),
	.combout(\Mux40~18_combout ),
	.cout());
// synopsys translate_off
defparam \Mux40~18 .lut_mask = 16'hDAD0;
defparam \Mux40~18 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X69_Y32_N21
dffeas \register[5][23] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\register~72_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~59_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\register[5][23]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \register[5][23] .is_wysiwyg = "true";
defparam \register[5][23] .power_up = "low";
// synopsys translate_on

// Location: FF_X69_Y32_N11
dffeas \register[4][23] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\register~72_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~60_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\register[4][23]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \register[4][23] .is_wysiwyg = "true";
defparam \register[4][23] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X69_Y32_N10
cycloneive_lcell_comb \Mux40~10 (
// Equation(s):
// \Mux40~10_combout  = (Selector91 & (((Selector10)))) # (!Selector91 & ((Selector10 & (\register[5][23]~q )) # (!Selector10 & ((\register[4][23]~q )))))

	.dataa(Selector91),
	.datab(\register[5][23]~q ),
	.datac(\register[4][23]~q ),
	.datad(Selector10),
	.cin(gnd),
	.combout(\Mux40~10_combout ),
	.cout());
// synopsys translate_off
defparam \Mux40~10 .lut_mask = 16'hEE50;
defparam \Mux40~10 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X68_Y31_N31
dffeas \register[7][23] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\register~72_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~43_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\register[7][23]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \register[7][23] .is_wysiwyg = "true";
defparam \register[7][23] .power_up = "low";
// synopsys translate_on

// Location: FF_X68_Y31_N13
dffeas \register[6][23] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\register~72_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~58_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\register[6][23]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \register[6][23] .is_wysiwyg = "true";
defparam \register[6][23] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X68_Y31_N12
cycloneive_lcell_comb \Mux40~11 (
// Equation(s):
// \Mux40~11_combout  = (\Mux40~10_combout  & ((\register[7][23]~q ) # ((!Selector91)))) # (!\Mux40~10_combout  & (((\register[6][23]~q  & Selector91))))

	.dataa(\Mux40~10_combout ),
	.datab(\register[7][23]~q ),
	.datac(\register[6][23]~q ),
	.datad(Selector91),
	.cin(gnd),
	.combout(\Mux40~11_combout ),
	.cout());
// synopsys translate_off
defparam \Mux40~11 .lut_mask = 16'hD8AA;
defparam \Mux40~11 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y36_N14
cycloneive_lcell_comb \register~73 (
// Equation(s):
// \register~73_combout  = (WideOr01 & ((\wdat[22]~18_combout ) # ((plif_memwbrtnaddr_l_22 & plif_memwbregsrc_l_1))))

	.dataa(plif_memwbrtnaddr_l_22),
	.datab(WideOr0),
	.datac(plif_memwbregsrc_l_1),
	.datad(wdat_22),
	.cin(gnd),
	.combout(\register~73_combout ),
	.cout());
// synopsys translate_off
defparam \register~73 .lut_mask = 16'hCC80;
defparam \register~73 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X67_Y30_N30
cycloneive_lcell_comb \register[29][22]~feeder (
// Equation(s):
// \register[29][22]~feeder_combout  = \register~73_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(\register~73_combout ),
	.cin(gnd),
	.combout(\register[29][22]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \register[29][22]~feeder .lut_mask = 16'hFF00;
defparam \register[29][22]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X67_Y30_N31
dffeas \register[29][22] (
	.clk(!CLK),
	.d(\register[29][22]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~28_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\register[29][22]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \register[29][22] .is_wysiwyg = "true";
defparam \register[29][22] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X62_Y36_N2
cycloneive_lcell_comb \register[25][22]~feeder (
// Equation(s):
// \register[25][22]~feeder_combout  = \register~73_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(\register~73_combout ),
	.datad(gnd),
	.cin(gnd),
	.combout(\register[25][22]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \register[25][22]~feeder .lut_mask = 16'hF0F0;
defparam \register[25][22]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X62_Y36_N3
dffeas \register[25][22] (
	.clk(!CLK),
	.d(\register[25][22]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~24_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\register[25][22]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \register[25][22] .is_wysiwyg = "true";
defparam \register[25][22] .power_up = "low";
// synopsys translate_on

// Location: FF_X62_Y34_N17
dffeas \register[17][22] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\register~73_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~26_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\register[17][22]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \register[17][22] .is_wysiwyg = "true";
defparam \register[17][22] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X68_Y36_N8
cycloneive_lcell_comb \register[21][22]~feeder (
// Equation(s):
// \register[21][22]~feeder_combout  = \register~73_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(\register~73_combout ),
	.datad(gnd),
	.cin(gnd),
	.combout(\register[21][22]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \register[21][22]~feeder .lut_mask = 16'hF0F0;
defparam \register[21][22]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X68_Y36_N9
dffeas \register[21][22] (
	.clk(!CLK),
	.d(\register[21][22]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~22_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\register[21][22]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \register[21][22] .is_wysiwyg = "true";
defparam \register[21][22] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X62_Y34_N16
cycloneive_lcell_comb \Mux41~0 (
// Equation(s):
// \Mux41~0_combout  = (Selector7 & (Selector8)) # (!Selector7 & ((Selector8 & ((\register[21][22]~q ))) # (!Selector8 & (\register[17][22]~q ))))

	.dataa(Selector7),
	.datab(Selector8),
	.datac(\register[17][22]~q ),
	.datad(\register[21][22]~q ),
	.cin(gnd),
	.combout(\Mux41~0_combout ),
	.cout());
// synopsys translate_off
defparam \Mux41~0 .lut_mask = 16'hDC98;
defparam \Mux41~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X67_Y30_N16
cycloneive_lcell_comb \Mux41~1 (
// Equation(s):
// \Mux41~1_combout  = (Selector7 & ((\Mux41~0_combout  & (\register[29][22]~q )) # (!\Mux41~0_combout  & ((\register[25][22]~q ))))) # (!Selector7 & (((\Mux41~0_combout ))))

	.dataa(\register[29][22]~q ),
	.datab(Selector7),
	.datac(\register[25][22]~q ),
	.datad(\Mux41~0_combout ),
	.cin(gnd),
	.combout(\Mux41~1_combout ),
	.cout());
// synopsys translate_off
defparam \Mux41~1 .lut_mask = 16'hBBC0;
defparam \Mux41~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X66_Y37_N0
cycloneive_lcell_comb \register[28][22]~feeder (
// Equation(s):
// \register[28][22]~feeder_combout  = \register~73_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(\register~73_combout ),
	.cin(gnd),
	.combout(\register[28][22]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \register[28][22]~feeder .lut_mask = 16'hFF00;
defparam \register[28][22]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X66_Y37_N1
dffeas \register[28][22] (
	.clk(!CLK),
	.d(\register[28][22]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~57_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\register[28][22]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \register[28][22] .is_wysiwyg = "true";
defparam \register[28][22] .power_up = "low";
// synopsys translate_on

// Location: FF_X65_Y37_N9
dffeas \register[16][22] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\register~73_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~36_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\register[16][22]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \register[16][22] .is_wysiwyg = "true";
defparam \register[16][22] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X66_Y37_N18
cycloneive_lcell_comb \register[24][22]~feeder (
// Equation(s):
// \register[24][22]~feeder_combout  = \register~73_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(\register~73_combout ),
	.cin(gnd),
	.combout(\register[24][22]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \register[24][22]~feeder .lut_mask = 16'hFF00;
defparam \register[24][22]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X66_Y37_N19
dffeas \register[24][22] (
	.clk(!CLK),
	.d(\register[24][22]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~34_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\register[24][22]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \register[24][22] .is_wysiwyg = "true";
defparam \register[24][22] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X65_Y37_N8
cycloneive_lcell_comb \Mux41~4 (
// Equation(s):
// \Mux41~4_combout  = (Selector8 & (Selector7)) # (!Selector8 & ((Selector7 & ((\register[24][22]~q ))) # (!Selector7 & (\register[16][22]~q ))))

	.dataa(Selector8),
	.datab(Selector7),
	.datac(\register[16][22]~q ),
	.datad(\register[24][22]~q ),
	.cin(gnd),
	.combout(\Mux41~4_combout ),
	.cout());
// synopsys translate_off
defparam \Mux41~4 .lut_mask = 16'hDC98;
defparam \Mux41~4 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X62_Y37_N19
dffeas \register[20][22] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\register~73_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~35_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\register[20][22]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \register[20][22] .is_wysiwyg = "true";
defparam \register[20][22] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X65_Y37_N10
cycloneive_lcell_comb \Mux41~5 (
// Equation(s):
// \Mux41~5_combout  = (Selector8 & ((\Mux41~4_combout  & (\register[28][22]~q )) # (!\Mux41~4_combout  & ((\register[20][22]~q ))))) # (!Selector8 & (((\Mux41~4_combout ))))

	.dataa(Selector8),
	.datab(\register[28][22]~q ),
	.datac(\Mux41~4_combout ),
	.datad(\register[20][22]~q ),
	.cin(gnd),
	.combout(\Mux41~5_combout ),
	.cout());
// synopsys translate_off
defparam \Mux41~5 .lut_mask = 16'hDAD0;
defparam \Mux41~5 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X69_Y35_N25
dffeas \register[22][22] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\register~73_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~55_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\register[22][22]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \register[22][22] .is_wysiwyg = "true";
defparam \register[22][22] .power_up = "low";
// synopsys translate_on

// Location: FF_X68_Y37_N7
dffeas \register[30][22] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\register~73_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~56_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\register[30][22]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \register[30][22] .is_wysiwyg = "true";
defparam \register[30][22] .power_up = "low";
// synopsys translate_on

// Location: FF_X69_Y35_N11
dffeas \register[18][22] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\register~73_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~33_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\register[18][22]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \register[18][22] .is_wysiwyg = "true";
defparam \register[18][22] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X69_Y35_N10
cycloneive_lcell_comb \Mux41~2 (
// Equation(s):
// \Mux41~2_combout  = (Selector8 & (((Selector7)))) # (!Selector8 & ((Selector7 & (\register[26][22]~q )) # (!Selector7 & ((\register[18][22]~q )))))

	.dataa(\register[26][22]~q ),
	.datab(Selector8),
	.datac(\register[18][22]~q ),
	.datad(Selector7),
	.cin(gnd),
	.combout(\Mux41~2_combout ),
	.cout());
// synopsys translate_off
defparam \Mux41~2 .lut_mask = 16'hEE30;
defparam \Mux41~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X68_Y37_N6
cycloneive_lcell_comb \Mux41~3 (
// Equation(s):
// \Mux41~3_combout  = (Selector8 & ((\Mux41~2_combout  & ((\register[30][22]~q ))) # (!\Mux41~2_combout  & (\register[22][22]~q )))) # (!Selector8 & (((\Mux41~2_combout ))))

	.dataa(Selector8),
	.datab(\register[22][22]~q ),
	.datac(\register[30][22]~q ),
	.datad(\Mux41~2_combout ),
	.cin(gnd),
	.combout(\Mux41~3_combout ),
	.cout());
// synopsys translate_off
defparam \Mux41~3 .lut_mask = 16'hF588;
defparam \Mux41~3 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X67_Y30_N26
cycloneive_lcell_comb \Mux41~6 (
// Equation(s):
// \Mux41~6_combout  = (Selector10 & (Selector91)) # (!Selector10 & ((Selector91 & ((\Mux41~3_combout ))) # (!Selector91 & (\Mux41~5_combout ))))

	.dataa(Selector10),
	.datab(Selector91),
	.datac(\Mux41~5_combout ),
	.datad(\Mux41~3_combout ),
	.cin(gnd),
	.combout(\Mux41~6_combout ),
	.cout());
// synopsys translate_off
defparam \Mux41~6 .lut_mask = 16'hDC98;
defparam \Mux41~6 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X62_Y39_N23
dffeas \register[27][22] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\register~73_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~38_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\register[27][22]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \register[27][22] .is_wysiwyg = "true";
defparam \register[27][22] .power_up = "low";
// synopsys translate_on

// Location: FF_X62_Y39_N21
dffeas \register[31][22] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\register~73_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~40_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\register[31][22]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \register[31][22] .is_wysiwyg = "true";
defparam \register[31][22] .power_up = "low";
// synopsys translate_on

// Location: FF_X62_Y38_N17
dffeas \register[19][22] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\register~73_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~39_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\register[19][22]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \register[19][22] .is_wysiwyg = "true";
defparam \register[19][22] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X62_Y38_N16
cycloneive_lcell_comb \Mux41~7 (
// Equation(s):
// \Mux41~7_combout  = (Selector8 & ((\register[23][22]~q ) # ((Selector7)))) # (!Selector8 & (((\register[19][22]~q  & !Selector7))))

	.dataa(\register[23][22]~q ),
	.datab(Selector8),
	.datac(\register[19][22]~q ),
	.datad(Selector7),
	.cin(gnd),
	.combout(\Mux41~7_combout ),
	.cout());
// synopsys translate_off
defparam \Mux41~7 .lut_mask = 16'hCCB8;
defparam \Mux41~7 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y39_N20
cycloneive_lcell_comb \Mux41~8 (
// Equation(s):
// \Mux41~8_combout  = (Selector7 & ((\Mux41~7_combout  & ((\register[31][22]~q ))) # (!\Mux41~7_combout  & (\register[27][22]~q )))) # (!Selector7 & (((\Mux41~7_combout ))))

	.dataa(\register[27][22]~q ),
	.datab(Selector7),
	.datac(\register[31][22]~q ),
	.datad(\Mux41~7_combout ),
	.cin(gnd),
	.combout(\Mux41~8_combout ),
	.cout());
// synopsys translate_off
defparam \Mux41~8 .lut_mask = 16'hF388;
defparam \Mux41~8 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X61_Y36_N15
dffeas \register[15][22] (
	.clk(!CLK),
	.d(\register~73_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~53_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\register[15][22]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \register[15][22] .is_wysiwyg = "true";
defparam \register[15][22] .power_up = "low";
// synopsys translate_on

// Location: FF_X62_Y30_N5
dffeas \register[13][22] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\register~73_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~62_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\register[13][22]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \register[13][22] .is_wysiwyg = "true";
defparam \register[13][22] .power_up = "low";
// synopsys translate_on

// Location: FF_X62_Y30_N27
dffeas \register[12][22] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\register~73_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~52_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\register[12][22]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \register[12][22] .is_wysiwyg = "true";
defparam \register[12][22] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X62_Y30_N26
cycloneive_lcell_comb \Mux41~17 (
// Equation(s):
// \Mux41~17_combout  = (Selector10 & ((\register[13][22]~q ) # ((Selector91)))) # (!Selector10 & (((\register[12][22]~q  & !Selector91))))

	.dataa(Selector10),
	.datab(\register[13][22]~q ),
	.datac(\register[12][22]~q ),
	.datad(Selector91),
	.cin(gnd),
	.combout(\Mux41~17_combout ),
	.cout());
// synopsys translate_off
defparam \Mux41~17 .lut_mask = 16'hAAD8;
defparam \Mux41~17 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X62_Y32_N31
dffeas \register[14][22] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\register~73_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~61_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\register[14][22]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \register[14][22] .is_wysiwyg = "true";
defparam \register[14][22] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X67_Y30_N22
cycloneive_lcell_comb \Mux41~18 (
// Equation(s):
// \Mux41~18_combout  = (\Mux41~17_combout  & ((\register[15][22]~q ) # ((!Selector91)))) # (!\Mux41~17_combout  & (((Selector91 & \register[14][22]~q ))))

	.dataa(\register[15][22]~q ),
	.datab(\Mux41~17_combout ),
	.datac(Selector91),
	.datad(\register[14][22]~q ),
	.cin(gnd),
	.combout(\Mux41~18_combout ),
	.cout());
// synopsys translate_off
defparam \Mux41~18 .lut_mask = 16'hBC8C;
defparam \Mux41~18 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X66_Y32_N27
dffeas \register[2][22] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\register~73_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~50_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\register[2][22]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \register[2][22] .is_wysiwyg = "true";
defparam \register[2][22] .power_up = "low";
// synopsys translate_on

// Location: FF_X69_Y33_N19
dffeas \register[1][22] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\register~73_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~49_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\register[1][22]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \register[1][22] .is_wysiwyg = "true";
defparam \register[1][22] .power_up = "low";
// synopsys translate_on

// Location: FF_X69_Y33_N5
dffeas \register[3][22] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\register~73_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~48_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\register[3][22]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \register[3][22] .is_wysiwyg = "true";
defparam \register[3][22] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X69_Y33_N18
cycloneive_lcell_comb \Mux41~14 (
// Equation(s):
// \Mux41~14_combout  = (Selector9 & ((plif_ifidinstr_l_17 & ((\register[3][22]~q ))) # (!plif_ifidinstr_l_17 & (\register[1][22]~q )))) # (!Selector9 & (((\register[1][22]~q ))))

	.dataa(Selector9),
	.datab(plif_ifidinstr_l_17),
	.datac(\register[1][22]~q ),
	.datad(\register[3][22]~q ),
	.cin(gnd),
	.combout(\Mux41~14_combout ),
	.cout());
// synopsys translate_off
defparam \Mux41~14 .lut_mask = 16'hF870;
defparam \Mux41~14 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X66_Y32_N26
cycloneive_lcell_comb \Mux41~15 (
// Equation(s):
// \Mux41~15_combout  = (Selector10 & (((\Mux41~14_combout )))) # (!Selector10 & (Selector91 & (\register[2][22]~q )))

	.dataa(Selector10),
	.datab(Selector91),
	.datac(\register[2][22]~q ),
	.datad(\Mux41~14_combout ),
	.cin(gnd),
	.combout(\Mux41~15_combout ),
	.cout());
// synopsys translate_off
defparam \Mux41~15 .lut_mask = 16'hEA40;
defparam \Mux41~15 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X66_Y32_N25
dffeas \register[7][22] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\register~73_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~43_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\register[7][22]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \register[7][22] .is_wysiwyg = "true";
defparam \register[7][22] .power_up = "low";
// synopsys translate_on

// Location: FF_X69_Y31_N1
dffeas \register[5][22] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\register~73_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~59_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\register[5][22]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \register[5][22] .is_wysiwyg = "true";
defparam \register[5][22] .power_up = "low";
// synopsys translate_on

// Location: FF_X69_Y31_N3
dffeas \register[4][22] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\register~73_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~60_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\register[4][22]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \register[4][22] .is_wysiwyg = "true";
defparam \register[4][22] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X69_Y31_N2
cycloneive_lcell_comb \Mux41~12 (
// Equation(s):
// \Mux41~12_combout  = (Selector10 & ((\register[5][22]~q ) # ((Selector91)))) # (!Selector10 & (((\register[4][22]~q  & !Selector91))))

	.dataa(Selector10),
	.datab(\register[5][22]~q ),
	.datac(\register[4][22]~q ),
	.datad(Selector91),
	.cin(gnd),
	.combout(\Mux41~12_combout ),
	.cout());
// synopsys translate_off
defparam \Mux41~12 .lut_mask = 16'hAAD8;
defparam \Mux41~12 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X66_Y32_N24
cycloneive_lcell_comb \Mux41~13 (
// Equation(s):
// \Mux41~13_combout  = (Selector91 & ((\Mux41~12_combout  & ((\register[7][22]~q ))) # (!\Mux41~12_combout  & (\register[6][22]~q )))) # (!Selector91 & (((\Mux41~12_combout ))))

	.dataa(\register[6][22]~q ),
	.datab(Selector91),
	.datac(\register[7][22]~q ),
	.datad(\Mux41~12_combout ),
	.cin(gnd),
	.combout(\Mux41~13_combout ),
	.cout());
// synopsys translate_off
defparam \Mux41~13 .lut_mask = 16'hF388;
defparam \Mux41~13 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X66_Y32_N12
cycloneive_lcell_comb \Mux41~16 (
// Equation(s):
// \Mux41~16_combout  = (Selector8 & ((Selector7) # ((\Mux41~13_combout )))) # (!Selector8 & (!Selector7 & (\Mux41~15_combout )))

	.dataa(Selector8),
	.datab(Selector7),
	.datac(\Mux41~15_combout ),
	.datad(\Mux41~13_combout ),
	.cin(gnd),
	.combout(\Mux41~16_combout ),
	.cout());
// synopsys translate_off
defparam \Mux41~16 .lut_mask = 16'hBA98;
defparam \Mux41~16 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X65_Y40_N15
dffeas \register[11][22] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\register~73_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~47_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\register[11][22]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \register[11][22] .is_wysiwyg = "true";
defparam \register[11][22] .power_up = "low";
// synopsys translate_on

// Location: FF_X65_Y40_N21
dffeas \register[9][22] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\register~73_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~44_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\register[9][22]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \register[9][22] .is_wysiwyg = "true";
defparam \register[9][22] .power_up = "low";
// synopsys translate_on

// Location: FF_X62_Y40_N15
dffeas \register[8][22] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\register~73_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~46_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\register[8][22]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \register[8][22] .is_wysiwyg = "true";
defparam \register[8][22] .power_up = "low";
// synopsys translate_on

// Location: FF_X62_Y40_N1
dffeas \register[10][22] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\register~73_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~45_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\register[10][22]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \register[10][22] .is_wysiwyg = "true";
defparam \register[10][22] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X62_Y40_N0
cycloneive_lcell_comb \Mux41~10 (
// Equation(s):
// \Mux41~10_combout  = (Selector91 & (((\register[10][22]~q ) # (Selector10)))) # (!Selector91 & (\register[8][22]~q  & ((!Selector10))))

	.dataa(Selector91),
	.datab(\register[8][22]~q ),
	.datac(\register[10][22]~q ),
	.datad(Selector10),
	.cin(gnd),
	.combout(\Mux41~10_combout ),
	.cout());
// synopsys translate_off
defparam \Mux41~10 .lut_mask = 16'hAAE4;
defparam \Mux41~10 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X65_Y40_N20
cycloneive_lcell_comb \Mux41~11 (
// Equation(s):
// \Mux41~11_combout  = (Selector10 & ((\Mux41~10_combout  & (\register[11][22]~q )) # (!\Mux41~10_combout  & ((\register[9][22]~q ))))) # (!Selector10 & (((\Mux41~10_combout ))))

	.dataa(Selector10),
	.datab(\register[11][22]~q ),
	.datac(\register[9][22]~q ),
	.datad(\Mux41~10_combout ),
	.cin(gnd),
	.combout(\Mux41~11_combout ),
	.cout());
// synopsys translate_off
defparam \Mux41~11 .lut_mask = 16'hDDA0;
defparam \Mux41~11 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y36_N28
cycloneive_lcell_comb \register~74 (
// Equation(s):
// \register~74_combout  = (WideOr01 & ((\wdat[21]~20_combout ) # ((plif_memwbrtnaddr_l_21 & plif_memwbregsrc_l_1))))

	.dataa(wdat_21),
	.datab(plif_memwbrtnaddr_l_21),
	.datac(plif_memwbregsrc_l_1),
	.datad(WideOr0),
	.cin(gnd),
	.combout(\register~74_combout ),
	.cout());
// synopsys translate_off
defparam \register~74 .lut_mask = 16'hEA00;
defparam \register~74 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X69_Y38_N15
dffeas \register[20][21] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\register~74_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~35_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\register[20][21]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \register[20][21] .is_wysiwyg = "true";
defparam \register[20][21] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X69_Y38_N14
cycloneive_lcell_comb \Mux42~4 (
// Equation(s):
// \Mux42~4_combout  = (Selector8 & (((\register[20][21]~q ) # (Selector7)))) # (!Selector8 & (\register[16][21]~q  & ((!Selector7))))

	.dataa(\register[16][21]~q ),
	.datab(Selector8),
	.datac(\register[20][21]~q ),
	.datad(Selector7),
	.cin(gnd),
	.combout(\Mux42~4_combout ),
	.cout());
// synopsys translate_off
defparam \Mux42~4 .lut_mask = 16'hCCE2;
defparam \Mux42~4 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X69_Y34_N21
dffeas \register[24][21] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\register~74_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~34_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\register[24][21]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \register[24][21] .is_wysiwyg = "true";
defparam \register[24][21] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X68_Y34_N4
cycloneive_lcell_comb \Mux42~5 (
// Equation(s):
// \Mux42~5_combout  = (\Mux42~4_combout  & ((\register[28][21]~q ) # ((!Selector7)))) # (!\Mux42~4_combout  & (((\register[24][21]~q  & Selector7))))

	.dataa(\register[28][21]~q ),
	.datab(\Mux42~4_combout ),
	.datac(\register[24][21]~q ),
	.datad(Selector7),
	.cin(gnd),
	.combout(\Mux42~5_combout ),
	.cout());
// synopsys translate_off
defparam \Mux42~5 .lut_mask = 16'hB8CC;
defparam \Mux42~5 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X68_Y34_N2
cycloneive_lcell_comb \register[30][21]~feeder (
// Equation(s):
// \register[30][21]~feeder_combout  = \register~74_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(\register~74_combout ),
	.cin(gnd),
	.combout(\register[30][21]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \register[30][21]~feeder .lut_mask = 16'hFF00;
defparam \register[30][21]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X68_Y34_N3
dffeas \register[30][21] (
	.clk(!CLK),
	.d(\register[30][21]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~56_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\register[30][21]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \register[30][21] .is_wysiwyg = "true";
defparam \register[30][21] .power_up = "low";
// synopsys translate_on

// Location: FF_X69_Y39_N15
dffeas \register[26][21] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\register~74_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~54_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\register[26][21]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \register[26][21] .is_wysiwyg = "true";
defparam \register[26][21] .power_up = "low";
// synopsys translate_on

// Location: FF_X69_Y39_N9
dffeas \register[18][21] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\register~74_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~33_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\register[18][21]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \register[18][21] .is_wysiwyg = "true";
defparam \register[18][21] .power_up = "low";
// synopsys translate_on

// Location: FF_X67_Y37_N19
dffeas \register[22][21] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\register~74_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~55_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\register[22][21]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \register[22][21] .is_wysiwyg = "true";
defparam \register[22][21] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X69_Y39_N8
cycloneive_lcell_comb \Mux42~2 (
// Equation(s):
// \Mux42~2_combout  = (Selector8 & ((Selector7) # ((\register[22][21]~q )))) # (!Selector8 & (!Selector7 & (\register[18][21]~q )))

	.dataa(Selector8),
	.datab(Selector7),
	.datac(\register[18][21]~q ),
	.datad(\register[22][21]~q ),
	.cin(gnd),
	.combout(\Mux42~2_combout ),
	.cout());
// synopsys translate_off
defparam \Mux42~2 .lut_mask = 16'hBA98;
defparam \Mux42~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X68_Y34_N20
cycloneive_lcell_comb \Mux42~3 (
// Equation(s):
// \Mux42~3_combout  = (Selector7 & ((\Mux42~2_combout  & (\register[30][21]~q )) # (!\Mux42~2_combout  & ((\register[26][21]~q ))))) # (!Selector7 & (((\Mux42~2_combout ))))

	.dataa(Selector7),
	.datab(\register[30][21]~q ),
	.datac(\register[26][21]~q ),
	.datad(\Mux42~2_combout ),
	.cin(gnd),
	.combout(\Mux42~3_combout ),
	.cout());
// synopsys translate_off
defparam \Mux42~3 .lut_mask = 16'hDDA0;
defparam \Mux42~3 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X68_Y34_N18
cycloneive_lcell_comb \Mux42~6 (
// Equation(s):
// \Mux42~6_combout  = (Selector10 & (Selector91)) # (!Selector10 & ((Selector91 & ((\Mux42~3_combout ))) # (!Selector91 & (\Mux42~5_combout ))))

	.dataa(Selector10),
	.datab(Selector91),
	.datac(\Mux42~5_combout ),
	.datad(\Mux42~3_combout ),
	.cin(gnd),
	.combout(\Mux42~6_combout ),
	.cout());
// synopsys translate_off
defparam \Mux42~6 .lut_mask = 16'hDC98;
defparam \Mux42~6 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X62_Y34_N7
dffeas \register[17][21] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\register~74_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~26_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\register[17][21]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \register[17][21] .is_wysiwyg = "true";
defparam \register[17][21] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X60_Y34_N12
cycloneive_lcell_comb \register[25][21]~feeder (
// Equation(s):
// \register[25][21]~feeder_combout  = \register~74_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(\register~74_combout ),
	.datad(gnd),
	.cin(gnd),
	.combout(\register[25][21]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \register[25][21]~feeder .lut_mask = 16'hF0F0;
defparam \register[25][21]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X60_Y34_N13
dffeas \register[25][21] (
	.clk(!CLK),
	.d(\register[25][21]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~24_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\register[25][21]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \register[25][21] .is_wysiwyg = "true";
defparam \register[25][21] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X62_Y34_N6
cycloneive_lcell_comb \Mux42~0 (
// Equation(s):
// \Mux42~0_combout  = (Selector7 & ((Selector8) # ((\register[25][21]~q )))) # (!Selector7 & (!Selector8 & (\register[17][21]~q )))

	.dataa(Selector7),
	.datab(Selector8),
	.datac(\register[17][21]~q ),
	.datad(\register[25][21]~q ),
	.cin(gnd),
	.combout(\Mux42~0_combout ),
	.cout());
// synopsys translate_off
defparam \Mux42~0 .lut_mask = 16'hBA98;
defparam \Mux42~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X63_Y34_N9
dffeas \register[21][21] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\register~74_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~22_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\register[21][21]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \register[21][21] .is_wysiwyg = "true";
defparam \register[21][21] .power_up = "low";
// synopsys translate_on

// Location: FF_X61_Y34_N21
dffeas \register[29][21] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\register~74_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~28_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\register[29][21]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \register[29][21] .is_wysiwyg = "true";
defparam \register[29][21] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X61_Y34_N20
cycloneive_lcell_comb \Mux42~1 (
// Equation(s):
// \Mux42~1_combout  = (\Mux42~0_combout  & (((\register[29][21]~q ) # (!Selector8)))) # (!\Mux42~0_combout  & (\register[21][21]~q  & ((Selector8))))

	.dataa(\Mux42~0_combout ),
	.datab(\register[21][21]~q ),
	.datac(\register[29][21]~q ),
	.datad(Selector8),
	.cin(gnd),
	.combout(\Mux42~1_combout ),
	.cout());
// synopsys translate_off
defparam \Mux42~1 .lut_mask = 16'hE4AA;
defparam \Mux42~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X60_Y35_N23
dffeas \register[23][21] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\register~74_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~37_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\register[23][21]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \register[23][21] .is_wysiwyg = "true";
defparam \register[23][21] .power_up = "low";
// synopsys translate_on

// Location: FF_X62_Y35_N3
dffeas \register[31][21] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\register~74_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~40_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\register[31][21]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \register[31][21] .is_wysiwyg = "true";
defparam \register[31][21] .power_up = "low";
// synopsys translate_on

// Location: FF_X60_Y38_N25
dffeas \register[19][21] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\register~74_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~39_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\register[19][21]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \register[19][21] .is_wysiwyg = "true";
defparam \register[19][21] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X59_Y38_N24
cycloneive_lcell_comb \register[27][21]~feeder (
// Equation(s):
// \register[27][21]~feeder_combout  = \register~74_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(\register~74_combout ),
	.cin(gnd),
	.combout(\register[27][21]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \register[27][21]~feeder .lut_mask = 16'hFF00;
defparam \register[27][21]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X59_Y38_N25
dffeas \register[27][21] (
	.clk(!CLK),
	.d(\register[27][21]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~38_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\register[27][21]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \register[27][21] .is_wysiwyg = "true";
defparam \register[27][21] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X60_Y38_N24
cycloneive_lcell_comb \Mux42~7 (
// Equation(s):
// \Mux42~7_combout  = (Selector8 & (Selector7)) # (!Selector8 & ((Selector7 & ((\register[27][21]~q ))) # (!Selector7 & (\register[19][21]~q ))))

	.dataa(Selector8),
	.datab(Selector7),
	.datac(\register[19][21]~q ),
	.datad(\register[27][21]~q ),
	.cin(gnd),
	.combout(\Mux42~7_combout ),
	.cout());
// synopsys translate_off
defparam \Mux42~7 .lut_mask = 16'hDC98;
defparam \Mux42~7 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y35_N2
cycloneive_lcell_comb \Mux42~8 (
// Equation(s):
// \Mux42~8_combout  = (Selector8 & ((\Mux42~7_combout  & ((\register[31][21]~q ))) # (!\Mux42~7_combout  & (\register[23][21]~q )))) # (!Selector8 & (((\Mux42~7_combout ))))

	.dataa(\register[23][21]~q ),
	.datab(Selector8),
	.datac(\register[31][21]~q ),
	.datad(\Mux42~7_combout ),
	.cin(gnd),
	.combout(\Mux42~8_combout ),
	.cout());
// synopsys translate_off
defparam \Mux42~8 .lut_mask = 16'hF388;
defparam \Mux42~8 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y36_N12
cycloneive_lcell_comb \register[15][21]~feeder (
// Equation(s):
// \register[15][21]~feeder_combout  = \register~74_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(\register~74_combout ),
	.cin(gnd),
	.combout(\register[15][21]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \register[15][21]~feeder .lut_mask = 16'hFF00;
defparam \register[15][21]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X61_Y36_N13
dffeas \register[15][21] (
	.clk(!CLK),
	.d(\register[15][21]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~53_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\register[15][21]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \register[15][21] .is_wysiwyg = "true";
defparam \register[15][21] .power_up = "low";
// synopsys translate_on

// Location: FF_X60_Y34_N11
dffeas \register[14][21] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\register~74_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~61_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\register[14][21]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \register[14][21] .is_wysiwyg = "true";
defparam \register[14][21] .power_up = "low";
// synopsys translate_on

// Location: FF_X62_Y30_N21
dffeas \register[13][21] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\register~74_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~62_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\register[13][21]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \register[13][21] .is_wysiwyg = "true";
defparam \register[13][21] .power_up = "low";
// synopsys translate_on

// Location: FF_X62_Y30_N3
dffeas \register[12][21] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\register~74_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~52_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\register[12][21]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \register[12][21] .is_wysiwyg = "true";
defparam \register[12][21] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X62_Y30_N20
cycloneive_lcell_comb \Mux42~17 (
// Equation(s):
// \Mux42~17_combout  = (Selector10 & ((Selector91) # ((\register[13][21]~q )))) # (!Selector10 & (!Selector91 & ((\register[12][21]~q ))))

	.dataa(Selector10),
	.datab(Selector91),
	.datac(\register[13][21]~q ),
	.datad(\register[12][21]~q ),
	.cin(gnd),
	.combout(\Mux42~17_combout ),
	.cout());
// synopsys translate_off
defparam \Mux42~17 .lut_mask = 16'hB9A8;
defparam \Mux42~17 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y34_N10
cycloneive_lcell_comb \Mux42~18 (
// Equation(s):
// \Mux42~18_combout  = (Selector91 & ((\Mux42~17_combout  & (\register[15][21]~q )) # (!\Mux42~17_combout  & ((\register[14][21]~q ))))) # (!Selector91 & (((\Mux42~17_combout ))))

	.dataa(\register[15][21]~q ),
	.datab(Selector91),
	.datac(\register[14][21]~q ),
	.datad(\Mux42~17_combout ),
	.cin(gnd),
	.combout(\Mux42~18_combout ),
	.cout());
// synopsys translate_off
defparam \Mux42~18 .lut_mask = 16'hBBC0;
defparam \Mux42~18 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X68_Y31_N11
dffeas \register[7][21] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\register~74_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~43_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\register[7][21]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \register[7][21] .is_wysiwyg = "true";
defparam \register[7][21] .power_up = "low";
// synopsys translate_on

// Location: FF_X68_Y31_N25
dffeas \register[6][21] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\register~74_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~58_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\register[6][21]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \register[6][21] .is_wysiwyg = "true";
defparam \register[6][21] .power_up = "low";
// synopsys translate_on

// Location: FF_X67_Y32_N19
dffeas \register[4][21] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\register~74_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~60_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\register[4][21]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \register[4][21] .is_wysiwyg = "true";
defparam \register[4][21] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X67_Y32_N18
cycloneive_lcell_comb \Mux42~10 (
// Equation(s):
// \Mux42~10_combout  = (Selector91 & (((Selector10)))) # (!Selector91 & ((Selector10 & (\register[5][21]~q )) # (!Selector10 & ((\register[4][21]~q )))))

	.dataa(\register[5][21]~q ),
	.datab(Selector91),
	.datac(\register[4][21]~q ),
	.datad(Selector10),
	.cin(gnd),
	.combout(\Mux42~10_combout ),
	.cout());
// synopsys translate_off
defparam \Mux42~10 .lut_mask = 16'hEE30;
defparam \Mux42~10 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X68_Y31_N24
cycloneive_lcell_comb \Mux42~11 (
// Equation(s):
// \Mux42~11_combout  = (Selector91 & ((\Mux42~10_combout  & (\register[7][21]~q )) # (!\Mux42~10_combout  & ((\register[6][21]~q ))))) # (!Selector91 & (((\Mux42~10_combout ))))

	.dataa(\register[7][21]~q ),
	.datab(Selector91),
	.datac(\register[6][21]~q ),
	.datad(\Mux42~10_combout ),
	.cin(gnd),
	.combout(\Mux42~11_combout ),
	.cout());
// synopsys translate_off
defparam \Mux42~11 .lut_mask = 16'hBBC0;
defparam \Mux42~11 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X67_Y34_N27
dffeas \register[11][21] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\register~74_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~47_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\register[11][21]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \register[11][21] .is_wysiwyg = "true";
defparam \register[11][21] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X63_Y34_N14
cycloneive_lcell_comb \register[9][21]~feeder (
// Equation(s):
// \register[9][21]~feeder_combout  = \register~74_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(\register~74_combout ),
	.datad(gnd),
	.cin(gnd),
	.combout(\register[9][21]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \register[9][21]~feeder .lut_mask = 16'hF0F0;
defparam \register[9][21]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X63_Y34_N15
dffeas \register[9][21] (
	.clk(!CLK),
	.d(\register[9][21]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~44_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\register[9][21]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \register[9][21] .is_wysiwyg = "true";
defparam \register[9][21] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X67_Y34_N26
cycloneive_lcell_comb \Mux42~13 (
// Equation(s):
// \Mux42~13_combout  = (\Mux42~12_combout  & (((\register[11][21]~q )) # (!Selector10))) # (!\Mux42~12_combout  & (Selector10 & ((\register[9][21]~q ))))

	.dataa(\Mux42~12_combout ),
	.datab(Selector10),
	.datac(\register[11][21]~q ),
	.datad(\register[9][21]~q ),
	.cin(gnd),
	.combout(\Mux42~13_combout ),
	.cout());
// synopsys translate_off
defparam \Mux42~13 .lut_mask = 16'hE6A2;
defparam \Mux42~13 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X67_Y34_N21
dffeas \register[2][21] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\register~74_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~50_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\register[2][21]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \register[2][21] .is_wysiwyg = "true";
defparam \register[2][21] .power_up = "low";
// synopsys translate_on

// Location: FF_X65_Y33_N5
dffeas \register[3][21] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\register~74_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~48_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\register[3][21]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \register[3][21] .is_wysiwyg = "true";
defparam \register[3][21] .power_up = "low";
// synopsys translate_on

// Location: FF_X65_Y33_N3
dffeas \register[1][21] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\register~74_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~49_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\register[1][21]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \register[1][21] .is_wysiwyg = "true";
defparam \register[1][21] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X65_Y33_N2
cycloneive_lcell_comb \Mux42~14 (
// Equation(s):
// \Mux42~14_combout  = (Selector10 & ((Selector91 & (\register[3][21]~q )) # (!Selector91 & ((\register[1][21]~q )))))

	.dataa(Selector91),
	.datab(\register[3][21]~q ),
	.datac(\register[1][21]~q ),
	.datad(Selector10),
	.cin(gnd),
	.combout(\Mux42~14_combout ),
	.cout());
// synopsys translate_off
defparam \Mux42~14 .lut_mask = 16'hD800;
defparam \Mux42~14 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X68_Y34_N10
cycloneive_lcell_comb \Mux42~15 (
// Equation(s):
// \Mux42~15_combout  = (\Mux42~14_combout ) # ((!Selector10 & (\register[2][21]~q  & Selector91)))

	.dataa(Selector10),
	.datab(\register[2][21]~q ),
	.datac(\Mux42~14_combout ),
	.datad(Selector91),
	.cin(gnd),
	.combout(\Mux42~15_combout ),
	.cout());
// synopsys translate_off
defparam \Mux42~15 .lut_mask = 16'hF4F0;
defparam \Mux42~15 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X68_Y34_N8
cycloneive_lcell_comb \Mux42~16 (
// Equation(s):
// \Mux42~16_combout  = (Selector7 & ((Selector8) # ((\Mux42~13_combout )))) # (!Selector7 & (!Selector8 & ((\Mux42~15_combout ))))

	.dataa(Selector7),
	.datab(Selector8),
	.datac(\Mux42~13_combout ),
	.datad(\Mux42~15_combout ),
	.cin(gnd),
	.combout(\Mux42~16_combout ),
	.cout());
// synopsys translate_off
defparam \Mux42~16 .lut_mask = 16'hB9A8;
defparam \Mux42~16 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y35_N10
cycloneive_lcell_comb \register~75 (
// Equation(s):
// \register~75_combout  = (WideOr01 & ((\wdat[20]~22_combout ) # ((plif_memwbregsrc_l_1 & plif_memwbrtnaddr_l_20))))

	.dataa(WideOr0),
	.datab(plif_memwbregsrc_l_1),
	.datac(wdat_20),
	.datad(plif_memwbrtnaddr_l_20),
	.cin(gnd),
	.combout(\register~75_combout ),
	.cout());
// synopsys translate_off
defparam \register~75 .lut_mask = 16'hA8A0;
defparam \register~75 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X67_Y39_N2
cycloneive_lcell_comb \register[30][20]~feeder (
// Equation(s):
// \register[30][20]~feeder_combout  = \register~75_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(\register~75_combout ),
	.cin(gnd),
	.combout(\register[30][20]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \register[30][20]~feeder .lut_mask = 16'hFF00;
defparam \register[30][20]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X67_Y39_N3
dffeas \register[30][20] (
	.clk(!CLK),
	.d(\register[30][20]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~56_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\register[30][20]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \register[30][20] .is_wysiwyg = "true";
defparam \register[30][20] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X68_Y39_N22
cycloneive_lcell_comb \register[22][20]~feeder (
// Equation(s):
// \register[22][20]~feeder_combout  = \register~75_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(\register~75_combout ),
	.datad(gnd),
	.cin(gnd),
	.combout(\register[22][20]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \register[22][20]~feeder .lut_mask = 16'hF0F0;
defparam \register[22][20]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X68_Y39_N23
dffeas \register[22][20] (
	.clk(!CLK),
	.d(\register[22][20]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~55_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\register[22][20]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \register[22][20] .is_wysiwyg = "true";
defparam \register[22][20] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X67_Y39_N16
cycloneive_lcell_comb \Mux43~3 (
// Equation(s):
// \Mux43~3_combout  = (\Mux43~2_combout  & ((\register[30][20]~q ) # ((!Selector8)))) # (!\Mux43~2_combout  & (((Selector8 & \register[22][20]~q ))))

	.dataa(\Mux43~2_combout ),
	.datab(\register[30][20]~q ),
	.datac(Selector8),
	.datad(\register[22][20]~q ),
	.cin(gnd),
	.combout(\Mux43~3_combout ),
	.cout());
// synopsys translate_off
defparam \Mux43~3 .lut_mask = 16'hDA8A;
defparam \Mux43~3 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X66_Y39_N5
dffeas \register[28][20] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\register~75_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~57_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\register[28][20]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \register[28][20] .is_wysiwyg = "true";
defparam \register[28][20] .power_up = "low";
// synopsys translate_on

// Location: FF_X65_Y39_N15
dffeas \register[20][20] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\register~75_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~35_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\register[20][20]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \register[20][20] .is_wysiwyg = "true";
defparam \register[20][20] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X66_Y39_N14
cycloneive_lcell_comb \Mux43~5 (
// Equation(s):
// \Mux43~5_combout  = (\Mux43~4_combout  & ((\register[28][20]~q ) # ((!Selector8)))) # (!\Mux43~4_combout  & (((\register[20][20]~q  & Selector8))))

	.dataa(\Mux43~4_combout ),
	.datab(\register[28][20]~q ),
	.datac(\register[20][20]~q ),
	.datad(Selector8),
	.cin(gnd),
	.combout(\Mux43~5_combout ),
	.cout());
// synopsys translate_off
defparam \Mux43~5 .lut_mask = 16'hD8AA;
defparam \Mux43~5 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y39_N12
cycloneive_lcell_comb \Mux43~6 (
// Equation(s):
// \Mux43~6_combout  = (Selector91 & ((Selector10) # ((\Mux43~3_combout )))) # (!Selector91 & (!Selector10 & ((\Mux43~5_combout ))))

	.dataa(Selector91),
	.datab(Selector10),
	.datac(\Mux43~3_combout ),
	.datad(\Mux43~5_combout ),
	.cin(gnd),
	.combout(\Mux43~6_combout ),
	.cout());
// synopsys translate_off
defparam \Mux43~6 .lut_mask = 16'hB9A8;
defparam \Mux43~6 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y39_N30
cycloneive_lcell_comb \register[31][20]~feeder (
// Equation(s):
// \register[31][20]~feeder_combout  = \register~75_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(\register~75_combout ),
	.cin(gnd),
	.combout(\register[31][20]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \register[31][20]~feeder .lut_mask = 16'hFF00;
defparam \register[31][20]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X60_Y39_N31
dffeas \register[31][20] (
	.clk(!CLK),
	.d(\register[31][20]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~40_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\register[31][20]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \register[31][20] .is_wysiwyg = "true";
defparam \register[31][20] .power_up = "low";
// synopsys translate_on

// Location: FF_X62_Y39_N11
dffeas \register[27][20] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\register~75_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~38_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\register[27][20]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \register[27][20] .is_wysiwyg = "true";
defparam \register[27][20] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X60_Y40_N8
cycloneive_lcell_comb \register[23][20]~feeder (
// Equation(s):
// \register[23][20]~feeder_combout  = \register~75_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(\register~75_combout ),
	.cin(gnd),
	.combout(\register[23][20]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \register[23][20]~feeder .lut_mask = 16'hFF00;
defparam \register[23][20]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X60_Y40_N9
dffeas \register[23][20] (
	.clk(!CLK),
	.d(\register[23][20]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~37_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\register[23][20]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \register[23][20] .is_wysiwyg = "true";
defparam \register[23][20] .power_up = "low";
// synopsys translate_on

// Location: FF_X62_Y38_N23
dffeas \register[19][20] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\register~75_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~39_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\register[19][20]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \register[19][20] .is_wysiwyg = "true";
defparam \register[19][20] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X62_Y38_N22
cycloneive_lcell_comb \Mux43~7 (
// Equation(s):
// \Mux43~7_combout  = (Selector8 & ((\register[23][20]~q ) # ((Selector7)))) # (!Selector8 & (((\register[19][20]~q  & !Selector7))))

	.dataa(Selector8),
	.datab(\register[23][20]~q ),
	.datac(\register[19][20]~q ),
	.datad(Selector7),
	.cin(gnd),
	.combout(\Mux43~7_combout ),
	.cout());
// synopsys translate_off
defparam \Mux43~7 .lut_mask = 16'hAAD8;
defparam \Mux43~7 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y39_N8
cycloneive_lcell_comb \Mux43~8 (
// Equation(s):
// \Mux43~8_combout  = (Selector7 & ((\Mux43~7_combout  & (\register[31][20]~q )) # (!\Mux43~7_combout  & ((\register[27][20]~q ))))) # (!Selector7 & (((\Mux43~7_combout ))))

	.dataa(\register[31][20]~q ),
	.datab(Selector7),
	.datac(\register[27][20]~q ),
	.datad(\Mux43~7_combout ),
	.cin(gnd),
	.combout(\Mux43~8_combout ),
	.cout());
// synopsys translate_off
defparam \Mux43~8 .lut_mask = 16'hBBC0;
defparam \Mux43~8 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y34_N12
cycloneive_lcell_comb \register[29][20]~feeder (
// Equation(s):
// \register[29][20]~feeder_combout  = \register~75_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(\register~75_combout ),
	.cin(gnd),
	.combout(\register[29][20]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \register[29][20]~feeder .lut_mask = 16'hFF00;
defparam \register[29][20]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X61_Y34_N13
dffeas \register[29][20] (
	.clk(!CLK),
	.d(\register[29][20]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~28_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\register[29][20]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \register[29][20] .is_wysiwyg = "true";
defparam \register[29][20] .power_up = "low";
// synopsys translate_on

// Location: FF_X60_Y34_N5
dffeas \register[25][20] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\register~75_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~24_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\register[25][20]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \register[25][20] .is_wysiwyg = "true";
defparam \register[25][20] .power_up = "low";
// synopsys translate_on

// Location: FF_X60_Y37_N11
dffeas \register[17][20] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\register~75_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~26_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\register[17][20]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \register[17][20] .is_wysiwyg = "true";
defparam \register[17][20] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X61_Y34_N22
cycloneive_lcell_comb \register[21][20]~feeder (
// Equation(s):
// \register[21][20]~feeder_combout  = \register~75_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(\register~75_combout ),
	.cin(gnd),
	.combout(\register[21][20]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \register[21][20]~feeder .lut_mask = 16'hFF00;
defparam \register[21][20]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X61_Y34_N23
dffeas \register[21][20] (
	.clk(!CLK),
	.d(\register[21][20]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~22_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\register[21][20]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \register[21][20] .is_wysiwyg = "true";
defparam \register[21][20] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X60_Y37_N10
cycloneive_lcell_comb \Mux43~0 (
// Equation(s):
// \Mux43~0_combout  = (Selector8 & ((Selector7) # ((\register[21][20]~q )))) # (!Selector8 & (!Selector7 & (\register[17][20]~q )))

	.dataa(Selector8),
	.datab(Selector7),
	.datac(\register[17][20]~q ),
	.datad(\register[21][20]~q ),
	.cin(gnd),
	.combout(\Mux43~0_combout ),
	.cout());
// synopsys translate_off
defparam \Mux43~0 .lut_mask = 16'hBA98;
defparam \Mux43~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y34_N10
cycloneive_lcell_comb \Mux43~1 (
// Equation(s):
// \Mux43~1_combout  = (Selector7 & ((\Mux43~0_combout  & (\register[29][20]~q )) # (!\Mux43~0_combout  & ((\register[25][20]~q ))))) # (!Selector7 & (((\Mux43~0_combout ))))

	.dataa(\register[29][20]~q ),
	.datab(\register[25][20]~q ),
	.datac(Selector7),
	.datad(\Mux43~0_combout ),
	.cin(gnd),
	.combout(\Mux43~1_combout ),
	.cout());
// synopsys translate_off
defparam \Mux43~1 .lut_mask = 16'hAFC0;
defparam \Mux43~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X68_Y31_N5
dffeas \register[6][20] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\register~75_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~58_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\register[6][20]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \register[6][20] .is_wysiwyg = "true";
defparam \register[6][20] .power_up = "low";
// synopsys translate_on

// Location: FF_X68_Y31_N19
dffeas \register[7][20] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\register~75_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~43_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\register[7][20]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \register[7][20] .is_wysiwyg = "true";
defparam \register[7][20] .power_up = "low";
// synopsys translate_on

// Location: FF_X67_Y32_N9
dffeas \register[5][20] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\register~75_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~59_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\register[5][20]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \register[5][20] .is_wysiwyg = "true";
defparam \register[5][20] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X67_Y32_N8
cycloneive_lcell_comb \Mux43~12 (
// Equation(s):
// \Mux43~12_combout  = (Selector91 & (((Selector10)))) # (!Selector91 & ((Selector10 & ((\register[5][20]~q ))) # (!Selector10 & (\register[4][20]~q ))))

	.dataa(\register[4][20]~q ),
	.datab(Selector91),
	.datac(\register[5][20]~q ),
	.datad(Selector10),
	.cin(gnd),
	.combout(\Mux43~12_combout ),
	.cout());
// synopsys translate_off
defparam \Mux43~12 .lut_mask = 16'hFC22;
defparam \Mux43~12 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X68_Y31_N18
cycloneive_lcell_comb \Mux43~13 (
// Equation(s):
// \Mux43~13_combout  = (Selector91 & ((\Mux43~12_combout  & ((\register[7][20]~q ))) # (!\Mux43~12_combout  & (\register[6][20]~q )))) # (!Selector91 & (((\Mux43~12_combout ))))

	.dataa(Selector91),
	.datab(\register[6][20]~q ),
	.datac(\register[7][20]~q ),
	.datad(\Mux43~12_combout ),
	.cin(gnd),
	.combout(\Mux43~13_combout ),
	.cout());
// synopsys translate_off
defparam \Mux43~13 .lut_mask = 16'hF588;
defparam \Mux43~13 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X65_Y36_N25
dffeas \register[3][20] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\register~75_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~48_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\register[3][20]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \register[3][20] .is_wysiwyg = "true";
defparam \register[3][20] .power_up = "low";
// synopsys translate_on

// Location: FF_X65_Y36_N27
dffeas \register[1][20] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\register~75_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~49_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\register[1][20]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \register[1][20] .is_wysiwyg = "true";
defparam \register[1][20] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X65_Y36_N26
cycloneive_lcell_comb \Mux43~14 (
// Equation(s):
// \Mux43~14_combout  = (Selector10 & ((Selector91 & (\register[3][20]~q )) # (!Selector91 & ((\register[1][20]~q )))))

	.dataa(Selector10),
	.datab(\register[3][20]~q ),
	.datac(\register[1][20]~q ),
	.datad(Selector91),
	.cin(gnd),
	.combout(\Mux43~14_combout ),
	.cout());
// synopsys translate_off
defparam \Mux43~14 .lut_mask = 16'h88A0;
defparam \Mux43~14 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X66_Y34_N27
dffeas \register[2][20] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\register~75_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~50_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\register[2][20]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \register[2][20] .is_wysiwyg = "true";
defparam \register[2][20] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X60_Y39_N24
cycloneive_lcell_comb \Mux43~15 (
// Equation(s):
// \Mux43~15_combout  = (\Mux43~14_combout ) # ((Selector91 & (!Selector10 & \register[2][20]~q )))

	.dataa(Selector91),
	.datab(Selector10),
	.datac(\Mux43~14_combout ),
	.datad(\register[2][20]~q ),
	.cin(gnd),
	.combout(\Mux43~15_combout ),
	.cout());
// synopsys translate_off
defparam \Mux43~15 .lut_mask = 16'hF2F0;
defparam \Mux43~15 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y39_N6
cycloneive_lcell_comb \Mux43~16 (
// Equation(s):
// \Mux43~16_combout  = (Selector7 & (((Selector8)))) # (!Selector7 & ((Selector8 & (\Mux43~13_combout )) # (!Selector8 & ((\Mux43~15_combout )))))

	.dataa(\Mux43~13_combout ),
	.datab(Selector7),
	.datac(Selector8),
	.datad(\Mux43~15_combout ),
	.cin(gnd),
	.combout(\Mux43~16_combout ),
	.cout());
// synopsys translate_off
defparam \Mux43~16 .lut_mask = 16'hE3E0;
defparam \Mux43~16 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X65_Y40_N3
dffeas \register[11][20] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\register~75_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~47_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\register[11][20]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \register[11][20] .is_wysiwyg = "true";
defparam \register[11][20] .power_up = "low";
// synopsys translate_on

// Location: FF_X65_Y40_N13
dffeas \register[9][20] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\register~75_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~44_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\register[9][20]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \register[9][20] .is_wysiwyg = "true";
defparam \register[9][20] .power_up = "low";
// synopsys translate_on

// Location: FF_X62_Y41_N25
dffeas \register[10][20] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\register~75_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~45_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\register[10][20]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \register[10][20] .is_wysiwyg = "true";
defparam \register[10][20] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X62_Y41_N24
cycloneive_lcell_comb \Mux43~10 (
// Equation(s):
// \Mux43~10_combout  = (Selector91 & (((\register[10][20]~q ) # (Selector10)))) # (!Selector91 & (\register[8][20]~q  & ((!Selector10))))

	.dataa(\register[8][20]~q ),
	.datab(Selector91),
	.datac(\register[10][20]~q ),
	.datad(Selector10),
	.cin(gnd),
	.combout(\Mux43~10_combout ),
	.cout());
// synopsys translate_off
defparam \Mux43~10 .lut_mask = 16'hCCE2;
defparam \Mux43~10 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X65_Y40_N12
cycloneive_lcell_comb \Mux43~11 (
// Equation(s):
// \Mux43~11_combout  = (Selector10 & ((\Mux43~10_combout  & (\register[11][20]~q )) # (!\Mux43~10_combout  & ((\register[9][20]~q ))))) # (!Selector10 & (((\Mux43~10_combout ))))

	.dataa(Selector10),
	.datab(\register[11][20]~q ),
	.datac(\register[9][20]~q ),
	.datad(\Mux43~10_combout ),
	.cin(gnd),
	.combout(\Mux43~11_combout ),
	.cout());
// synopsys translate_off
defparam \Mux43~11 .lut_mask = 16'hDDA0;
defparam \Mux43~11 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X62_Y30_N15
dffeas \register[12][20] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\register~75_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~52_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\register[12][20]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \register[12][20] .is_wysiwyg = "true";
defparam \register[12][20] .power_up = "low";
// synopsys translate_on

// Location: FF_X62_Y30_N17
dffeas \register[13][20] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\register~75_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~62_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\register[13][20]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \register[13][20] .is_wysiwyg = "true";
defparam \register[13][20] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X62_Y30_N16
cycloneive_lcell_comb \Mux43~17 (
// Equation(s):
// \Mux43~17_combout  = (Selector10 & (((\register[13][20]~q ) # (Selector91)))) # (!Selector10 & (\register[12][20]~q  & ((!Selector91))))

	.dataa(Selector10),
	.datab(\register[12][20]~q ),
	.datac(\register[13][20]~q ),
	.datad(Selector91),
	.cin(gnd),
	.combout(\Mux43~17_combout ),
	.cout());
// synopsys translate_off
defparam \Mux43~17 .lut_mask = 16'hAAE4;
defparam \Mux43~17 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y34_N26
cycloneive_lcell_comb \register[14][20]~feeder (
// Equation(s):
// \register[14][20]~feeder_combout  = \register~75_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(\register~75_combout ),
	.cin(gnd),
	.combout(\register[14][20]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \register[14][20]~feeder .lut_mask = 16'hFF00;
defparam \register[14][20]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X60_Y34_N27
dffeas \register[14][20] (
	.clk(!CLK),
	.d(\register[14][20]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~61_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\register[14][20]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \register[14][20] .is_wysiwyg = "true";
defparam \register[14][20] .power_up = "low";
// synopsys translate_on

// Location: FF_X61_Y35_N11
dffeas \register[15][20] (
	.clk(!CLK),
	.d(\register~75_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~53_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\register[15][20]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \register[15][20] .is_wysiwyg = "true";
defparam \register[15][20] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X60_Y34_N28
cycloneive_lcell_comb \Mux43~18 (
// Equation(s):
// \Mux43~18_combout  = (\Mux43~17_combout  & (((\register[15][20]~q )) # (!Selector91))) # (!\Mux43~17_combout  & (Selector91 & (\register[14][20]~q )))

	.dataa(\Mux43~17_combout ),
	.datab(Selector91),
	.datac(\register[14][20]~q ),
	.datad(\register[15][20]~q ),
	.cin(gnd),
	.combout(\Mux43~18_combout ),
	.cout());
// synopsys translate_off
defparam \Mux43~18 .lut_mask = 16'hEA62;
defparam \Mux43~18 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y36_N6
cycloneive_lcell_comb \register~76 (
// Equation(s):
// \register~76_combout  = (WideOr01 & ((\wdat[19]~24_combout ) # ((plif_memwbrtnaddr_l_19 & plif_memwbregsrc_l_1))))

	.dataa(plif_memwbrtnaddr_l_19),
	.datab(wdat_19),
	.datac(plif_memwbregsrc_l_1),
	.datad(WideOr0),
	.cin(gnd),
	.combout(\register~76_combout ),
	.cout());
// synopsys translate_off
defparam \register~76 .lut_mask = 16'hEC00;
defparam \register~76 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y39_N20
cycloneive_lcell_comb \register[31][19]~feeder (
// Equation(s):
// \register[31][19]~feeder_combout  = \register~76_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(\register~76_combout ),
	.cin(gnd),
	.combout(\register[31][19]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \register[31][19]~feeder .lut_mask = 16'hFF00;
defparam \register[31][19]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X60_Y39_N21
dffeas \register[31][19] (
	.clk(!CLK),
	.d(\register[31][19]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~40_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\register[31][19]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \register[31][19] .is_wysiwyg = "true";
defparam \register[31][19] .power_up = "low";
// synopsys translate_on

// Location: FF_X60_Y35_N1
dffeas \register[23][19] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\register~76_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~37_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\register[23][19]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \register[23][19] .is_wysiwyg = "true";
defparam \register[23][19] .power_up = "low";
// synopsys translate_on

// Location: FF_X60_Y35_N19
dffeas \register[19][19] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\register~76_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~39_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\register[19][19]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \register[19][19] .is_wysiwyg = "true";
defparam \register[19][19] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X60_Y35_N18
cycloneive_lcell_comb \Mux44~7 (
// Equation(s):
// \Mux44~7_combout  = (Selector7 & ((\register[27][19]~q ) # ((Selector8)))) # (!Selector7 & (((\register[19][19]~q  & !Selector8))))

	.dataa(\register[27][19]~q ),
	.datab(Selector7),
	.datac(\register[19][19]~q ),
	.datad(Selector8),
	.cin(gnd),
	.combout(\Mux44~7_combout ),
	.cout());
// synopsys translate_off
defparam \Mux44~7 .lut_mask = 16'hCCB8;
defparam \Mux44~7 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y39_N22
cycloneive_lcell_comb \Mux44~8 (
// Equation(s):
// \Mux44~8_combout  = (Selector8 & ((\Mux44~7_combout  & (\register[31][19]~q )) # (!\Mux44~7_combout  & ((\register[23][19]~q ))))) # (!Selector8 & (((\Mux44~7_combout ))))

	.dataa(\register[31][19]~q ),
	.datab(\register[23][19]~q ),
	.datac(Selector8),
	.datad(\Mux44~7_combout ),
	.cin(gnd),
	.combout(\Mux44~8_combout ),
	.cout());
// synopsys translate_off
defparam \Mux44~8 .lut_mask = 16'hAFC0;
defparam \Mux44~8 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X63_Y34_N25
dffeas \register[21][19] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\register~76_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~22_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\register[21][19]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \register[21][19] .is_wysiwyg = "true";
defparam \register[21][19] .power_up = "low";
// synopsys translate_on

// Location: FF_X62_Y34_N13
dffeas \register[17][19] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\register~76_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~26_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\register[17][19]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \register[17][19] .is_wysiwyg = "true";
defparam \register[17][19] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X62_Y36_N20
cycloneive_lcell_comb \register[25][19]~feeder (
// Equation(s):
// \register[25][19]~feeder_combout  = \register~76_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(\register~76_combout ),
	.datad(gnd),
	.cin(gnd),
	.combout(\register[25][19]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \register[25][19]~feeder .lut_mask = 16'hF0F0;
defparam \register[25][19]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X62_Y36_N21
dffeas \register[25][19] (
	.clk(!CLK),
	.d(\register[25][19]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~24_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\register[25][19]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \register[25][19] .is_wysiwyg = "true";
defparam \register[25][19] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X62_Y34_N12
cycloneive_lcell_comb \Mux44~0 (
// Equation(s):
// \Mux44~0_combout  = (Selector7 & ((Selector8) # ((\register[25][19]~q )))) # (!Selector7 & (!Selector8 & (\register[17][19]~q )))

	.dataa(Selector7),
	.datab(Selector8),
	.datac(\register[17][19]~q ),
	.datad(\register[25][19]~q ),
	.cin(gnd),
	.combout(\Mux44~0_combout ),
	.cout());
// synopsys translate_off
defparam \Mux44~0 .lut_mask = 16'hBA98;
defparam \Mux44~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y34_N0
cycloneive_lcell_comb \register[29][19]~feeder (
// Equation(s):
// \register[29][19]~feeder_combout  = \register~76_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(\register~76_combout ),
	.cin(gnd),
	.combout(\register[29][19]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \register[29][19]~feeder .lut_mask = 16'hFF00;
defparam \register[29][19]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X61_Y34_N1
dffeas \register[29][19] (
	.clk(!CLK),
	.d(\register[29][19]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~28_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\register[29][19]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \register[29][19] .is_wysiwyg = "true";
defparam \register[29][19] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X61_Y34_N26
cycloneive_lcell_comb \Mux44~1 (
// Equation(s):
// \Mux44~1_combout  = (Selector8 & ((\Mux44~0_combout  & ((\register[29][19]~q ))) # (!\Mux44~0_combout  & (\register[21][19]~q )))) # (!Selector8 & (((\Mux44~0_combout ))))

	.dataa(\register[21][19]~q ),
	.datab(Selector8),
	.datac(\Mux44~0_combout ),
	.datad(\register[29][19]~q ),
	.cin(gnd),
	.combout(\Mux44~1_combout ),
	.cout());
// synopsys translate_off
defparam \Mux44~1 .lut_mask = 16'hF838;
defparam \Mux44~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X66_Y39_N21
dffeas \register[24][19] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\register~76_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~34_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\register[24][19]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \register[24][19] .is_wysiwyg = "true";
defparam \register[24][19] .power_up = "low";
// synopsys translate_on

// Location: FF_X66_Y39_N27
dffeas \register[28][19] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\register~76_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~57_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\register[28][19]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \register[28][19] .is_wysiwyg = "true";
defparam \register[28][19] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X69_Y38_N10
cycloneive_lcell_comb \register[16][19]~feeder (
// Equation(s):
// \register[16][19]~feeder_combout  = \register~76_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(\register~76_combout ),
	.cin(gnd),
	.combout(\register[16][19]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \register[16][19]~feeder .lut_mask = 16'hFF00;
defparam \register[16][19]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X69_Y38_N11
dffeas \register[16][19] (
	.clk(!CLK),
	.d(\register[16][19]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~36_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\register[16][19]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \register[16][19] .is_wysiwyg = "true";
defparam \register[16][19] .power_up = "low";
// synopsys translate_on

// Location: FF_X69_Y38_N1
dffeas \register[20][19] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\register~76_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~35_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\register[20][19]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \register[20][19] .is_wysiwyg = "true";
defparam \register[20][19] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X69_Y38_N0
cycloneive_lcell_comb \Mux44~4 (
// Equation(s):
// \Mux44~4_combout  = (Selector8 & (((\register[20][19]~q ) # (Selector7)))) # (!Selector8 & (\register[16][19]~q  & ((!Selector7))))

	.dataa(Selector8),
	.datab(\register[16][19]~q ),
	.datac(\register[20][19]~q ),
	.datad(Selector7),
	.cin(gnd),
	.combout(\Mux44~4_combout ),
	.cout());
// synopsys translate_off
defparam \Mux44~4 .lut_mask = 16'hAAE4;
defparam \Mux44~4 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X66_Y39_N26
cycloneive_lcell_comb \Mux44~5 (
// Equation(s):
// \Mux44~5_combout  = (Selector7 & ((\Mux44~4_combout  & ((\register[28][19]~q ))) # (!\Mux44~4_combout  & (\register[24][19]~q )))) # (!Selector7 & (((\Mux44~4_combout ))))

	.dataa(Selector7),
	.datab(\register[24][19]~q ),
	.datac(\register[28][19]~q ),
	.datad(\Mux44~4_combout ),
	.cin(gnd),
	.combout(\Mux44~5_combout ),
	.cout());
// synopsys translate_off
defparam \Mux44~5 .lut_mask = 16'hF588;
defparam \Mux44~5 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X68_Y39_N19
dffeas \register[30][19] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\register~76_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~56_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\register[30][19]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \register[30][19] .is_wysiwyg = "true";
defparam \register[30][19] .power_up = "low";
// synopsys translate_on

// Location: FF_X69_Y39_N27
dffeas \register[26][19] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\register~76_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~54_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\register[26][19]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \register[26][19] .is_wysiwyg = "true";
defparam \register[26][19] .power_up = "low";
// synopsys translate_on

// Location: FF_X68_Y39_N25
dffeas \register[22][19] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\register~76_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~55_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\register[22][19]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \register[22][19] .is_wysiwyg = "true";
defparam \register[22][19] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X68_Y39_N24
cycloneive_lcell_comb \Mux44~2 (
// Equation(s):
// \Mux44~2_combout  = (Selector8 & (((\register[22][19]~q ) # (Selector7)))) # (!Selector8 & (\register[18][19]~q  & ((!Selector7))))

	.dataa(\register[18][19]~q ),
	.datab(Selector8),
	.datac(\register[22][19]~q ),
	.datad(Selector7),
	.cin(gnd),
	.combout(\Mux44~2_combout ),
	.cout());
// synopsys translate_off
defparam \Mux44~2 .lut_mask = 16'hCCE2;
defparam \Mux44~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X69_Y39_N26
cycloneive_lcell_comb \Mux44~3 (
// Equation(s):
// \Mux44~3_combout  = (Selector7 & ((\Mux44~2_combout  & (\register[30][19]~q )) # (!\Mux44~2_combout  & ((\register[26][19]~q ))))) # (!Selector7 & (((\Mux44~2_combout ))))

	.dataa(Selector7),
	.datab(\register[30][19]~q ),
	.datac(\register[26][19]~q ),
	.datad(\Mux44~2_combout ),
	.cin(gnd),
	.combout(\Mux44~3_combout ),
	.cout());
// synopsys translate_off
defparam \Mux44~3 .lut_mask = 16'hDDA0;
defparam \Mux44~3 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y39_N10
cycloneive_lcell_comb \Mux44~6 (
// Equation(s):
// \Mux44~6_combout  = (Selector91 & ((Selector10) # ((\Mux44~3_combout )))) # (!Selector91 & (!Selector10 & (\Mux44~5_combout )))

	.dataa(Selector91),
	.datab(Selector10),
	.datac(\Mux44~5_combout ),
	.datad(\Mux44~3_combout ),
	.cin(gnd),
	.combout(\Mux44~6_combout ),
	.cout());
// synopsys translate_off
defparam \Mux44~6 .lut_mask = 16'hBA98;
defparam \Mux44~6 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X61_Y36_N7
dffeas \register[15][19] (
	.clk(!CLK),
	.d(\register~76_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~53_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\register[15][19]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \register[15][19] .is_wysiwyg = "true";
defparam \register[15][19] .power_up = "low";
// synopsys translate_on

// Location: FF_X60_Y36_N15
dffeas \register[12][19] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\register~76_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~52_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\register[12][19]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \register[12][19] .is_wysiwyg = "true";
defparam \register[12][19] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X60_Y36_N14
cycloneive_lcell_comb \Mux44~17 (
// Equation(s):
// \Mux44~17_combout  = (Selector10 & ((\register[13][19]~q ) # ((Selector91)))) # (!Selector10 & (((\register[12][19]~q  & !Selector91))))

	.dataa(\register[13][19]~q ),
	.datab(Selector10),
	.datac(\register[12][19]~q ),
	.datad(Selector91),
	.cin(gnd),
	.combout(\Mux44~17_combout ),
	.cout());
// synopsys translate_off
defparam \Mux44~17 .lut_mask = 16'hCCB8;
defparam \Mux44~17 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X60_Y36_N29
dffeas \register[14][19] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\register~76_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~61_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\register[14][19]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \register[14][19] .is_wysiwyg = "true";
defparam \register[14][19] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X60_Y36_N28
cycloneive_lcell_comb \Mux44~18 (
// Equation(s):
// \Mux44~18_combout  = (\Mux44~17_combout  & ((\register[15][19]~q ) # ((!Selector91)))) # (!\Mux44~17_combout  & (((\register[14][19]~q  & Selector91))))

	.dataa(\register[15][19]~q ),
	.datab(\Mux44~17_combout ),
	.datac(\register[14][19]~q ),
	.datad(Selector91),
	.cin(gnd),
	.combout(\Mux44~18_combout ),
	.cout());
// synopsys translate_off
defparam \Mux44~18 .lut_mask = 16'hB8CC;
defparam \Mux44~18 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X68_Y32_N3
dffeas \register[7][19] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\register~76_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~43_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\register[7][19]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \register[7][19] .is_wysiwyg = "true";
defparam \register[7][19] .power_up = "low";
// synopsys translate_on

// Location: FF_X68_Y32_N29
dffeas \register[6][19] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\register~76_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~58_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\register[6][19]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \register[6][19] .is_wysiwyg = "true";
defparam \register[6][19] .power_up = "low";
// synopsys translate_on

// Location: FF_X67_Y32_N29
dffeas \register[5][19] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\register~76_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~59_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\register[5][19]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \register[5][19] .is_wysiwyg = "true";
defparam \register[5][19] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X67_Y32_N28
cycloneive_lcell_comb \Mux44~10 (
// Equation(s):
// \Mux44~10_combout  = (Selector91 & (((Selector10)))) # (!Selector91 & ((Selector10 & ((\register[5][19]~q ))) # (!Selector10 & (\register[4][19]~q ))))

	.dataa(\register[4][19]~q ),
	.datab(Selector91),
	.datac(\register[5][19]~q ),
	.datad(Selector10),
	.cin(gnd),
	.combout(\Mux44~10_combout ),
	.cout());
// synopsys translate_off
defparam \Mux44~10 .lut_mask = 16'hFC22;
defparam \Mux44~10 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X68_Y32_N28
cycloneive_lcell_comb \Mux44~11 (
// Equation(s):
// \Mux44~11_combout  = (Selector91 & ((\Mux44~10_combout  & (\register[7][19]~q )) # (!\Mux44~10_combout  & ((\register[6][19]~q ))))) # (!Selector91 & (((\Mux44~10_combout ))))

	.dataa(Selector91),
	.datab(\register[7][19]~q ),
	.datac(\register[6][19]~q ),
	.datad(\Mux44~10_combout ),
	.cin(gnd),
	.combout(\Mux44~11_combout ),
	.cout());
// synopsys translate_off
defparam \Mux44~11 .lut_mask = 16'hDDA0;
defparam \Mux44~11 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X65_Y36_N17
dffeas \register[3][19] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\register~76_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~48_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\register[3][19]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \register[3][19] .is_wysiwyg = "true";
defparam \register[3][19] .power_up = "low";
// synopsys translate_on

// Location: FF_X65_Y36_N7
dffeas \register[1][19] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\register~76_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~49_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\register[1][19]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \register[1][19] .is_wysiwyg = "true";
defparam \register[1][19] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X65_Y36_N6
cycloneive_lcell_comb \Mux44~14 (
// Equation(s):
// \Mux44~14_combout  = (Selector10 & ((Selector91 & (\register[3][19]~q )) # (!Selector91 & ((\register[1][19]~q )))))

	.dataa(Selector10),
	.datab(\register[3][19]~q ),
	.datac(\register[1][19]~q ),
	.datad(Selector91),
	.cin(gnd),
	.combout(\Mux44~14_combout ),
	.cout());
// synopsys translate_off
defparam \Mux44~14 .lut_mask = 16'h88A0;
defparam \Mux44~14 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y36_N0
cycloneive_lcell_comb \Mux44~15 (
// Equation(s):
// \Mux44~15_combout  = (\Mux44~14_combout ) # ((\register[2][19]~q  & (Selector91 & !Selector10)))

	.dataa(\register[2][19]~q ),
	.datab(Selector91),
	.datac(\Mux44~14_combout ),
	.datad(Selector10),
	.cin(gnd),
	.combout(\Mux44~15_combout ),
	.cout());
// synopsys translate_off
defparam \Mux44~15 .lut_mask = 16'hF0F8;
defparam \Mux44~15 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X66_Y40_N9
dffeas \register[10][19] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\register~76_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~45_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\register[10][19]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \register[10][19] .is_wysiwyg = "true";
defparam \register[10][19] .power_up = "low";
// synopsys translate_on

// Location: FF_X66_Y40_N19
dffeas \register[8][19] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\register~76_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~46_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\register[8][19]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \register[8][19] .is_wysiwyg = "true";
defparam \register[8][19] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X66_Y40_N18
cycloneive_lcell_comb \Mux44~12 (
// Equation(s):
// \Mux44~12_combout  = (Selector10 & (((Selector91)))) # (!Selector10 & ((Selector91 & (\register[10][19]~q )) # (!Selector91 & ((\register[8][19]~q )))))

	.dataa(Selector10),
	.datab(\register[10][19]~q ),
	.datac(\register[8][19]~q ),
	.datad(Selector91),
	.cin(gnd),
	.combout(\Mux44~12_combout ),
	.cout());
// synopsys translate_off
defparam \Mux44~12 .lut_mask = 16'hEE50;
defparam \Mux44~12 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X65_Y40_N31
dffeas \register[11][19] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\register~76_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~47_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\register[11][19]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \register[11][19] .is_wysiwyg = "true";
defparam \register[11][19] .power_up = "low";
// synopsys translate_on

// Location: FF_X65_Y40_N17
dffeas \register[9][19] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\register~76_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~44_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\register[9][19]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \register[9][19] .is_wysiwyg = "true";
defparam \register[9][19] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X65_Y40_N30
cycloneive_lcell_comb \Mux44~13 (
// Equation(s):
// \Mux44~13_combout  = (Selector10 & ((\Mux44~12_combout  & (\register[11][19]~q )) # (!\Mux44~12_combout  & ((\register[9][19]~q ))))) # (!Selector10 & (\Mux44~12_combout ))

	.dataa(Selector10),
	.datab(\Mux44~12_combout ),
	.datac(\register[11][19]~q ),
	.datad(\register[9][19]~q ),
	.cin(gnd),
	.combout(\Mux44~13_combout ),
	.cout());
// synopsys translate_off
defparam \Mux44~13 .lut_mask = 16'hE6C4;
defparam \Mux44~13 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y39_N18
cycloneive_lcell_comb \Mux44~16 (
// Equation(s):
// \Mux44~16_combout  = (Selector7 & (((Selector8) # (\Mux44~13_combout )))) # (!Selector7 & (\Mux44~15_combout  & (!Selector8)))

	.dataa(\Mux44~15_combout ),
	.datab(Selector7),
	.datac(Selector8),
	.datad(\Mux44~13_combout ),
	.cin(gnd),
	.combout(\Mux44~16_combout ),
	.cout());
// synopsys translate_off
defparam \Mux44~16 .lut_mask = 16'hCEC2;
defparam \Mux44~16 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y36_N16
cycloneive_lcell_comb \register~77 (
// Equation(s):
// \register~77_combout  = (WideOr01 & ((\wdat[18]~26_combout ) # ((plif_memwbregsrc_l_1 & plif_memwbrtnaddr_l_18))))

	.dataa(plif_memwbregsrc_l_1),
	.datab(WideOr0),
	.datac(plif_memwbrtnaddr_l_18),
	.datad(wdat_18),
	.cin(gnd),
	.combout(\register~77_combout ),
	.cout());
// synopsys translate_off
defparam \register~77 .lut_mask = 16'hCC80;
defparam \register~77 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X68_Y39_N20
cycloneive_lcell_comb \register[22][18]~feeder (
// Equation(s):
// \register[22][18]~feeder_combout  = \register~77_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(\register~77_combout ),
	.datad(gnd),
	.cin(gnd),
	.combout(\register[22][18]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \register[22][18]~feeder .lut_mask = 16'hF0F0;
defparam \register[22][18]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X68_Y39_N21
dffeas \register[22][18] (
	.clk(!CLK),
	.d(\register[22][18]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~55_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\register[22][18]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \register[22][18] .is_wysiwyg = "true";
defparam \register[22][18] .power_up = "low";
// synopsys translate_on

// Location: FF_X68_Y39_N11
dffeas \register[30][18] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\register~77_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~56_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\register[30][18]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \register[30][18] .is_wysiwyg = "true";
defparam \register[30][18] .power_up = "low";
// synopsys translate_on

// Location: FF_X69_Y39_N19
dffeas \register[26][18] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\register~77_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~54_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\register[26][18]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \register[26][18] .is_wysiwyg = "true";
defparam \register[26][18] .power_up = "low";
// synopsys translate_on

// Location: FF_X69_Y39_N21
dffeas \register[18][18] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\register~77_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~33_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\register[18][18]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \register[18][18] .is_wysiwyg = "true";
defparam \register[18][18] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X69_Y39_N18
cycloneive_lcell_comb \Mux45~2 (
// Equation(s):
// \Mux45~2_combout  = (Selector8 & (Selector7)) # (!Selector8 & ((Selector7 & (\register[26][18]~q )) # (!Selector7 & ((\register[18][18]~q )))))

	.dataa(Selector8),
	.datab(Selector7),
	.datac(\register[26][18]~q ),
	.datad(\register[18][18]~q ),
	.cin(gnd),
	.combout(\Mux45~2_combout ),
	.cout());
// synopsys translate_off
defparam \Mux45~2 .lut_mask = 16'hD9C8;
defparam \Mux45~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X68_Y39_N10
cycloneive_lcell_comb \Mux45~3 (
// Equation(s):
// \Mux45~3_combout  = (Selector8 & ((\Mux45~2_combout  & ((\register[30][18]~q ))) # (!\Mux45~2_combout  & (\register[22][18]~q )))) # (!Selector8 & (((\Mux45~2_combout ))))

	.dataa(Selector8),
	.datab(\register[22][18]~q ),
	.datac(\register[30][18]~q ),
	.datad(\Mux45~2_combout ),
	.cin(gnd),
	.combout(\Mux45~3_combout ),
	.cout());
// synopsys translate_off
defparam \Mux45~3 .lut_mask = 16'hF588;
defparam \Mux45~3 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X66_Y39_N0
cycloneive_lcell_comb \register[24][18]~feeder (
// Equation(s):
// \register[24][18]~feeder_combout  = \register~77_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(\register~77_combout ),
	.datad(gnd),
	.cin(gnd),
	.combout(\register[24][18]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \register[24][18]~feeder .lut_mask = 16'hF0F0;
defparam \register[24][18]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X66_Y39_N1
dffeas \register[24][18] (
	.clk(!CLK),
	.d(\register[24][18]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~34_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\register[24][18]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \register[24][18] .is_wysiwyg = "true";
defparam \register[24][18] .power_up = "low";
// synopsys translate_on

// Location: FF_X65_Y39_N21
dffeas \register[16][18] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\register~77_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~36_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\register[16][18]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \register[16][18] .is_wysiwyg = "true";
defparam \register[16][18] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X65_Y39_N20
cycloneive_lcell_comb \Mux45~4 (
// Equation(s):
// \Mux45~4_combout  = (Selector7 & ((\register[24][18]~q ) # ((Selector8)))) # (!Selector7 & (((\register[16][18]~q  & !Selector8))))

	.dataa(Selector7),
	.datab(\register[24][18]~q ),
	.datac(\register[16][18]~q ),
	.datad(Selector8),
	.cin(gnd),
	.combout(\Mux45~4_combout ),
	.cout());
// synopsys translate_off
defparam \Mux45~4 .lut_mask = 16'hAAD8;
defparam \Mux45~4 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X65_Y39_N3
dffeas \register[20][18] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\register~77_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~35_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\register[20][18]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \register[20][18] .is_wysiwyg = "true";
defparam \register[20][18] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X66_Y39_N8
cycloneive_lcell_comb \Mux45~5 (
// Equation(s):
// \Mux45~5_combout  = (\Mux45~4_combout  & ((\register[28][18]~q ) # ((!Selector8)))) # (!\Mux45~4_combout  & (((\register[20][18]~q  & Selector8))))

	.dataa(\register[28][18]~q ),
	.datab(\Mux45~4_combout ),
	.datac(\register[20][18]~q ),
	.datad(Selector8),
	.cin(gnd),
	.combout(\Mux45~5_combout ),
	.cout());
// synopsys translate_off
defparam \Mux45~5 .lut_mask = 16'hB8CC;
defparam \Mux45~5 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X66_Y39_N22
cycloneive_lcell_comb \Mux45~6 (
// Equation(s):
// \Mux45~6_combout  = (Selector10 & (((Selector91)))) # (!Selector10 & ((Selector91 & (\Mux45~3_combout )) # (!Selector91 & ((\Mux45~5_combout )))))

	.dataa(Selector10),
	.datab(\Mux45~3_combout ),
	.datac(\Mux45~5_combout ),
	.datad(Selector91),
	.cin(gnd),
	.combout(\Mux45~6_combout ),
	.cout());
// synopsys translate_off
defparam \Mux45~6 .lut_mask = 16'hEE50;
defparam \Mux45~6 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y36_N10
cycloneive_lcell_comb \register[25][18]~feeder (
// Equation(s):
// \register[25][18]~feeder_combout  = \register~77_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(\register~77_combout ),
	.datad(gnd),
	.cin(gnd),
	.combout(\register[25][18]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \register[25][18]~feeder .lut_mask = 16'hF0F0;
defparam \register[25][18]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X62_Y36_N11
dffeas \register[25][18] (
	.clk(!CLK),
	.d(\register[25][18]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~24_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\register[25][18]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \register[25][18] .is_wysiwyg = "true";
defparam \register[25][18] .power_up = "low";
// synopsys translate_on

// Location: FF_X63_Y33_N1
dffeas \register[29][18] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\register~77_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~28_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\register[29][18]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \register[29][18] .is_wysiwyg = "true";
defparam \register[29][18] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X62_Y34_N22
cycloneive_lcell_comb \register[17][18]~feeder (
// Equation(s):
// \register[17][18]~feeder_combout  = \register~77_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(\register~77_combout ),
	.datad(gnd),
	.cin(gnd),
	.combout(\register[17][18]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \register[17][18]~feeder .lut_mask = 16'hF0F0;
defparam \register[17][18]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X62_Y34_N23
dffeas \register[17][18] (
	.clk(!CLK),
	.d(\register[17][18]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~26_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\register[17][18]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \register[17][18] .is_wysiwyg = "true";
defparam \register[17][18] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X63_Y36_N12
cycloneive_lcell_comb \register[21][18]~feeder (
// Equation(s):
// \register[21][18]~feeder_combout  = \register~77_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(\register~77_combout ),
	.cin(gnd),
	.combout(\register[21][18]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \register[21][18]~feeder .lut_mask = 16'hFF00;
defparam \register[21][18]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X63_Y36_N13
dffeas \register[21][18] (
	.clk(!CLK),
	.d(\register[21][18]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~22_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\register[21][18]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \register[21][18] .is_wysiwyg = "true";
defparam \register[21][18] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X62_Y34_N0
cycloneive_lcell_comb \Mux45~0 (
// Equation(s):
// \Mux45~0_combout  = (Selector7 & (Selector8)) # (!Selector7 & ((Selector8 & ((\register[21][18]~q ))) # (!Selector8 & (\register[17][18]~q ))))

	.dataa(Selector7),
	.datab(Selector8),
	.datac(\register[17][18]~q ),
	.datad(\register[21][18]~q ),
	.cin(gnd),
	.combout(\Mux45~0_combout ),
	.cout());
// synopsys translate_off
defparam \Mux45~0 .lut_mask = 16'hDC98;
defparam \Mux45~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X63_Y33_N0
cycloneive_lcell_comb \Mux45~1 (
// Equation(s):
// \Mux45~1_combout  = (Selector7 & ((\Mux45~0_combout  & ((\register[29][18]~q ))) # (!\Mux45~0_combout  & (\register[25][18]~q )))) # (!Selector7 & (((\Mux45~0_combout ))))

	.dataa(\register[25][18]~q ),
	.datab(Selector7),
	.datac(\register[29][18]~q ),
	.datad(\Mux45~0_combout ),
	.cin(gnd),
	.combout(\Mux45~1_combout ),
	.cout());
// synopsys translate_off
defparam \Mux45~1 .lut_mask = 16'hF388;
defparam \Mux45~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y38_N30
cycloneive_lcell_comb \register[27][18]~feeder (
// Equation(s):
// \register[27][18]~feeder_combout  = \register~77_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(\register~77_combout ),
	.datad(gnd),
	.cin(gnd),
	.combout(\register[27][18]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \register[27][18]~feeder .lut_mask = 16'hF0F0;
defparam \register[27][18]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X60_Y38_N31
dffeas \register[27][18] (
	.clk(!CLK),
	.d(\register[27][18]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~38_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\register[27][18]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \register[27][18] .is_wysiwyg = "true";
defparam \register[27][18] .power_up = "low";
// synopsys translate_on

// Location: FF_X62_Y34_N27
dffeas \register[31][18] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\register~77_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~40_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\register[31][18]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \register[31][18] .is_wysiwyg = "true";
defparam \register[31][18] .power_up = "low";
// synopsys translate_on

// Location: FF_X62_Y38_N21
dffeas \register[23][18] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\register~77_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~37_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\register[23][18]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \register[23][18] .is_wysiwyg = "true";
defparam \register[23][18] .power_up = "low";
// synopsys translate_on

// Location: FF_X60_Y38_N5
dffeas \register[19][18] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\register~77_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~39_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\register[19][18]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \register[19][18] .is_wysiwyg = "true";
defparam \register[19][18] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X62_Y38_N20
cycloneive_lcell_comb \Mux45~7 (
// Equation(s):
// \Mux45~7_combout  = (Selector7 & (Selector8)) # (!Selector7 & ((Selector8 & (\register[23][18]~q )) # (!Selector8 & ((\register[19][18]~q )))))

	.dataa(Selector7),
	.datab(Selector8),
	.datac(\register[23][18]~q ),
	.datad(\register[19][18]~q ),
	.cin(gnd),
	.combout(\Mux45~7_combout ),
	.cout());
// synopsys translate_off
defparam \Mux45~7 .lut_mask = 16'hD9C8;
defparam \Mux45~7 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y34_N26
cycloneive_lcell_comb \Mux45~8 (
// Equation(s):
// \Mux45~8_combout  = (Selector7 & ((\Mux45~7_combout  & ((\register[31][18]~q ))) # (!\Mux45~7_combout  & (\register[27][18]~q )))) # (!Selector7 & (((\Mux45~7_combout ))))

	.dataa(Selector7),
	.datab(\register[27][18]~q ),
	.datac(\register[31][18]~q ),
	.datad(\Mux45~7_combout ),
	.cin(gnd),
	.combout(\Mux45~8_combout ),
	.cout());
// synopsys translate_off
defparam \Mux45~8 .lut_mask = 16'hF588;
defparam \Mux45~8 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X65_Y40_N4
cycloneive_lcell_comb \register[9][18]~feeder (
// Equation(s):
// \register[9][18]~feeder_combout  = \register~77_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(\register~77_combout ),
	.datad(gnd),
	.cin(gnd),
	.combout(\register[9][18]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \register[9][18]~feeder .lut_mask = 16'hF0F0;
defparam \register[9][18]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X65_Y40_N5
dffeas \register[9][18] (
	.clk(!CLK),
	.d(\register[9][18]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~44_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\register[9][18]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \register[9][18] .is_wysiwyg = "true";
defparam \register[9][18] .power_up = "low";
// synopsys translate_on

// Location: FF_X66_Y40_N5
dffeas \register[10][18] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\register~77_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~45_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\register[10][18]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \register[10][18] .is_wysiwyg = "true";
defparam \register[10][18] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X66_Y40_N4
cycloneive_lcell_comb \Mux45~10 (
// Equation(s):
// \Mux45~10_combout  = (Selector91 & (((\register[10][18]~q ) # (Selector10)))) # (!Selector91 & (\register[8][18]~q  & ((!Selector10))))

	.dataa(\register[8][18]~q ),
	.datab(Selector91),
	.datac(\register[10][18]~q ),
	.datad(Selector10),
	.cin(gnd),
	.combout(\Mux45~10_combout ),
	.cout());
// synopsys translate_off
defparam \Mux45~10 .lut_mask = 16'hCCE2;
defparam \Mux45~10 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X65_Y40_N23
dffeas \register[11][18] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\register~77_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~47_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\register[11][18]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \register[11][18] .is_wysiwyg = "true";
defparam \register[11][18] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X66_Y40_N20
cycloneive_lcell_comb \Mux45~11 (
// Equation(s):
// \Mux45~11_combout  = (Selector10 & ((\Mux45~10_combout  & ((\register[11][18]~q ))) # (!\Mux45~10_combout  & (\register[9][18]~q )))) # (!Selector10 & (((\Mux45~10_combout ))))

	.dataa(Selector10),
	.datab(\register[9][18]~q ),
	.datac(\Mux45~10_combout ),
	.datad(\register[11][18]~q ),
	.cin(gnd),
	.combout(\Mux45~11_combout ),
	.cout());
// synopsys translate_off
defparam \Mux45~11 .lut_mask = 16'hF858;
defparam \Mux45~11 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X60_Y36_N23
dffeas \register[12][18] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\register~77_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~52_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\register[12][18]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \register[12][18] .is_wysiwyg = "true";
defparam \register[12][18] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X60_Y36_N22
cycloneive_lcell_comb \Mux45~17 (
// Equation(s):
// \Mux45~17_combout  = (Selector10 & ((\register[13][18]~q ) # ((Selector91)))) # (!Selector10 & (((\register[12][18]~q  & !Selector91))))

	.dataa(\register[13][18]~q ),
	.datab(Selector10),
	.datac(\register[12][18]~q ),
	.datad(Selector91),
	.cin(gnd),
	.combout(\Mux45~17_combout ),
	.cout());
// synopsys translate_off
defparam \Mux45~17 .lut_mask = 16'hCCB8;
defparam \Mux45~17 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X60_Y36_N25
dffeas \register[14][18] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\register~77_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~61_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\register[14][18]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \register[14][18] .is_wysiwyg = "true";
defparam \register[14][18] .power_up = "low";
// synopsys translate_on

// Location: FF_X61_Y36_N17
dffeas \register[15][18] (
	.clk(!CLK),
	.d(\register~77_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~53_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\register[15][18]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \register[15][18] .is_wysiwyg = "true";
defparam \register[15][18] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X60_Y36_N24
cycloneive_lcell_comb \Mux45~18 (
// Equation(s):
// \Mux45~18_combout  = (\Mux45~17_combout  & (((\register[15][18]~q )) # (!Selector91))) # (!\Mux45~17_combout  & (Selector91 & (\register[14][18]~q )))

	.dataa(\Mux45~17_combout ),
	.datab(Selector91),
	.datac(\register[14][18]~q ),
	.datad(\register[15][18]~q ),
	.cin(gnd),
	.combout(\Mux45~18_combout ),
	.cout());
// synopsys translate_off
defparam \Mux45~18 .lut_mask = 16'hEA62;
defparam \Mux45~18 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X66_Y32_N19
dffeas \register[7][18] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\register~77_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~43_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\register[7][18]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \register[7][18] .is_wysiwyg = "true";
defparam \register[7][18] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X67_Y33_N0
cycloneive_lcell_comb \register[6][18]~feeder (
// Equation(s):
// \register[6][18]~feeder_combout  = \register~77_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(\register~77_combout ),
	.datad(gnd),
	.cin(gnd),
	.combout(\register[6][18]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \register[6][18]~feeder .lut_mask = 16'hF0F0;
defparam \register[6][18]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X67_Y33_N1
dffeas \register[6][18] (
	.clk(!CLK),
	.d(\register[6][18]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~58_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\register[6][18]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \register[6][18] .is_wysiwyg = "true";
defparam \register[6][18] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X66_Y32_N18
cycloneive_lcell_comb \Mux45~13 (
// Equation(s):
// \Mux45~13_combout  = (\Mux45~12_combout  & (((\register[7][18]~q )) # (!Selector91))) # (!\Mux45~12_combout  & (Selector91 & ((\register[6][18]~q ))))

	.dataa(\Mux45~12_combout ),
	.datab(Selector91),
	.datac(\register[7][18]~q ),
	.datad(\register[6][18]~q ),
	.cin(gnd),
	.combout(\Mux45~13_combout ),
	.cout());
// synopsys translate_off
defparam \Mux45~13 .lut_mask = 16'hE6A2;
defparam \Mux45~13 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X66_Y32_N21
dffeas \register[2][18] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\register~77_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~50_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\register[2][18]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \register[2][18] .is_wysiwyg = "true";
defparam \register[2][18] .power_up = "low";
// synopsys translate_on

// Location: FF_X65_Y33_N13
dffeas \register[3][18] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\register~77_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~48_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\register[3][18]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \register[3][18] .is_wysiwyg = "true";
defparam \register[3][18] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X65_Y33_N12
cycloneive_lcell_comb \Mux45~14 (
// Equation(s):
// \Mux45~14_combout  = (Selector10 & ((Selector91 & ((\register[3][18]~q ))) # (!Selector91 & (\register[1][18]~q ))))

	.dataa(\register[1][18]~q ),
	.datab(Selector91),
	.datac(\register[3][18]~q ),
	.datad(Selector10),
	.cin(gnd),
	.combout(\Mux45~14_combout ),
	.cout());
// synopsys translate_off
defparam \Mux45~14 .lut_mask = 16'hE200;
defparam \Mux45~14 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X66_Y32_N20
cycloneive_lcell_comb \Mux45~15 (
// Equation(s):
// \Mux45~15_combout  = (\Mux45~14_combout ) # ((!Selector10 & (Selector91 & \register[2][18]~q )))

	.dataa(Selector10),
	.datab(Selector91),
	.datac(\register[2][18]~q ),
	.datad(\Mux45~14_combout ),
	.cin(gnd),
	.combout(\Mux45~15_combout ),
	.cout());
// synopsys translate_off
defparam \Mux45~15 .lut_mask = 16'hFF40;
defparam \Mux45~15 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X66_Y39_N2
cycloneive_lcell_comb \Mux45~16 (
// Equation(s):
// \Mux45~16_combout  = (Selector7 & (Selector8)) # (!Selector7 & ((Selector8 & (\Mux45~13_combout )) # (!Selector8 & ((\Mux45~15_combout )))))

	.dataa(Selector7),
	.datab(Selector8),
	.datac(\Mux45~13_combout ),
	.datad(\Mux45~15_combout ),
	.cin(gnd),
	.combout(\Mux45~16_combout ),
	.cout());
// synopsys translate_off
defparam \Mux45~16 .lut_mask = 16'hD9C8;
defparam \Mux45~16 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y36_N2
cycloneive_lcell_comb \register~78 (
// Equation(s):
// \register~78_combout  = (WideOr01 & ((\wdat[17]~28_combout ) # ((plif_memwbregsrc_l_1 & plif_memwbrtnaddr_l_17))))

	.dataa(plif_memwbregsrc_l_1),
	.datab(plif_memwbrtnaddr_l_17),
	.datac(wdat_17),
	.datad(WideOr0),
	.cin(gnd),
	.combout(\register~78_combout ),
	.cout());
// synopsys translate_off
defparam \register~78 .lut_mask = 16'hF800;
defparam \register~78 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X68_Y39_N3
dffeas \register[30][17] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\register~78_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~56_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\register[30][17]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \register[30][17] .is_wysiwyg = "true";
defparam \register[30][17] .power_up = "low";
// synopsys translate_on

// Location: FF_X69_Y39_N29
dffeas \register[18][17] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\register~78_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~33_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\register[18][17]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \register[18][17] .is_wysiwyg = "true";
defparam \register[18][17] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X69_Y39_N28
cycloneive_lcell_comb \Mux46~2 (
// Equation(s):
// \Mux46~2_combout  = (Selector7 & (((Selector8)))) # (!Selector7 & ((Selector8 & (\register[22][17]~q )) # (!Selector8 & ((\register[18][17]~q )))))

	.dataa(\register[22][17]~q ),
	.datab(Selector7),
	.datac(\register[18][17]~q ),
	.datad(Selector8),
	.cin(gnd),
	.combout(\Mux46~2_combout ),
	.cout());
// synopsys translate_off
defparam \Mux46~2 .lut_mask = 16'hEE30;
defparam \Mux46~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X68_Y39_N2
cycloneive_lcell_comb \Mux46~3 (
// Equation(s):
// \Mux46~3_combout  = (Selector7 & ((\Mux46~2_combout  & ((\register[30][17]~q ))) # (!\Mux46~2_combout  & (\register[26][17]~q )))) # (!Selector7 & (((\Mux46~2_combout ))))

	.dataa(\register[26][17]~q ),
	.datab(Selector7),
	.datac(\register[30][17]~q ),
	.datad(\Mux46~2_combout ),
	.cin(gnd),
	.combout(\Mux46~3_combout ),
	.cout());
// synopsys translate_off
defparam \Mux46~3 .lut_mask = 16'hF388;
defparam \Mux46~3 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X61_Y40_N17
dffeas \register[24][17] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\register~78_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~34_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\register[24][17]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \register[24][17] .is_wysiwyg = "true";
defparam \register[24][17] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X69_Y38_N18
cycloneive_lcell_comb \register[16][17]~feeder (
// Equation(s):
// \register[16][17]~feeder_combout  = \register~78_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(\register~78_combout ),
	.datad(gnd),
	.cin(gnd),
	.combout(\register[16][17]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \register[16][17]~feeder .lut_mask = 16'hF0F0;
defparam \register[16][17]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X69_Y38_N19
dffeas \register[16][17] (
	.clk(!CLK),
	.d(\register[16][17]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~36_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\register[16][17]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \register[16][17] .is_wysiwyg = "true";
defparam \register[16][17] .power_up = "low";
// synopsys translate_on

// Location: FF_X69_Y38_N17
dffeas \register[20][17] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\register~78_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~35_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\register[20][17]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \register[20][17] .is_wysiwyg = "true";
defparam \register[20][17] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X69_Y38_N16
cycloneive_lcell_comb \Mux46~4 (
// Equation(s):
// \Mux46~4_combout  = (Selector8 & (((\register[20][17]~q ) # (Selector7)))) # (!Selector8 & (\register[16][17]~q  & ((!Selector7))))

	.dataa(Selector8),
	.datab(\register[16][17]~q ),
	.datac(\register[20][17]~q ),
	.datad(Selector7),
	.cin(gnd),
	.combout(\Mux46~4_combout ),
	.cout());
// synopsys translate_off
defparam \Mux46~4 .lut_mask = 16'hAAE4;
defparam \Mux46~4 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X67_Y40_N16
cycloneive_lcell_comb \Mux46~5 (
// Equation(s):
// \Mux46~5_combout  = (Selector7 & ((\Mux46~4_combout  & (\register[28][17]~q )) # (!\Mux46~4_combout  & ((\register[24][17]~q ))))) # (!Selector7 & (((\Mux46~4_combout ))))

	.dataa(\register[28][17]~q ),
	.datab(Selector7),
	.datac(\register[24][17]~q ),
	.datad(\Mux46~4_combout ),
	.cin(gnd),
	.combout(\Mux46~5_combout ),
	.cout());
// synopsys translate_off
defparam \Mux46~5 .lut_mask = 16'hBBC0;
defparam \Mux46~5 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X67_Y40_N18
cycloneive_lcell_comb \Mux46~6 (
// Equation(s):
// \Mux46~6_combout  = (Selector91 & ((\Mux46~3_combout ) # ((Selector10)))) # (!Selector91 & (((!Selector10 & \Mux46~5_combout ))))

	.dataa(\Mux46~3_combout ),
	.datab(Selector91),
	.datac(Selector10),
	.datad(\Mux46~5_combout ),
	.cin(gnd),
	.combout(\Mux46~6_combout ),
	.cout());
// synopsys translate_off
defparam \Mux46~6 .lut_mask = 16'hCBC8;
defparam \Mux46~6 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X67_Y40_N4
cycloneive_lcell_comb \register[31][17]~feeder (
// Equation(s):
// \register[31][17]~feeder_combout  = \register~78_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(\register~78_combout ),
	.cin(gnd),
	.combout(\register[31][17]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \register[31][17]~feeder .lut_mask = 16'hFF00;
defparam \register[31][17]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X67_Y40_N5
dffeas \register[31][17] (
	.clk(!CLK),
	.d(\register[31][17]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~40_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\register[31][17]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \register[31][17] .is_wysiwyg = "true";
defparam \register[31][17] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X65_Y32_N6
cycloneive_lcell_comb \register[23][17]~feeder (
// Equation(s):
// \register[23][17]~feeder_combout  = \register~78_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(\register~78_combout ),
	.datad(gnd),
	.cin(gnd),
	.combout(\register[23][17]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \register[23][17]~feeder .lut_mask = 16'hF0F0;
defparam \register[23][17]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X65_Y32_N7
dffeas \register[23][17] (
	.clk(!CLK),
	.d(\register[23][17]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~37_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\register[23][17]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \register[23][17] .is_wysiwyg = "true";
defparam \register[23][17] .power_up = "low";
// synopsys translate_on

// Location: FF_X62_Y39_N29
dffeas \register[27][17] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\register~78_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~38_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\register[27][17]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \register[27][17] .is_wysiwyg = "true";
defparam \register[27][17] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X62_Y39_N28
cycloneive_lcell_comb \Mux46~7 (
// Equation(s):
// \Mux46~7_combout  = (Selector8 & (((Selector7)))) # (!Selector8 & ((Selector7 & ((\register[27][17]~q ))) # (!Selector7 & (\register[19][17]~q ))))

	.dataa(\register[19][17]~q ),
	.datab(Selector8),
	.datac(\register[27][17]~q ),
	.datad(Selector7),
	.cin(gnd),
	.combout(\Mux46~7_combout ),
	.cout());
// synopsys translate_off
defparam \Mux46~7 .lut_mask = 16'hFC22;
defparam \Mux46~7 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X67_Y40_N30
cycloneive_lcell_comb \Mux46~8 (
// Equation(s):
// \Mux46~8_combout  = (Selector8 & ((\Mux46~7_combout  & (\register[31][17]~q )) # (!\Mux46~7_combout  & ((\register[23][17]~q ))))) # (!Selector8 & (((\Mux46~7_combout ))))

	.dataa(Selector8),
	.datab(\register[31][17]~q ),
	.datac(\register[23][17]~q ),
	.datad(\Mux46~7_combout ),
	.cin(gnd),
	.combout(\Mux46~8_combout ),
	.cout());
// synopsys translate_off
defparam \Mux46~8 .lut_mask = 16'hDDA0;
defparam \Mux46~8 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X63_Y34_N7
dffeas \register[21][17] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\register~78_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~22_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\register[21][17]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \register[21][17] .is_wysiwyg = "true";
defparam \register[21][17] .power_up = "low";
// synopsys translate_on

// Location: FF_X60_Y37_N1
dffeas \register[17][17] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\register~78_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~26_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\register[17][17]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \register[17][17] .is_wysiwyg = "true";
defparam \register[17][17] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X56_Y40_N12
cycloneive_lcell_comb \register[25][17]~feeder (
// Equation(s):
// \register[25][17]~feeder_combout  = \register~78_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(\register~78_combout ),
	.datad(gnd),
	.cin(gnd),
	.combout(\register[25][17]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \register[25][17]~feeder .lut_mask = 16'hF0F0;
defparam \register[25][17]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X56_Y40_N13
dffeas \register[25][17] (
	.clk(!CLK),
	.d(\register[25][17]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~24_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\register[25][17]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \register[25][17] .is_wysiwyg = "true";
defparam \register[25][17] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X60_Y37_N0
cycloneive_lcell_comb \Mux46~0 (
// Equation(s):
// \Mux46~0_combout  = (Selector8 & (Selector7)) # (!Selector8 & ((Selector7 & ((\register[25][17]~q ))) # (!Selector7 & (\register[17][17]~q ))))

	.dataa(Selector8),
	.datab(Selector7),
	.datac(\register[17][17]~q ),
	.datad(\register[25][17]~q ),
	.cin(gnd),
	.combout(\Mux46~0_combout ),
	.cout());
// synopsys translate_off
defparam \Mux46~0 .lut_mask = 16'hDC98;
defparam \Mux46~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y34_N28
cycloneive_lcell_comb \register[29][17]~feeder (
// Equation(s):
// \register[29][17]~feeder_combout  = \register~78_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(\register~78_combout ),
	.datad(gnd),
	.cin(gnd),
	.combout(\register[29][17]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \register[29][17]~feeder .lut_mask = 16'hF0F0;
defparam \register[29][17]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X61_Y34_N29
dffeas \register[29][17] (
	.clk(!CLK),
	.d(\register[29][17]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~28_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\register[29][17]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \register[29][17] .is_wysiwyg = "true";
defparam \register[29][17] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X61_Y34_N2
cycloneive_lcell_comb \Mux46~1 (
// Equation(s):
// \Mux46~1_combout  = (Selector8 & ((\Mux46~0_combout  & ((\register[29][17]~q ))) # (!\Mux46~0_combout  & (\register[21][17]~q )))) # (!Selector8 & (((\Mux46~0_combout ))))

	.dataa(Selector8),
	.datab(\register[21][17]~q ),
	.datac(\Mux46~0_combout ),
	.datad(\register[29][17]~q ),
	.cin(gnd),
	.combout(\Mux46~1_combout ),
	.cout());
// synopsys translate_off
defparam \Mux46~1 .lut_mask = 16'hF858;
defparam \Mux46~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X68_Y32_N15
dffeas \register[7][17] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\register~78_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~43_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\register[7][17]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \register[7][17] .is_wysiwyg = "true";
defparam \register[7][17] .power_up = "low";
// synopsys translate_on

// Location: FF_X68_Y32_N13
dffeas \register[6][17] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\register~78_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~58_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\register[6][17]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \register[6][17] .is_wysiwyg = "true";
defparam \register[6][17] .power_up = "low";
// synopsys translate_on

// Location: FF_X67_Y32_N11
dffeas \register[4][17] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\register~78_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~60_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\register[4][17]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \register[4][17] .is_wysiwyg = "true";
defparam \register[4][17] .power_up = "low";
// synopsys translate_on

// Location: FF_X67_Y32_N21
dffeas \register[5][17] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\register~78_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~59_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\register[5][17]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \register[5][17] .is_wysiwyg = "true";
defparam \register[5][17] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X67_Y32_N10
cycloneive_lcell_comb \Mux46~10 (
// Equation(s):
// \Mux46~10_combout  = (Selector10 & ((Selector91) # ((\register[5][17]~q )))) # (!Selector10 & (!Selector91 & (\register[4][17]~q )))

	.dataa(Selector10),
	.datab(Selector91),
	.datac(\register[4][17]~q ),
	.datad(\register[5][17]~q ),
	.cin(gnd),
	.combout(\Mux46~10_combout ),
	.cout());
// synopsys translate_off
defparam \Mux46~10 .lut_mask = 16'hBA98;
defparam \Mux46~10 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X68_Y32_N12
cycloneive_lcell_comb \Mux46~11 (
// Equation(s):
// \Mux46~11_combout  = (Selector91 & ((\Mux46~10_combout  & (\register[7][17]~q )) # (!\Mux46~10_combout  & ((\register[6][17]~q ))))) # (!Selector91 & (((\Mux46~10_combout ))))

	.dataa(Selector91),
	.datab(\register[7][17]~q ),
	.datac(\register[6][17]~q ),
	.datad(\Mux46~10_combout ),
	.cin(gnd),
	.combout(\Mux46~11_combout ),
	.cout());
// synopsys translate_off
defparam \Mux46~11 .lut_mask = 16'hDDA0;
defparam \Mux46~11 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X61_Y36_N3
dffeas \register[15][17] (
	.clk(!CLK),
	.d(\register~78_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~53_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\register[15][17]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \register[15][17] .is_wysiwyg = "true";
defparam \register[15][17] .power_up = "low";
// synopsys translate_on

// Location: FF_X60_Y36_N21
dffeas \register[14][17] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\register~78_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~61_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\register[14][17]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \register[14][17] .is_wysiwyg = "true";
defparam \register[14][17] .power_up = "low";
// synopsys translate_on

// Location: FF_X60_Y36_N11
dffeas \register[12][17] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\register~78_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~52_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\register[12][17]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \register[12][17] .is_wysiwyg = "true";
defparam \register[12][17] .power_up = "low";
// synopsys translate_on

// Location: FF_X59_Y36_N19
dffeas \register[13][17] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\register~78_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~62_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\register[13][17]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \register[13][17] .is_wysiwyg = "true";
defparam \register[13][17] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X60_Y36_N10
cycloneive_lcell_comb \Mux46~17 (
// Equation(s):
// \Mux46~17_combout  = (Selector91 & (Selector10)) # (!Selector91 & ((Selector10 & ((\register[13][17]~q ))) # (!Selector10 & (\register[12][17]~q ))))

	.dataa(Selector91),
	.datab(Selector10),
	.datac(\register[12][17]~q ),
	.datad(\register[13][17]~q ),
	.cin(gnd),
	.combout(\Mux46~17_combout ),
	.cout());
// synopsys translate_off
defparam \Mux46~17 .lut_mask = 16'hDC98;
defparam \Mux46~17 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y36_N20
cycloneive_lcell_comb \Mux46~18 (
// Equation(s):
// \Mux46~18_combout  = (Selector91 & ((\Mux46~17_combout  & (\register[15][17]~q )) # (!\Mux46~17_combout  & ((\register[14][17]~q ))))) # (!Selector91 & (((\Mux46~17_combout ))))

	.dataa(\register[15][17]~q ),
	.datab(Selector91),
	.datac(\register[14][17]~q ),
	.datad(\Mux46~17_combout ),
	.cin(gnd),
	.combout(\Mux46~18_combout ),
	.cout());
// synopsys translate_off
defparam \Mux46~18 .lut_mask = 16'hBBC0;
defparam \Mux46~18 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X63_Y40_N1
dffeas \register[9][17] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\register~78_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~44_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\register[9][17]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \register[9][17] .is_wysiwyg = "true";
defparam \register[9][17] .power_up = "low";
// synopsys translate_on

// Location: FF_X63_Y40_N15
dffeas \register[11][17] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\register~78_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~47_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\register[11][17]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \register[11][17] .is_wysiwyg = "true";
defparam \register[11][17] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X63_Y40_N14
cycloneive_lcell_comb \Mux46~13 (
// Equation(s):
// \Mux46~13_combout  = (\Mux46~12_combout  & (((\register[11][17]~q ) # (!Selector10)))) # (!\Mux46~12_combout  & (\register[9][17]~q  & ((Selector10))))

	.dataa(\Mux46~12_combout ),
	.datab(\register[9][17]~q ),
	.datac(\register[11][17]~q ),
	.datad(Selector10),
	.cin(gnd),
	.combout(\Mux46~13_combout ),
	.cout());
// synopsys translate_off
defparam \Mux46~13 .lut_mask = 16'hE4AA;
defparam \Mux46~13 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X69_Y33_N7
dffeas \register[1][17] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\register~78_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~49_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\register[1][17]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \register[1][17] .is_wysiwyg = "true";
defparam \register[1][17] .power_up = "low";
// synopsys translate_on

// Location: FF_X69_Y33_N13
dffeas \register[3][17] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\register~78_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~48_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\register[3][17]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \register[3][17] .is_wysiwyg = "true";
defparam \register[3][17] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X69_Y33_N6
cycloneive_lcell_comb \Mux46~14 (
// Equation(s):
// \Mux46~14_combout  = (Selector9 & ((plif_ifidinstr_l_17 & ((\register[3][17]~q ))) # (!plif_ifidinstr_l_17 & (\register[1][17]~q )))) # (!Selector9 & (((\register[1][17]~q ))))

	.dataa(Selector9),
	.datab(plif_ifidinstr_l_17),
	.datac(\register[1][17]~q ),
	.datad(\register[3][17]~q ),
	.cin(gnd),
	.combout(\Mux46~14_combout ),
	.cout());
// synopsys translate_off
defparam \Mux46~14 .lut_mask = 16'hF870;
defparam \Mux46~14 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X66_Y32_N6
cycloneive_lcell_comb \register[2][17]~feeder (
// Equation(s):
// \register[2][17]~feeder_combout  = \register~78_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(\register~78_combout ),
	.cin(gnd),
	.combout(\register[2][17]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \register[2][17]~feeder .lut_mask = 16'hFF00;
defparam \register[2][17]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X66_Y32_N7
dffeas \register[2][17] (
	.clk(!CLK),
	.d(\register[2][17]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~50_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\register[2][17]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \register[2][17] .is_wysiwyg = "true";
defparam \register[2][17] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X67_Y40_N6
cycloneive_lcell_comb \Mux46~15 (
// Equation(s):
// \Mux46~15_combout  = (Selector10 & (\Mux46~14_combout )) # (!Selector10 & (((Selector91 & \register[2][17]~q ))))

	.dataa(Selector10),
	.datab(\Mux46~14_combout ),
	.datac(Selector91),
	.datad(\register[2][17]~q ),
	.cin(gnd),
	.combout(\Mux46~15_combout ),
	.cout());
// synopsys translate_off
defparam \Mux46~15 .lut_mask = 16'hD888;
defparam \Mux46~15 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X67_Y40_N0
cycloneive_lcell_comb \Mux46~16 (
// Equation(s):
// \Mux46~16_combout  = (Selector8 & (Selector7)) # (!Selector8 & ((Selector7 & (\Mux46~13_combout )) # (!Selector7 & ((\Mux46~15_combout )))))

	.dataa(Selector8),
	.datab(Selector7),
	.datac(\Mux46~13_combout ),
	.datad(\Mux46~15_combout ),
	.cin(gnd),
	.combout(\Mux46~16_combout ),
	.cout());
// synopsys translate_off
defparam \Mux46~16 .lut_mask = 16'hD9C8;
defparam \Mux46~16 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y36_N10
cycloneive_lcell_comb \register~79 (
// Equation(s):
// \register~79_combout  = (WideOr01 & ((\wdat[16]~30_combout ) # ((plif_memwbrtnaddr_l_16 & plif_memwbregsrc_l_1))))

	.dataa(wdat_16),
	.datab(plif_memwbrtnaddr_l_16),
	.datac(plif_memwbregsrc_l_1),
	.datad(WideOr0),
	.cin(gnd),
	.combout(\register~79_combout ),
	.cout());
// synopsys translate_off
defparam \register~79 .lut_mask = 16'hEA00;
defparam \register~79 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X63_Y35_N10
cycloneive_lcell_comb \register[27][16]~feeder (
// Equation(s):
// \register[27][16]~feeder_combout  = \register~79_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(\register~79_combout ),
	.datad(gnd),
	.cin(gnd),
	.combout(\register[27][16]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \register[27][16]~feeder .lut_mask = 16'hF0F0;
defparam \register[27][16]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X63_Y35_N11
dffeas \register[27][16] (
	.clk(!CLK),
	.d(\register[27][16]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~38_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\register[27][16]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \register[27][16] .is_wysiwyg = "true";
defparam \register[27][16] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X67_Y40_N22
cycloneive_lcell_comb \register[31][16]~feeder (
// Equation(s):
// \register[31][16]~feeder_combout  = \register~79_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(\register~79_combout ),
	.cin(gnd),
	.combout(\register[31][16]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \register[31][16]~feeder .lut_mask = 16'hFF00;
defparam \register[31][16]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X67_Y40_N23
dffeas \register[31][16] (
	.clk(!CLK),
	.d(\register[31][16]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~40_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\register[31][16]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \register[31][16] .is_wysiwyg = "true";
defparam \register[31][16] .power_up = "low";
// synopsys translate_on

// Location: FF_X62_Y31_N21
dffeas \register[23][16] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\register~79_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~37_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\register[23][16]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \register[23][16] .is_wysiwyg = "true";
defparam \register[23][16] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X62_Y31_N20
cycloneive_lcell_comb \Mux47~7 (
// Equation(s):
// \Mux47~7_combout  = (Selector7 & (((Selector8)))) # (!Selector7 & ((Selector8 & ((\register[23][16]~q ))) # (!Selector8 & (\register[19][16]~q ))))

	.dataa(\register[19][16]~q ),
	.datab(Selector7),
	.datac(\register[23][16]~q ),
	.datad(Selector8),
	.cin(gnd),
	.combout(\Mux47~7_combout ),
	.cout());
// synopsys translate_off
defparam \Mux47~7 .lut_mask = 16'hFC22;
defparam \Mux47~7 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X67_Y40_N28
cycloneive_lcell_comb \Mux47~8 (
// Equation(s):
// \Mux47~8_combout  = (Selector7 & ((\Mux47~7_combout  & ((\register[31][16]~q ))) # (!\Mux47~7_combout  & (\register[27][16]~q )))) # (!Selector7 & (((\Mux47~7_combout ))))

	.dataa(\register[27][16]~q ),
	.datab(Selector7),
	.datac(\register[31][16]~q ),
	.datad(\Mux47~7_combout ),
	.cin(gnd),
	.combout(\Mux47~8_combout ),
	.cout());
// synopsys translate_off
defparam \Mux47~8 .lut_mask = 16'hF388;
defparam \Mux47~8 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X67_Y37_N21
dffeas \register[22][16] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\register~79_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~55_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\register[22][16]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \register[22][16] .is_wysiwyg = "true";
defparam \register[22][16] .power_up = "low";
// synopsys translate_on

// Location: FF_X68_Y37_N19
dffeas \register[30][16] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\register~79_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~56_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\register[30][16]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \register[30][16] .is_wysiwyg = "true";
defparam \register[30][16] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X68_Y37_N18
cycloneive_lcell_comb \Mux47~3 (
// Equation(s):
// \Mux47~3_combout  = (\Mux47~2_combout  & (((\register[30][16]~q ) # (!Selector8)))) # (!\Mux47~2_combout  & (\register[22][16]~q  & ((Selector8))))

	.dataa(\Mux47~2_combout ),
	.datab(\register[22][16]~q ),
	.datac(\register[30][16]~q ),
	.datad(Selector8),
	.cin(gnd),
	.combout(\Mux47~3_combout ),
	.cout());
// synopsys translate_off
defparam \Mux47~3 .lut_mask = 16'hE4AA;
defparam \Mux47~3 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X65_Y37_N17
dffeas \register[20][16] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\register~79_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~35_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\register[20][16]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \register[20][16] .is_wysiwyg = "true";
defparam \register[20][16] .power_up = "low";
// synopsys translate_on

// Location: FF_X68_Y34_N1
dffeas \register[28][16] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\register~79_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~57_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\register[28][16]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \register[28][16] .is_wysiwyg = "true";
defparam \register[28][16] .power_up = "low";
// synopsys translate_on

// Location: FF_X61_Y37_N17
dffeas \register[24][16] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\register~79_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~34_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\register[24][16]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \register[24][16] .is_wysiwyg = "true";
defparam \register[24][16] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X65_Y37_N2
cycloneive_lcell_comb \register[16][16]~feeder (
// Equation(s):
// \register[16][16]~feeder_combout  = \register~79_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(\register~79_combout ),
	.datad(gnd),
	.cin(gnd),
	.combout(\register[16][16]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \register[16][16]~feeder .lut_mask = 16'hF0F0;
defparam \register[16][16]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X65_Y37_N3
dffeas \register[16][16] (
	.clk(!CLK),
	.d(\register[16][16]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~36_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\register[16][16]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \register[16][16] .is_wysiwyg = "true";
defparam \register[16][16] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X61_Y37_N16
cycloneive_lcell_comb \Mux47~4 (
// Equation(s):
// \Mux47~4_combout  = (Selector7 & ((Selector8) # ((\register[24][16]~q )))) # (!Selector7 & (!Selector8 & ((\register[16][16]~q ))))

	.dataa(Selector7),
	.datab(Selector8),
	.datac(\register[24][16]~q ),
	.datad(\register[16][16]~q ),
	.cin(gnd),
	.combout(\Mux47~4_combout ),
	.cout());
// synopsys translate_off
defparam \Mux47~4 .lut_mask = 16'hB9A8;
defparam \Mux47~4 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X66_Y37_N26
cycloneive_lcell_comb \Mux47~5 (
// Equation(s):
// \Mux47~5_combout  = (Selector8 & ((\Mux47~4_combout  & ((\register[28][16]~q ))) # (!\Mux47~4_combout  & (\register[20][16]~q )))) # (!Selector8 & (((\Mux47~4_combout ))))

	.dataa(Selector8),
	.datab(\register[20][16]~q ),
	.datac(\register[28][16]~q ),
	.datad(\Mux47~4_combout ),
	.cin(gnd),
	.combout(\Mux47~5_combout ),
	.cout());
// synopsys translate_off
defparam \Mux47~5 .lut_mask = 16'hF588;
defparam \Mux47~5 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X67_Y40_N8
cycloneive_lcell_comb \Mux47~6 (
// Equation(s):
// \Mux47~6_combout  = (Selector91 & ((\Mux47~3_combout ) # ((Selector10)))) # (!Selector91 & (((!Selector10 & \Mux47~5_combout ))))

	.dataa(\Mux47~3_combout ),
	.datab(Selector91),
	.datac(Selector10),
	.datad(\Mux47~5_combout ),
	.cin(gnd),
	.combout(\Mux47~6_combout ),
	.cout());
// synopsys translate_off
defparam \Mux47~6 .lut_mask = 16'hCBC8;
defparam \Mux47~6 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X61_Y37_N27
dffeas \register[25][16] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\register~79_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~24_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\register[25][16]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \register[25][16] .is_wysiwyg = "true";
defparam \register[25][16] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X61_Y34_N4
cycloneive_lcell_comb \register[29][16]~feeder (
// Equation(s):
// \register[29][16]~feeder_combout  = \register~79_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(\register~79_combout ),
	.cin(gnd),
	.combout(\register[29][16]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \register[29][16]~feeder .lut_mask = 16'hFF00;
defparam \register[29][16]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X61_Y34_N5
dffeas \register[29][16] (
	.clk(!CLK),
	.d(\register[29][16]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~28_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\register[29][16]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \register[29][16] .is_wysiwyg = "true";
defparam \register[29][16] .power_up = "low";
// synopsys translate_on

// Location: FF_X60_Y37_N31
dffeas \register[17][16] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\register~79_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~26_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\register[17][16]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \register[17][16] .is_wysiwyg = "true";
defparam \register[17][16] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X60_Y37_N30
cycloneive_lcell_comb \Mux47~0 (
// Equation(s):
// \Mux47~0_combout  = (Selector7 & (((Selector8)))) # (!Selector7 & ((Selector8 & (\register[21][16]~q )) # (!Selector8 & ((\register[17][16]~q )))))

	.dataa(\register[21][16]~q ),
	.datab(Selector7),
	.datac(\register[17][16]~q ),
	.datad(Selector8),
	.cin(gnd),
	.combout(\Mux47~0_combout ),
	.cout());
// synopsys translate_off
defparam \Mux47~0 .lut_mask = 16'hEE30;
defparam \Mux47~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y34_N6
cycloneive_lcell_comb \Mux47~1 (
// Equation(s):
// \Mux47~1_combout  = (Selector7 & ((\Mux47~0_combout  & ((\register[29][16]~q ))) # (!\Mux47~0_combout  & (\register[25][16]~q )))) # (!Selector7 & (((\Mux47~0_combout ))))

	.dataa(Selector7),
	.datab(\register[25][16]~q ),
	.datac(\register[29][16]~q ),
	.datad(\Mux47~0_combout ),
	.cin(gnd),
	.combout(\Mux47~1_combout ),
	.cout());
// synopsys translate_off
defparam \Mux47~1 .lut_mask = 16'hF588;
defparam \Mux47~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X62_Y40_N5
dffeas \register[10][16] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\register~79_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~45_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\register[10][16]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \register[10][16] .is_wysiwyg = "true";
defparam \register[10][16] .power_up = "low";
// synopsys translate_on

// Location: FF_X62_Y40_N3
dffeas \register[8][16] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\register~79_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~46_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\register[8][16]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \register[8][16] .is_wysiwyg = "true";
defparam \register[8][16] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X62_Y40_N2
cycloneive_lcell_comb \Mux47~10 (
// Equation(s):
// \Mux47~10_combout  = (Selector91 & ((\register[10][16]~q ) # ((Selector10)))) # (!Selector91 & (((\register[8][16]~q  & !Selector10))))

	.dataa(Selector91),
	.datab(\register[10][16]~q ),
	.datac(\register[8][16]~q ),
	.datad(Selector10),
	.cin(gnd),
	.combout(\Mux47~10_combout ),
	.cout());
// synopsys translate_off
defparam \Mux47~10 .lut_mask = 16'hAAD8;
defparam \Mux47~10 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X63_Y40_N9
dffeas \register[9][16] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\register~79_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~44_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\register[9][16]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \register[9][16] .is_wysiwyg = "true";
defparam \register[9][16] .power_up = "low";
// synopsys translate_on

// Location: FF_X63_Y40_N31
dffeas \register[11][16] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\register~79_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~47_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\register[11][16]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \register[11][16] .is_wysiwyg = "true";
defparam \register[11][16] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X63_Y40_N30
cycloneive_lcell_comb \Mux47~11 (
// Equation(s):
// \Mux47~11_combout  = (\Mux47~10_combout  & (((\register[11][16]~q ) # (!Selector10)))) # (!\Mux47~10_combout  & (\register[9][16]~q  & ((Selector10))))

	.dataa(\Mux47~10_combout ),
	.datab(\register[9][16]~q ),
	.datac(\register[11][16]~q ),
	.datad(Selector10),
	.cin(gnd),
	.combout(\Mux47~11_combout ),
	.cout());
// synopsys translate_off
defparam \Mux47~11 .lut_mask = 16'hE4AA;
defparam \Mux47~11 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y36_N8
cycloneive_lcell_comb \register[15][16]~feeder (
// Equation(s):
// \register[15][16]~feeder_combout  = \register~79_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(\register~79_combout ),
	.cin(gnd),
	.combout(\register[15][16]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \register[15][16]~feeder .lut_mask = 16'hFF00;
defparam \register[15][16]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X61_Y36_N9
dffeas \register[15][16] (
	.clk(!CLK),
	.d(\register[15][16]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~53_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\register[15][16]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \register[15][16] .is_wysiwyg = "true";
defparam \register[15][16] .power_up = "low";
// synopsys translate_on

// Location: FF_X60_Y36_N5
dffeas \register[14][16] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\register~79_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~61_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\register[14][16]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \register[14][16] .is_wysiwyg = "true";
defparam \register[14][16] .power_up = "low";
// synopsys translate_on

// Location: FF_X60_Y36_N3
dffeas \register[12][16] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\register~79_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~52_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\register[12][16]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \register[12][16] .is_wysiwyg = "true";
defparam \register[12][16] .power_up = "low";
// synopsys translate_on

// Location: FF_X59_Y36_N29
dffeas \register[13][16] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\register~79_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~62_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\register[13][16]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \register[13][16] .is_wysiwyg = "true";
defparam \register[13][16] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X60_Y36_N2
cycloneive_lcell_comb \Mux47~17 (
// Equation(s):
// \Mux47~17_combout  = (Selector91 & (Selector10)) # (!Selector91 & ((Selector10 & ((\register[13][16]~q ))) # (!Selector10 & (\register[12][16]~q ))))

	.dataa(Selector91),
	.datab(Selector10),
	.datac(\register[12][16]~q ),
	.datad(\register[13][16]~q ),
	.cin(gnd),
	.combout(\Mux47~17_combout ),
	.cout());
// synopsys translate_off
defparam \Mux47~17 .lut_mask = 16'hDC98;
defparam \Mux47~17 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y36_N4
cycloneive_lcell_comb \Mux47~18 (
// Equation(s):
// \Mux47~18_combout  = (Selector91 & ((\Mux47~17_combout  & (\register[15][16]~q )) # (!\Mux47~17_combout  & ((\register[14][16]~q ))))) # (!Selector91 & (((\Mux47~17_combout ))))

	.dataa(Selector91),
	.datab(\register[15][16]~q ),
	.datac(\register[14][16]~q ),
	.datad(\Mux47~17_combout ),
	.cin(gnd),
	.combout(\Mux47~18_combout ),
	.cout());
// synopsys translate_off
defparam \Mux47~18 .lut_mask = 16'hDDA0;
defparam \Mux47~18 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X68_Y32_N17
dffeas \register[6][16] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\register~79_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~58_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\register[6][16]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \register[6][16] .is_wysiwyg = "true";
defparam \register[6][16] .power_up = "low";
// synopsys translate_on

// Location: FF_X68_Y32_N31
dffeas \register[7][16] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\register~79_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~43_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\register[7][16]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \register[7][16] .is_wysiwyg = "true";
defparam \register[7][16] .power_up = "low";
// synopsys translate_on

// Location: FF_X69_Y32_N7
dffeas \register[4][16] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\register~79_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~60_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\register[4][16]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \register[4][16] .is_wysiwyg = "true";
defparam \register[4][16] .power_up = "low";
// synopsys translate_on

// Location: FF_X69_Y32_N29
dffeas \register[5][16] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\register~79_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~59_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\register[5][16]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \register[5][16] .is_wysiwyg = "true";
defparam \register[5][16] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X69_Y32_N6
cycloneive_lcell_comb \Mux47~12 (
// Equation(s):
// \Mux47~12_combout  = (Selector10 & ((Selector91) # ((\register[5][16]~q )))) # (!Selector10 & (!Selector91 & (\register[4][16]~q )))

	.dataa(Selector10),
	.datab(Selector91),
	.datac(\register[4][16]~q ),
	.datad(\register[5][16]~q ),
	.cin(gnd),
	.combout(\Mux47~12_combout ),
	.cout());
// synopsys translate_off
defparam \Mux47~12 .lut_mask = 16'hBA98;
defparam \Mux47~12 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X68_Y32_N30
cycloneive_lcell_comb \Mux47~13 (
// Equation(s):
// \Mux47~13_combout  = (Selector91 & ((\Mux47~12_combout  & ((\register[7][16]~q ))) # (!\Mux47~12_combout  & (\register[6][16]~q )))) # (!Selector91 & (((\Mux47~12_combout ))))

	.dataa(Selector91),
	.datab(\register[6][16]~q ),
	.datac(\register[7][16]~q ),
	.datad(\Mux47~12_combout ),
	.cin(gnd),
	.combout(\Mux47~13_combout ),
	.cout());
// synopsys translate_off
defparam \Mux47~13 .lut_mask = 16'hF588;
defparam \Mux47~13 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X66_Y32_N5
dffeas \register[2][16] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\register~79_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~50_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\register[2][16]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \register[2][16] .is_wysiwyg = "true";
defparam \register[2][16] .power_up = "low";
// synopsys translate_on

// Location: FF_X70_Y34_N7
dffeas \register[1][16] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\register~79_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~49_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\register[1][16]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \register[1][16] .is_wysiwyg = "true";
defparam \register[1][16] .power_up = "low";
// synopsys translate_on

// Location: FF_X70_Y34_N1
dffeas \register[3][16] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\register~79_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~48_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\register[3][16]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \register[3][16] .is_wysiwyg = "true";
defparam \register[3][16] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X70_Y34_N6
cycloneive_lcell_comb \Mux47~14 (
// Equation(s):
// \Mux47~14_combout  = (Selector10 & ((Selector91 & ((\register[3][16]~q ))) # (!Selector91 & (\register[1][16]~q ))))

	.dataa(Selector10),
	.datab(Selector91),
	.datac(\register[1][16]~q ),
	.datad(\register[3][16]~q ),
	.cin(gnd),
	.combout(\Mux47~14_combout ),
	.cout());
// synopsys translate_off
defparam \Mux47~14 .lut_mask = 16'hA820;
defparam \Mux47~14 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X66_Y32_N4
cycloneive_lcell_comb \Mux47~15 (
// Equation(s):
// \Mux47~15_combout  = (\Mux47~14_combout ) # ((!Selector10 & (Selector91 & \register[2][16]~q )))

	.dataa(Selector10),
	.datab(Selector91),
	.datac(\register[2][16]~q ),
	.datad(\Mux47~14_combout ),
	.cin(gnd),
	.combout(\Mux47~15_combout ),
	.cout());
// synopsys translate_off
defparam \Mux47~15 .lut_mask = 16'hFF40;
defparam \Mux47~15 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X67_Y40_N12
cycloneive_lcell_comb \Mux47~16 (
// Equation(s):
// \Mux47~16_combout  = (Selector8 & ((Selector7) # ((\Mux47~13_combout )))) # (!Selector8 & (!Selector7 & ((\Mux47~15_combout ))))

	.dataa(Selector8),
	.datab(Selector7),
	.datac(\Mux47~13_combout ),
	.datad(\Mux47~15_combout ),
	.cin(gnd),
	.combout(\Mux47~16_combout ),
	.cout());
// synopsys translate_off
defparam \Mux47~16 .lut_mask = 16'hB9A8;
defparam \Mux47~16 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y36_N22
cycloneive_lcell_comb \register~80 (
// Equation(s):
// \register~80_combout  = (WideOr01 & ((\wdat[15]~32_combout ) # ((plif_memwbrtnaddr_l_15 & plif_memwbregsrc_l_1))))

	.dataa(plif_memwbrtnaddr_l_15),
	.datab(WideOr0),
	.datac(plif_memwbregsrc_l_1),
	.datad(wdat_15),
	.cin(gnd),
	.combout(\register~80_combout ),
	.cout());
// synopsys translate_off
defparam \register~80 .lut_mask = 16'hCC80;
defparam \register~80 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X69_Y36_N22
cycloneive_lcell_comb \register[28][15]~feeder (
// Equation(s):
// \register[28][15]~feeder_combout  = \register~80_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(\register~80_combout ),
	.cin(gnd),
	.combout(\register[28][15]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \register[28][15]~feeder .lut_mask = 16'hFF00;
defparam \register[28][15]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X69_Y36_N23
dffeas \register[28][15] (
	.clk(!CLK),
	.d(\register[28][15]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~57_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\register[28][15]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \register[28][15] .is_wysiwyg = "true";
defparam \register[28][15] .power_up = "low";
// synopsys translate_on

// Location: FF_X69_Y34_N5
dffeas \register[16][15] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\register~80_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~36_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\register[16][15]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \register[16][15] .is_wysiwyg = "true";
defparam \register[16][15] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X69_Y38_N4
cycloneive_lcell_comb \register[20][15]~feeder (
// Equation(s):
// \register[20][15]~feeder_combout  = \register~80_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(\register~80_combout ),
	.datad(gnd),
	.cin(gnd),
	.combout(\register[20][15]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \register[20][15]~feeder .lut_mask = 16'hF0F0;
defparam \register[20][15]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X69_Y38_N5
dffeas \register[20][15] (
	.clk(!CLK),
	.d(\register[20][15]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~35_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\register[20][15]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \register[20][15] .is_wysiwyg = "true";
defparam \register[20][15] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X69_Y34_N4
cycloneive_lcell_comb \Mux48~4 (
// Equation(s):
// \Mux48~4_combout  = (Selector7 & (Selector8)) # (!Selector7 & ((Selector8 & ((\register[20][15]~q ))) # (!Selector8 & (\register[16][15]~q ))))

	.dataa(Selector7),
	.datab(Selector8),
	.datac(\register[16][15]~q ),
	.datad(\register[20][15]~q ),
	.cin(gnd),
	.combout(\Mux48~4_combout ),
	.cout());
// synopsys translate_off
defparam \Mux48~4 .lut_mask = 16'hDC98;
defparam \Mux48~4 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X69_Y34_N18
cycloneive_lcell_comb \register[24][15]~feeder (
// Equation(s):
// \register[24][15]~feeder_combout  = \register~80_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(\register~80_combout ),
	.datad(gnd),
	.cin(gnd),
	.combout(\register[24][15]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \register[24][15]~feeder .lut_mask = 16'hF0F0;
defparam \register[24][15]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X69_Y34_N19
dffeas \register[24][15] (
	.clk(!CLK),
	.d(\register[24][15]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~34_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\register[24][15]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \register[24][15] .is_wysiwyg = "true";
defparam \register[24][15] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X69_Y34_N22
cycloneive_lcell_comb \Mux48~5 (
// Equation(s):
// \Mux48~5_combout  = (Selector7 & ((\Mux48~4_combout  & (\register[28][15]~q )) # (!\Mux48~4_combout  & ((\register[24][15]~q ))))) # (!Selector7 & (((\Mux48~4_combout ))))

	.dataa(Selector7),
	.datab(\register[28][15]~q ),
	.datac(\Mux48~4_combout ),
	.datad(\register[24][15]~q ),
	.cin(gnd),
	.combout(\Mux48~5_combout ),
	.cout());
// synopsys translate_off
defparam \Mux48~5 .lut_mask = 16'hDAD0;
defparam \Mux48~5 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X68_Y38_N25
dffeas \register[26][15] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\register~80_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~54_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\register[26][15]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \register[26][15] .is_wysiwyg = "true";
defparam \register[26][15] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X69_Y36_N4
cycloneive_lcell_comb \register[30][15]~feeder (
// Equation(s):
// \register[30][15]~feeder_combout  = \register~80_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(\register~80_combout ),
	.cin(gnd),
	.combout(\register[30][15]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \register[30][15]~feeder .lut_mask = 16'hFF00;
defparam \register[30][15]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X69_Y36_N5
dffeas \register[30][15] (
	.clk(!CLK),
	.d(\register[30][15]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~56_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\register[30][15]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \register[30][15] .is_wysiwyg = "true";
defparam \register[30][15] .power_up = "low";
// synopsys translate_on

// Location: FF_X68_Y38_N3
dffeas \register[18][15] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\register~80_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~33_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\register[18][15]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \register[18][15] .is_wysiwyg = "true";
defparam \register[18][15] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X69_Y37_N16
cycloneive_lcell_comb \register[22][15]~feeder (
// Equation(s):
// \register[22][15]~feeder_combout  = \register~80_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(\register~80_combout ),
	.cin(gnd),
	.combout(\register[22][15]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \register[22][15]~feeder .lut_mask = 16'hFF00;
defparam \register[22][15]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X69_Y37_N17
dffeas \register[22][15] (
	.clk(!CLK),
	.d(\register[22][15]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~55_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\register[22][15]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \register[22][15] .is_wysiwyg = "true";
defparam \register[22][15] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X68_Y38_N2
cycloneive_lcell_comb \Mux48~2 (
// Equation(s):
// \Mux48~2_combout  = (Selector7 & (Selector8)) # (!Selector7 & ((Selector8 & ((\register[22][15]~q ))) # (!Selector8 & (\register[18][15]~q ))))

	.dataa(Selector7),
	.datab(Selector8),
	.datac(\register[18][15]~q ),
	.datad(\register[22][15]~q ),
	.cin(gnd),
	.combout(\Mux48~2_combout ),
	.cout());
// synopsys translate_off
defparam \Mux48~2 .lut_mask = 16'hDC98;
defparam \Mux48~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X69_Y34_N28
cycloneive_lcell_comb \Mux48~3 (
// Equation(s):
// \Mux48~3_combout  = (Selector7 & ((\Mux48~2_combout  & ((\register[30][15]~q ))) # (!\Mux48~2_combout  & (\register[26][15]~q )))) # (!Selector7 & (((\Mux48~2_combout ))))

	.dataa(Selector7),
	.datab(\register[26][15]~q ),
	.datac(\register[30][15]~q ),
	.datad(\Mux48~2_combout ),
	.cin(gnd),
	.combout(\Mux48~3_combout ),
	.cout());
// synopsys translate_off
defparam \Mux48~3 .lut_mask = 16'hF588;
defparam \Mux48~3 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X69_Y34_N0
cycloneive_lcell_comb \Mux48~6 (
// Equation(s):
// \Mux48~6_combout  = (Selector91 & ((Selector10) # ((\Mux48~3_combout )))) # (!Selector91 & (!Selector10 & (\Mux48~5_combout )))

	.dataa(Selector91),
	.datab(Selector10),
	.datac(\Mux48~5_combout ),
	.datad(\Mux48~3_combout ),
	.cin(gnd),
	.combout(\Mux48~6_combout ),
	.cout());
// synopsys translate_off
defparam \Mux48~6 .lut_mask = 16'hBA98;
defparam \Mux48~6 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y31_N0
cycloneive_lcell_comb \register[23][15]~feeder (
// Equation(s):
// \register[23][15]~feeder_combout  = \register~80_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(\register~80_combout ),
	.datad(gnd),
	.cin(gnd),
	.combout(\register[23][15]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \register[23][15]~feeder .lut_mask = 16'hF0F0;
defparam \register[23][15]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X62_Y31_N1
dffeas \register[23][15] (
	.clk(!CLK),
	.d(\register[23][15]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~37_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\register[23][15]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \register[23][15] .is_wysiwyg = "true";
defparam \register[23][15] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X61_Y38_N2
cycloneive_lcell_comb \register[31][15]~feeder (
// Equation(s):
// \register[31][15]~feeder_combout  = \register~80_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(\register~80_combout ),
	.datad(gnd),
	.cin(gnd),
	.combout(\register[31][15]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \register[31][15]~feeder .lut_mask = 16'hF0F0;
defparam \register[31][15]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X61_Y38_N3
dffeas \register[31][15] (
	.clk(!CLK),
	.d(\register[31][15]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~40_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\register[31][15]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \register[31][15] .is_wysiwyg = "true";
defparam \register[31][15] .power_up = "low";
// synopsys translate_on

// Location: FF_X60_Y38_N1
dffeas \register[27][15] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\register~80_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~38_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\register[27][15]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \register[27][15] .is_wysiwyg = "true";
defparam \register[27][15] .power_up = "low";
// synopsys translate_on

// Location: FF_X62_Y31_N15
dffeas \register[19][15] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\register~80_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~39_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\register[19][15]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \register[19][15] .is_wysiwyg = "true";
defparam \register[19][15] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X60_Y38_N0
cycloneive_lcell_comb \Mux48~7 (
// Equation(s):
// \Mux48~7_combout  = (Selector8 & (Selector7)) # (!Selector8 & ((Selector7 & (\register[27][15]~q )) # (!Selector7 & ((\register[19][15]~q )))))

	.dataa(Selector8),
	.datab(Selector7),
	.datac(\register[27][15]~q ),
	.datad(\register[19][15]~q ),
	.cin(gnd),
	.combout(\Mux48~7_combout ),
	.cout());
// synopsys translate_off
defparam \Mux48~7 .lut_mask = 16'hD9C8;
defparam \Mux48~7 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y38_N8
cycloneive_lcell_comb \Mux48~8 (
// Equation(s):
// \Mux48~8_combout  = (\Mux48~7_combout  & (((\register[31][15]~q ) # (!Selector8)))) # (!\Mux48~7_combout  & (\register[23][15]~q  & ((Selector8))))

	.dataa(\register[23][15]~q ),
	.datab(\register[31][15]~q ),
	.datac(\Mux48~7_combout ),
	.datad(Selector8),
	.cin(gnd),
	.combout(\Mux48~8_combout ),
	.cout());
// synopsys translate_off
defparam \Mux48~8 .lut_mask = 16'hCAF0;
defparam \Mux48~8 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y31_N4
cycloneive_lcell_comb \register[29][15]~feeder (
// Equation(s):
// \register[29][15]~feeder_combout  = \register~80_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(\register~80_combout ),
	.cin(gnd),
	.combout(\register[29][15]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \register[29][15]~feeder .lut_mask = 16'hFF00;
defparam \register[29][15]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X61_Y31_N5
dffeas \register[29][15] (
	.clk(!CLK),
	.d(\register[29][15]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~28_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\register[29][15]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \register[29][15] .is_wysiwyg = "true";
defparam \register[29][15] .power_up = "low";
// synopsys translate_on

// Location: FF_X62_Y33_N7
dffeas \register[21][15] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\register~80_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~22_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\register[21][15]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \register[21][15] .is_wysiwyg = "true";
defparam \register[21][15] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X59_Y40_N28
cycloneive_lcell_comb \register[25][15]~feeder (
// Equation(s):
// \register[25][15]~feeder_combout  = \register~80_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(\register~80_combout ),
	.datad(gnd),
	.cin(gnd),
	.combout(\register[25][15]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \register[25][15]~feeder .lut_mask = 16'hF0F0;
defparam \register[25][15]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X59_Y40_N29
dffeas \register[25][15] (
	.clk(!CLK),
	.d(\register[25][15]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~24_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\register[25][15]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \register[25][15] .is_wysiwyg = "true";
defparam \register[25][15] .power_up = "low";
// synopsys translate_on

// Location: FF_X62_Y34_N29
dffeas \register[17][15] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\register~80_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~26_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\register[17][15]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \register[17][15] .is_wysiwyg = "true";
defparam \register[17][15] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X62_Y34_N28
cycloneive_lcell_comb \Mux48~0 (
// Equation(s):
// \Mux48~0_combout  = (Selector7 & ((\register[25][15]~q ) # ((Selector8)))) # (!Selector7 & (((\register[17][15]~q  & !Selector8))))

	.dataa(Selector7),
	.datab(\register[25][15]~q ),
	.datac(\register[17][15]~q ),
	.datad(Selector8),
	.cin(gnd),
	.combout(\Mux48~0_combout ),
	.cout());
// synopsys translate_off
defparam \Mux48~0 .lut_mask = 16'hAAD8;
defparam \Mux48~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y31_N18
cycloneive_lcell_comb \Mux48~1 (
// Equation(s):
// \Mux48~1_combout  = (Selector8 & ((\Mux48~0_combout  & (\register[29][15]~q )) # (!\Mux48~0_combout  & ((\register[21][15]~q ))))) # (!Selector8 & (((\Mux48~0_combout ))))

	.dataa(Selector8),
	.datab(\register[29][15]~q ),
	.datac(\register[21][15]~q ),
	.datad(\Mux48~0_combout ),
	.cin(gnd),
	.combout(\Mux48~1_combout ),
	.cout());
// synopsys translate_off
defparam \Mux48~1 .lut_mask = 16'hDDA0;
defparam \Mux48~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X68_Y32_N19
dffeas \register[7][15] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\register~80_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~43_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\register[7][15]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \register[7][15] .is_wysiwyg = "true";
defparam \register[7][15] .power_up = "low";
// synopsys translate_on

// Location: FF_X68_Y32_N9
dffeas \register[6][15] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\register~80_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~58_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\register[6][15]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \register[6][15] .is_wysiwyg = "true";
defparam \register[6][15] .power_up = "low";
// synopsys translate_on

// Location: FF_X69_Y32_N5
dffeas \register[5][15] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\register~80_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~59_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\register[5][15]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \register[5][15] .is_wysiwyg = "true";
defparam \register[5][15] .power_up = "low";
// synopsys translate_on

// Location: FF_X69_Y32_N3
dffeas \register[4][15] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\register~80_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~60_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\register[4][15]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \register[4][15] .is_wysiwyg = "true";
defparam \register[4][15] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X69_Y32_N2
cycloneive_lcell_comb \Mux48~10 (
// Equation(s):
// \Mux48~10_combout  = (Selector91 & (((Selector10)))) # (!Selector91 & ((Selector10 & (\register[5][15]~q )) # (!Selector10 & ((\register[4][15]~q )))))

	.dataa(Selector91),
	.datab(\register[5][15]~q ),
	.datac(\register[4][15]~q ),
	.datad(Selector10),
	.cin(gnd),
	.combout(\Mux48~10_combout ),
	.cout());
// synopsys translate_off
defparam \Mux48~10 .lut_mask = 16'hEE50;
defparam \Mux48~10 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X68_Y32_N8
cycloneive_lcell_comb \Mux48~11 (
// Equation(s):
// \Mux48~11_combout  = (Selector91 & ((\Mux48~10_combout  & (\register[7][15]~q )) # (!\Mux48~10_combout  & ((\register[6][15]~q ))))) # (!Selector91 & (((\Mux48~10_combout ))))

	.dataa(Selector91),
	.datab(\register[7][15]~q ),
	.datac(\register[6][15]~q ),
	.datad(\Mux48~10_combout ),
	.cin(gnd),
	.combout(\Mux48~11_combout ),
	.cout());
// synopsys translate_off
defparam \Mux48~11 .lut_mask = 16'hDDA0;
defparam \Mux48~11 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X62_Y33_N13
dffeas \register[14][15] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\register~80_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~61_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\register[14][15]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \register[14][15] .is_wysiwyg = "true";
defparam \register[14][15] .power_up = "low";
// synopsys translate_on

// Location: FF_X63_Y30_N3
dffeas \register[12][15] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\register~80_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~52_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\register[12][15]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \register[12][15] .is_wysiwyg = "true";
defparam \register[12][15] .power_up = "low";
// synopsys translate_on

// Location: FF_X63_Y30_N1
dffeas \register[13][15] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\register~80_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~62_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\register[13][15]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \register[13][15] .is_wysiwyg = "true";
defparam \register[13][15] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X63_Y30_N0
cycloneive_lcell_comb \Mux48~17 (
// Equation(s):
// \Mux48~17_combout  = (Selector91 & (((Selector10)))) # (!Selector91 & ((Selector10 & ((\register[13][15]~q ))) # (!Selector10 & (\register[12][15]~q ))))

	.dataa(Selector91),
	.datab(\register[12][15]~q ),
	.datac(\register[13][15]~q ),
	.datad(Selector10),
	.cin(gnd),
	.combout(\Mux48~17_combout ),
	.cout());
// synopsys translate_off
defparam \Mux48~17 .lut_mask = 16'hFA44;
defparam \Mux48~17 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X61_Y36_N23
dffeas \register[15][15] (
	.clk(!CLK),
	.d(\register~80_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~53_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\register[15][15]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \register[15][15] .is_wysiwyg = "true";
defparam \register[15][15] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X62_Y33_N30
cycloneive_lcell_comb \Mux48~18 (
// Equation(s):
// \Mux48~18_combout  = (Selector91 & ((\Mux48~17_combout  & ((\register[15][15]~q ))) # (!\Mux48~17_combout  & (\register[14][15]~q )))) # (!Selector91 & (((\Mux48~17_combout ))))

	.dataa(\register[14][15]~q ),
	.datab(Selector91),
	.datac(\Mux48~17_combout ),
	.datad(\register[15][15]~q ),
	.cin(gnd),
	.combout(\Mux48~18_combout ),
	.cout());
// synopsys translate_off
defparam \Mux48~18 .lut_mask = 16'hF838;
defparam \Mux48~18 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X65_Y33_N1
dffeas \register[3][15] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\register~80_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~48_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\register[3][15]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \register[3][15] .is_wysiwyg = "true";
defparam \register[3][15] .power_up = "low";
// synopsys translate_on

// Location: FF_X65_Y33_N23
dffeas \register[1][15] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\register~80_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~49_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\register[1][15]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \register[1][15] .is_wysiwyg = "true";
defparam \register[1][15] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X65_Y33_N22
cycloneive_lcell_comb \Mux48~14 (
// Equation(s):
// \Mux48~14_combout  = (Selector10 & ((Selector91 & (\register[3][15]~q )) # (!Selector91 & ((\register[1][15]~q )))))

	.dataa(Selector91),
	.datab(\register[3][15]~q ),
	.datac(\register[1][15]~q ),
	.datad(Selector10),
	.cin(gnd),
	.combout(\Mux48~14_combout ),
	.cout());
// synopsys translate_off
defparam \Mux48~14 .lut_mask = 16'hD800;
defparam \Mux48~14 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X69_Y34_N30
cycloneive_lcell_comb \Mux48~15 (
// Equation(s):
// \Mux48~15_combout  = (\Mux48~14_combout ) # ((\register[2][15]~q  & (Selector91 & !Selector10)))

	.dataa(\register[2][15]~q ),
	.datab(Selector91),
	.datac(Selector10),
	.datad(\Mux48~14_combout ),
	.cin(gnd),
	.combout(\Mux48~15_combout ),
	.cout());
// synopsys translate_off
defparam \Mux48~15 .lut_mask = 16'hFF08;
defparam \Mux48~15 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X63_Y40_N19
dffeas \register[11][15] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\register~80_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~47_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\register[11][15]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \register[11][15] .is_wysiwyg = "true";
defparam \register[11][15] .power_up = "low";
// synopsys translate_on

// Location: FF_X63_Y40_N29
dffeas \register[9][15] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\register~80_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~44_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\register[9][15]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \register[9][15] .is_wysiwyg = "true";
defparam \register[9][15] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X63_Y40_N18
cycloneive_lcell_comb \Mux48~13 (
// Equation(s):
// \Mux48~13_combout  = (\Mux48~12_combout  & (((\register[11][15]~q )) # (!Selector10))) # (!\Mux48~12_combout  & (Selector10 & ((\register[9][15]~q ))))

	.dataa(\Mux48~12_combout ),
	.datab(Selector10),
	.datac(\register[11][15]~q ),
	.datad(\register[9][15]~q ),
	.cin(gnd),
	.combout(\Mux48~13_combout ),
	.cout());
// synopsys translate_off
defparam \Mux48~13 .lut_mask = 16'hE6A2;
defparam \Mux48~13 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X70_Y35_N0
cycloneive_lcell_comb \Mux48~16 (
// Equation(s):
// \Mux48~16_combout  = (Selector8 & (Selector7)) # (!Selector8 & ((Selector7 & ((\Mux48~13_combout ))) # (!Selector7 & (\Mux48~15_combout ))))

	.dataa(Selector8),
	.datab(Selector7),
	.datac(\Mux48~15_combout ),
	.datad(\Mux48~13_combout ),
	.cin(gnd),
	.combout(\Mux48~16_combout ),
	.cout());
// synopsys translate_off
defparam \Mux48~16 .lut_mask = 16'hDC98;
defparam \Mux48~16 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y36_N20
cycloneive_lcell_comb \register~81 (
// Equation(s):
// \register~81_combout  = (WideOr01 & ((\wdat[14]~34_combout ) # ((plif_memwbrtnaddr_l_14 & plif_memwbregsrc_l_1))))

	.dataa(plif_memwbrtnaddr_l_14),
	.datab(wdat_14),
	.datac(plif_memwbregsrc_l_1),
	.datad(WideOr0),
	.cin(gnd),
	.combout(\register~81_combout ),
	.cout());
// synopsys translate_off
defparam \register~81 .lut_mask = 16'hEC00;
defparam \register~81 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X60_Y38_N11
dffeas \register[27][14] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\register~81_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~38_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\register[27][14]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \register[27][14] .is_wysiwyg = "true";
defparam \register[27][14] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X66_Y30_N18
cycloneive_lcell_comb \register[31][14]~feeder (
// Equation(s):
// \register[31][14]~feeder_combout  = \register~81_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(\register~81_combout ),
	.cin(gnd),
	.combout(\register[31][14]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \register[31][14]~feeder .lut_mask = 16'hFF00;
defparam \register[31][14]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X66_Y30_N19
dffeas \register[31][14] (
	.clk(!CLK),
	.d(\register[31][14]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~40_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\register[31][14]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \register[31][14] .is_wysiwyg = "true";
defparam \register[31][14] .power_up = "low";
// synopsys translate_on

// Location: FF_X60_Y35_N21
dffeas \register[23][14] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\register~81_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~37_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\register[23][14]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \register[23][14] .is_wysiwyg = "true";
defparam \register[23][14] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X60_Y35_N20
cycloneive_lcell_comb \Mux49~7 (
// Equation(s):
// \Mux49~7_combout  = (Selector7 & (((Selector8)))) # (!Selector7 & ((Selector8 & ((\register[23][14]~q ))) # (!Selector8 & (\register[19][14]~q ))))

	.dataa(\register[19][14]~q ),
	.datab(Selector7),
	.datac(\register[23][14]~q ),
	.datad(Selector8),
	.cin(gnd),
	.combout(\Mux49~7_combout ),
	.cout());
// synopsys translate_off
defparam \Mux49~7 .lut_mask = 16'hFC22;
defparam \Mux49~7 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X66_Y30_N8
cycloneive_lcell_comb \Mux49~8 (
// Equation(s):
// \Mux49~8_combout  = (Selector7 & ((\Mux49~7_combout  & ((\register[31][14]~q ))) # (!\Mux49~7_combout  & (\register[27][14]~q )))) # (!Selector7 & (((\Mux49~7_combout ))))

	.dataa(\register[27][14]~q ),
	.datab(\register[31][14]~q ),
	.datac(Selector7),
	.datad(\Mux49~7_combout ),
	.cin(gnd),
	.combout(\Mux49~8_combout ),
	.cout());
// synopsys translate_off
defparam \Mux49~8 .lut_mask = 16'hCFA0;
defparam \Mux49~8 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X60_Y34_N3
dffeas \register[25][14] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\register~81_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~24_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\register[25][14]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \register[25][14] .is_wysiwyg = "true";
defparam \register[25][14] .power_up = "low";
// synopsys translate_on

// Location: FF_X61_Y34_N9
dffeas \register[29][14] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\register~81_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~28_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\register[29][14]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \register[29][14] .is_wysiwyg = "true";
defparam \register[29][14] .power_up = "low";
// synopsys translate_on

// Location: FF_X60_Y37_N29
dffeas \register[17][14] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\register~81_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~26_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\register[17][14]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \register[17][14] .is_wysiwyg = "true";
defparam \register[17][14] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X63_Y34_N12
cycloneive_lcell_comb \register[21][14]~feeder (
// Equation(s):
// \register[21][14]~feeder_combout  = \register~81_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(\register~81_combout ),
	.datad(gnd),
	.cin(gnd),
	.combout(\register[21][14]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \register[21][14]~feeder .lut_mask = 16'hF0F0;
defparam \register[21][14]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X63_Y34_N13
dffeas \register[21][14] (
	.clk(!CLK),
	.d(\register[21][14]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~22_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\register[21][14]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \register[21][14] .is_wysiwyg = "true";
defparam \register[21][14] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X60_Y37_N28
cycloneive_lcell_comb \Mux49~0 (
// Equation(s):
// \Mux49~0_combout  = (Selector8 & ((Selector7) # ((\register[21][14]~q )))) # (!Selector8 & (!Selector7 & (\register[17][14]~q )))

	.dataa(Selector8),
	.datab(Selector7),
	.datac(\register[17][14]~q ),
	.datad(\register[21][14]~q ),
	.cin(gnd),
	.combout(\Mux49~0_combout ),
	.cout());
// synopsys translate_off
defparam \Mux49~0 .lut_mask = 16'hBA98;
defparam \Mux49~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y34_N8
cycloneive_lcell_comb \Mux49~1 (
// Equation(s):
// \Mux49~1_combout  = (Selector7 & ((\Mux49~0_combout  & ((\register[29][14]~q ))) # (!\Mux49~0_combout  & (\register[25][14]~q )))) # (!Selector7 & (((\Mux49~0_combout ))))

	.dataa(\register[25][14]~q ),
	.datab(Selector7),
	.datac(\register[29][14]~q ),
	.datad(\Mux49~0_combout ),
	.cin(gnd),
	.combout(\Mux49~1_combout ),
	.cout());
// synopsys translate_off
defparam \Mux49~1 .lut_mask = 16'hF388;
defparam \Mux49~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X68_Y39_N13
dffeas \register[30][14] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\register~81_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~56_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\register[30][14]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \register[30][14] .is_wysiwyg = "true";
defparam \register[30][14] .power_up = "low";
// synopsys translate_on

// Location: FF_X68_Y35_N5
dffeas \register[26][14] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\register~81_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~54_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\register[26][14]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \register[26][14] .is_wysiwyg = "true";
defparam \register[26][14] .power_up = "low";
// synopsys translate_on

// Location: FF_X69_Y35_N3
dffeas \register[18][14] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\register~81_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~33_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\register[18][14]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \register[18][14] .is_wysiwyg = "true";
defparam \register[18][14] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X69_Y35_N2
cycloneive_lcell_comb \Mux49~2 (
// Equation(s):
// \Mux49~2_combout  = (Selector7 & ((\register[26][14]~q ) # ((Selector8)))) # (!Selector7 & (((\register[18][14]~q  & !Selector8))))

	.dataa(Selector7),
	.datab(\register[26][14]~q ),
	.datac(\register[18][14]~q ),
	.datad(Selector8),
	.cin(gnd),
	.combout(\Mux49~2_combout ),
	.cout());
// synopsys translate_off
defparam \Mux49~2 .lut_mask = 16'hAAD8;
defparam \Mux49~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X68_Y39_N12
cycloneive_lcell_comb \Mux49~3 (
// Equation(s):
// \Mux49~3_combout  = (Selector8 & ((\Mux49~2_combout  & ((\register[30][14]~q ))) # (!\Mux49~2_combout  & (\register[22][14]~q )))) # (!Selector8 & (((\Mux49~2_combout ))))

	.dataa(\register[22][14]~q ),
	.datab(Selector8),
	.datac(\register[30][14]~q ),
	.datad(\Mux49~2_combout ),
	.cin(gnd),
	.combout(\Mux49~3_combout ),
	.cout());
// synopsys translate_off
defparam \Mux49~3 .lut_mask = 16'hF388;
defparam \Mux49~3 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X65_Y37_N5
dffeas \register[20][14] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\register~81_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~35_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\register[20][14]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \register[20][14] .is_wysiwyg = "true";
defparam \register[20][14] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X68_Y34_N30
cycloneive_lcell_comb \register[28][14]~feeder (
// Equation(s):
// \register[28][14]~feeder_combout  = \register~81_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(\register~81_combout ),
	.cin(gnd),
	.combout(\register[28][14]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \register[28][14]~feeder .lut_mask = 16'hFF00;
defparam \register[28][14]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X68_Y34_N31
dffeas \register[28][14] (
	.clk(!CLK),
	.d(\register[28][14]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~57_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\register[28][14]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \register[28][14] .is_wysiwyg = "true";
defparam \register[28][14] .power_up = "low";
// synopsys translate_on

// Location: FF_X61_Y37_N3
dffeas \register[24][14] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\register~81_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~34_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\register[24][14]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \register[24][14] .is_wysiwyg = "true";
defparam \register[24][14] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X65_Y37_N18
cycloneive_lcell_comb \register[16][14]~feeder (
// Equation(s):
// \register[16][14]~feeder_combout  = \register~81_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(\register~81_combout ),
	.datad(gnd),
	.cin(gnd),
	.combout(\register[16][14]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \register[16][14]~feeder .lut_mask = 16'hF0F0;
defparam \register[16][14]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X65_Y37_N19
dffeas \register[16][14] (
	.clk(!CLK),
	.d(\register[16][14]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~36_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\register[16][14]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \register[16][14] .is_wysiwyg = "true";
defparam \register[16][14] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X61_Y37_N2
cycloneive_lcell_comb \Mux49~4 (
// Equation(s):
// \Mux49~4_combout  = (Selector7 & ((Selector8) # ((\register[24][14]~q )))) # (!Selector7 & (!Selector8 & ((\register[16][14]~q ))))

	.dataa(Selector7),
	.datab(Selector8),
	.datac(\register[24][14]~q ),
	.datad(\register[16][14]~q ),
	.cin(gnd),
	.combout(\Mux49~4_combout ),
	.cout());
// synopsys translate_off
defparam \Mux49~4 .lut_mask = 16'hB9A8;
defparam \Mux49~4 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X65_Y37_N12
cycloneive_lcell_comb \Mux49~5 (
// Equation(s):
// \Mux49~5_combout  = (Selector8 & ((\Mux49~4_combout  & ((\register[28][14]~q ))) # (!\Mux49~4_combout  & (\register[20][14]~q )))) # (!Selector8 & (((\Mux49~4_combout ))))

	.dataa(Selector8),
	.datab(\register[20][14]~q ),
	.datac(\register[28][14]~q ),
	.datad(\Mux49~4_combout ),
	.cin(gnd),
	.combout(\Mux49~5_combout ),
	.cout());
// synopsys translate_off
defparam \Mux49~5 .lut_mask = 16'hF588;
defparam \Mux49~5 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X66_Y30_N24
cycloneive_lcell_comb \Mux49~6 (
// Equation(s):
// \Mux49~6_combout  = (Selector91 & ((Selector10) # ((\Mux49~3_combout )))) # (!Selector91 & (!Selector10 & ((\Mux49~5_combout ))))

	.dataa(Selector91),
	.datab(Selector10),
	.datac(\Mux49~3_combout ),
	.datad(\Mux49~5_combout ),
	.cin(gnd),
	.combout(\Mux49~6_combout ),
	.cout());
// synopsys translate_off
defparam \Mux49~6 .lut_mask = 16'hB9A8;
defparam \Mux49~6 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X66_Y34_N15
dffeas \register[2][14] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\register~81_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~50_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\register[2][14]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \register[2][14] .is_wysiwyg = "true";
defparam \register[2][14] .power_up = "low";
// synopsys translate_on

// Location: FF_X70_Y34_N15
dffeas \register[1][14] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\register~81_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~49_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\register[1][14]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \register[1][14] .is_wysiwyg = "true";
defparam \register[1][14] .power_up = "low";
// synopsys translate_on

// Location: FF_X70_Y34_N17
dffeas \register[3][14] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\register~81_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~48_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\register[3][14]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \register[3][14] .is_wysiwyg = "true";
defparam \register[3][14] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X70_Y34_N14
cycloneive_lcell_comb \Mux49~14 (
// Equation(s):
// \Mux49~14_combout  = (Selector10 & ((Selector91 & ((\register[3][14]~q ))) # (!Selector91 & (\register[1][14]~q ))))

	.dataa(Selector10),
	.datab(Selector91),
	.datac(\register[1][14]~q ),
	.datad(\register[3][14]~q ),
	.cin(gnd),
	.combout(\Mux49~14_combout ),
	.cout());
// synopsys translate_off
defparam \Mux49~14 .lut_mask = 16'hA820;
defparam \Mux49~14 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X66_Y30_N0
cycloneive_lcell_comb \Mux49~15 (
// Equation(s):
// \Mux49~15_combout  = (\Mux49~14_combout ) # ((Selector91 & (\register[2][14]~q  & !Selector10)))

	.dataa(Selector91),
	.datab(\register[2][14]~q ),
	.datac(\Mux49~14_combout ),
	.datad(Selector10),
	.cin(gnd),
	.combout(\Mux49~15_combout ),
	.cout());
// synopsys translate_off
defparam \Mux49~15 .lut_mask = 16'hF0F8;
defparam \Mux49~15 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X69_Y32_N25
dffeas \register[5][14] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\register~81_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~59_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\register[5][14]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \register[5][14] .is_wysiwyg = "true";
defparam \register[5][14] .power_up = "low";
// synopsys translate_on

// Location: FF_X69_Y32_N15
dffeas \register[4][14] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\register~81_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~60_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\register[4][14]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \register[4][14] .is_wysiwyg = "true";
defparam \register[4][14] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X69_Y32_N14
cycloneive_lcell_comb \Mux49~12 (
// Equation(s):
// \Mux49~12_combout  = (Selector10 & ((\register[5][14]~q ) # ((Selector91)))) # (!Selector10 & (((\register[4][14]~q  & !Selector91))))

	.dataa(Selector10),
	.datab(\register[5][14]~q ),
	.datac(\register[4][14]~q ),
	.datad(Selector91),
	.cin(gnd),
	.combout(\Mux49~12_combout ),
	.cout());
// synopsys translate_off
defparam \Mux49~12 .lut_mask = 16'hAAD8;
defparam \Mux49~12 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X68_Y32_N7
dffeas \register[7][14] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\register~81_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~43_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\register[7][14]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \register[7][14] .is_wysiwyg = "true";
defparam \register[7][14] .power_up = "low";
// synopsys translate_on

// Location: FF_X68_Y32_N21
dffeas \register[6][14] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\register~81_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~58_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\register[6][14]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \register[6][14] .is_wysiwyg = "true";
defparam \register[6][14] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X68_Y32_N6
cycloneive_lcell_comb \Mux49~13 (
// Equation(s):
// \Mux49~13_combout  = (Selector91 & ((\Mux49~12_combout  & (\register[7][14]~q )) # (!\Mux49~12_combout  & ((\register[6][14]~q ))))) # (!Selector91 & (\Mux49~12_combout ))

	.dataa(Selector91),
	.datab(\Mux49~12_combout ),
	.datac(\register[7][14]~q ),
	.datad(\register[6][14]~q ),
	.cin(gnd),
	.combout(\Mux49~13_combout ),
	.cout());
// synopsys translate_off
defparam \Mux49~13 .lut_mask = 16'hE6C4;
defparam \Mux49~13 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X66_Y30_N6
cycloneive_lcell_comb \Mux49~16 (
// Equation(s):
// \Mux49~16_combout  = (Selector8 & (((Selector7) # (\Mux49~13_combout )))) # (!Selector8 & (\Mux49~15_combout  & (!Selector7)))

	.dataa(Selector8),
	.datab(\Mux49~15_combout ),
	.datac(Selector7),
	.datad(\Mux49~13_combout ),
	.cin(gnd),
	.combout(\Mux49~16_combout ),
	.cout());
// synopsys translate_off
defparam \Mux49~16 .lut_mask = 16'hAEA4;
defparam \Mux49~16 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X63_Y34_N10
cycloneive_lcell_comb \register[9][14]~feeder (
// Equation(s):
// \register[9][14]~feeder_combout  = \register~81_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(\register~81_combout ),
	.datad(gnd),
	.cin(gnd),
	.combout(\register[9][14]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \register[9][14]~feeder .lut_mask = 16'hF0F0;
defparam \register[9][14]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X63_Y34_N11
dffeas \register[9][14] (
	.clk(!CLK),
	.d(\register[9][14]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~44_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\register[9][14]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \register[9][14] .is_wysiwyg = "true";
defparam \register[9][14] .power_up = "low";
// synopsys translate_on

// Location: FF_X66_Y34_N29
dffeas \register[11][14] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\register~81_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~47_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\register[11][14]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \register[11][14] .is_wysiwyg = "true";
defparam \register[11][14] .power_up = "low";
// synopsys translate_on

// Location: FF_X62_Y40_N21
dffeas \register[10][14] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\register~81_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~45_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\register[10][14]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \register[10][14] .is_wysiwyg = "true";
defparam \register[10][14] .power_up = "low";
// synopsys translate_on

// Location: FF_X62_Y40_N23
dffeas \register[8][14] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\register~81_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~46_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\register[8][14]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \register[8][14] .is_wysiwyg = "true";
defparam \register[8][14] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X62_Y40_N22
cycloneive_lcell_comb \Mux49~10 (
// Equation(s):
// \Mux49~10_combout  = (Selector91 & ((\register[10][14]~q ) # ((Selector10)))) # (!Selector91 & (((\register[8][14]~q  & !Selector10))))

	.dataa(Selector91),
	.datab(\register[10][14]~q ),
	.datac(\register[8][14]~q ),
	.datad(Selector10),
	.cin(gnd),
	.combout(\Mux49~10_combout ),
	.cout());
// synopsys translate_off
defparam \Mux49~10 .lut_mask = 16'hAAD8;
defparam \Mux49~10 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X63_Y34_N20
cycloneive_lcell_comb \Mux49~11 (
// Equation(s):
// \Mux49~11_combout  = (Selector10 & ((\Mux49~10_combout  & ((\register[11][14]~q ))) # (!\Mux49~10_combout  & (\register[9][14]~q )))) # (!Selector10 & (((\Mux49~10_combout ))))

	.dataa(\register[9][14]~q ),
	.datab(Selector10),
	.datac(\register[11][14]~q ),
	.datad(\Mux49~10_combout ),
	.cin(gnd),
	.combout(\Mux49~11_combout ),
	.cout());
// synopsys translate_off
defparam \Mux49~11 .lut_mask = 16'hF388;
defparam \Mux49~11 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X60_Y34_N9
dffeas \register[14][14] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\register~81_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~61_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\register[14][14]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \register[14][14] .is_wysiwyg = "true";
defparam \register[14][14] .power_up = "low";
// synopsys translate_on

// Location: FF_X61_Y36_N21
dffeas \register[15][14] (
	.clk(!CLK),
	.d(\register~81_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~53_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\register[15][14]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \register[15][14] .is_wysiwyg = "true";
defparam \register[15][14] .power_up = "low";
// synopsys translate_on

// Location: FF_X63_Y30_N21
dffeas \register[13][14] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\register~81_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~62_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\register[13][14]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \register[13][14] .is_wysiwyg = "true";
defparam \register[13][14] .power_up = "low";
// synopsys translate_on

// Location: FF_X63_Y30_N31
dffeas \register[12][14] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\register~81_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~52_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\register[12][14]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \register[12][14] .is_wysiwyg = "true";
defparam \register[12][14] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X63_Y30_N30
cycloneive_lcell_comb \Mux49~17 (
// Equation(s):
// \Mux49~17_combout  = (Selector91 & (((Selector10)))) # (!Selector91 & ((Selector10 & (\register[13][14]~q )) # (!Selector10 & ((\register[12][14]~q )))))

	.dataa(Selector91),
	.datab(\register[13][14]~q ),
	.datac(\register[12][14]~q ),
	.datad(Selector10),
	.cin(gnd),
	.combout(\Mux49~17_combout ),
	.cout());
// synopsys translate_off
defparam \Mux49~17 .lut_mask = 16'hEE50;
defparam \Mux49~17 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X66_Y30_N28
cycloneive_lcell_comb \Mux49~18 (
// Equation(s):
// \Mux49~18_combout  = (Selector91 & ((\Mux49~17_combout  & ((\register[15][14]~q ))) # (!\Mux49~17_combout  & (\register[14][14]~q )))) # (!Selector91 & (((\Mux49~17_combout ))))

	.dataa(Selector91),
	.datab(\register[14][14]~q ),
	.datac(\register[15][14]~q ),
	.datad(\Mux49~17_combout ),
	.cin(gnd),
	.combout(\Mux49~18_combout ),
	.cout());
// synopsys translate_off
defparam \Mux49~18 .lut_mask = 16'hF588;
defparam \Mux49~18 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y36_N26
cycloneive_lcell_comb \register~82 (
// Equation(s):
// \register~82_combout  = (WideOr01 & ((\wdat[13]~36_combout ) # ((plif_memwbrtnaddr_l_13 & plif_memwbregsrc_l_1))))

	.dataa(plif_memwbrtnaddr_l_13),
	.datab(WideOr0),
	.datac(plif_memwbregsrc_l_1),
	.datad(wdat_13),
	.cin(gnd),
	.combout(\register~82_combout ),
	.cout());
// synopsys translate_off
defparam \register~82 .lut_mask = 16'hCC80;
defparam \register~82 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y38_N22
cycloneive_lcell_comb \register[29][13]~feeder (
// Equation(s):
// \register[29][13]~feeder_combout  = \register~82_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(\register~82_combout ),
	.datad(gnd),
	.cin(gnd),
	.combout(\register[29][13]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \register[29][13]~feeder .lut_mask = 16'hF0F0;
defparam \register[29][13]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X61_Y38_N23
dffeas \register[29][13] (
	.clk(!CLK),
	.d(\register[29][13]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~28_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\register[29][13]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \register[29][13] .is_wysiwyg = "true";
defparam \register[29][13] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X62_Y33_N16
cycloneive_lcell_comb \register[21][13]~feeder (
// Equation(s):
// \register[21][13]~feeder_combout  = \register~82_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(\register~82_combout ),
	.datad(gnd),
	.cin(gnd),
	.combout(\register[21][13]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \register[21][13]~feeder .lut_mask = 16'hF0F0;
defparam \register[21][13]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X62_Y33_N17
dffeas \register[21][13] (
	.clk(!CLK),
	.d(\register[21][13]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~22_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\register[21][13]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \register[21][13] .is_wysiwyg = "true";
defparam \register[21][13] .power_up = "low";
// synopsys translate_on

// Location: FF_X60_Y37_N19
dffeas \register[17][13] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\register~82_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~26_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\register[17][13]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \register[17][13] .is_wysiwyg = "true";
defparam \register[17][13] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X60_Y37_N18
cycloneive_lcell_comb \Mux50~0 (
// Equation(s):
// \Mux50~0_combout  = (Selector7 & ((\register[25][13]~q ) # ((Selector8)))) # (!Selector7 & (((\register[17][13]~q  & !Selector8))))

	.dataa(\register[25][13]~q ),
	.datab(Selector7),
	.datac(\register[17][13]~q ),
	.datad(Selector8),
	.cin(gnd),
	.combout(\Mux50~0_combout ),
	.cout());
// synopsys translate_off
defparam \Mux50~0 .lut_mask = 16'hCCB8;
defparam \Mux50~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y38_N20
cycloneive_lcell_comb \Mux50~1 (
// Equation(s):
// \Mux50~1_combout  = (\Mux50~0_combout  & ((\register[29][13]~q ) # ((!Selector8)))) # (!\Mux50~0_combout  & (((\register[21][13]~q  & Selector8))))

	.dataa(\register[29][13]~q ),
	.datab(\register[21][13]~q ),
	.datac(\Mux50~0_combout ),
	.datad(Selector8),
	.cin(gnd),
	.combout(\Mux50~1_combout ),
	.cout());
// synopsys translate_off
defparam \Mux50~1 .lut_mask = 16'hACF0;
defparam \Mux50~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y40_N26
cycloneive_lcell_comb \register[23][13]~feeder (
// Equation(s):
// \register[23][13]~feeder_combout  = \register~82_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(\register~82_combout ),
	.cin(gnd),
	.combout(\register[23][13]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \register[23][13]~feeder .lut_mask = 16'hFF00;
defparam \register[23][13]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X60_Y40_N27
dffeas \register[23][13] (
	.clk(!CLK),
	.d(\register[23][13]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~37_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\register[23][13]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \register[23][13] .is_wysiwyg = "true";
defparam \register[23][13] .power_up = "low";
// synopsys translate_on

// Location: FF_X61_Y38_N7
dffeas \register[31][13] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\register~82_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~40_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\register[31][13]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \register[31][13] .is_wysiwyg = "true";
defparam \register[31][13] .power_up = "low";
// synopsys translate_on

// Location: FF_X60_Y38_N19
dffeas \register[27][13] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\register~82_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~38_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\register[27][13]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \register[27][13] .is_wysiwyg = "true";
defparam \register[27][13] .power_up = "low";
// synopsys translate_on

// Location: FF_X60_Y38_N29
dffeas \register[19][13] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\register~82_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~39_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\register[19][13]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \register[19][13] .is_wysiwyg = "true";
defparam \register[19][13] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X60_Y38_N18
cycloneive_lcell_comb \Mux50~7 (
// Equation(s):
// \Mux50~7_combout  = (Selector8 & (Selector7)) # (!Selector8 & ((Selector7 & (\register[27][13]~q )) # (!Selector7 & ((\register[19][13]~q )))))

	.dataa(Selector8),
	.datab(Selector7),
	.datac(\register[27][13]~q ),
	.datad(\register[19][13]~q ),
	.cin(gnd),
	.combout(\Mux50~7_combout ),
	.cout());
// synopsys translate_off
defparam \Mux50~7 .lut_mask = 16'hD9C8;
defparam \Mux50~7 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y38_N6
cycloneive_lcell_comb \Mux50~8 (
// Equation(s):
// \Mux50~8_combout  = (Selector8 & ((\Mux50~7_combout  & ((\register[31][13]~q ))) # (!\Mux50~7_combout  & (\register[23][13]~q )))) # (!Selector8 & (((\Mux50~7_combout ))))

	.dataa(\register[23][13]~q ),
	.datab(Selector8),
	.datac(\register[31][13]~q ),
	.datad(\Mux50~7_combout ),
	.cin(gnd),
	.combout(\Mux50~8_combout ),
	.cout());
// synopsys translate_off
defparam \Mux50~8 .lut_mask = 16'hF388;
defparam \Mux50~8 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X65_Y38_N24
cycloneive_lcell_comb \register[24][13]~feeder (
// Equation(s):
// \register[24][13]~feeder_combout  = \register~82_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(\register~82_combout ),
	.datad(gnd),
	.cin(gnd),
	.combout(\register[24][13]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \register[24][13]~feeder .lut_mask = 16'hF0F0;
defparam \register[24][13]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X65_Y38_N25
dffeas \register[24][13] (
	.clk(!CLK),
	.d(\register[24][13]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~34_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\register[24][13]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \register[24][13] .is_wysiwyg = "true";
defparam \register[24][13] .power_up = "low";
// synopsys translate_on

// Location: FF_X65_Y34_N19
dffeas \register[20][13] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\register~82_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~35_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\register[20][13]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \register[20][13] .is_wysiwyg = "true";
defparam \register[20][13] .power_up = "low";
// synopsys translate_on

// Location: FF_X65_Y34_N25
dffeas \register[16][13] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\register~82_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~36_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\register[16][13]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \register[16][13] .is_wysiwyg = "true";
defparam \register[16][13] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X65_Y34_N18
cycloneive_lcell_comb \Mux50~4 (
// Equation(s):
// \Mux50~4_combout  = (Selector7 & (Selector8)) # (!Selector7 & ((Selector8 & (\register[20][13]~q )) # (!Selector8 & ((\register[16][13]~q )))))

	.dataa(Selector7),
	.datab(Selector8),
	.datac(\register[20][13]~q ),
	.datad(\register[16][13]~q ),
	.cin(gnd),
	.combout(\Mux50~4_combout ),
	.cout());
// synopsys translate_off
defparam \Mux50~4 .lut_mask = 16'hD9C8;
defparam \Mux50~4 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X65_Y38_N20
cycloneive_lcell_comb \Mux50~5 (
// Equation(s):
// \Mux50~5_combout  = (\Mux50~4_combout  & ((\register[28][13]~q ) # ((!Selector7)))) # (!\Mux50~4_combout  & (((\register[24][13]~q  & Selector7))))

	.dataa(\register[28][13]~q ),
	.datab(\register[24][13]~q ),
	.datac(\Mux50~4_combout ),
	.datad(Selector7),
	.cin(gnd),
	.combout(\Mux50~5_combout ),
	.cout());
// synopsys translate_off
defparam \Mux50~5 .lut_mask = 16'hACF0;
defparam \Mux50~5 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X68_Y38_N1
dffeas \register[26][13] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\register~82_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~54_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\register[26][13]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \register[26][13] .is_wysiwyg = "true";
defparam \register[26][13] .power_up = "low";
// synopsys translate_on

// Location: FF_X68_Y39_N29
dffeas \register[30][13] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\register~82_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~56_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\register[30][13]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \register[30][13] .is_wysiwyg = "true";
defparam \register[30][13] .power_up = "low";
// synopsys translate_on

// Location: FF_X68_Y38_N11
dffeas \register[18][13] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\register~82_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~33_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\register[18][13]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \register[18][13] .is_wysiwyg = "true";
defparam \register[18][13] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X68_Y38_N10
cycloneive_lcell_comb \Mux50~2 (
// Equation(s):
// \Mux50~2_combout  = (Selector8 & ((\register[22][13]~q ) # ((Selector7)))) # (!Selector8 & (((\register[18][13]~q  & !Selector7))))

	.dataa(\register[22][13]~q ),
	.datab(Selector8),
	.datac(\register[18][13]~q ),
	.datad(Selector7),
	.cin(gnd),
	.combout(\Mux50~2_combout ),
	.cout());
// synopsys translate_off
defparam \Mux50~2 .lut_mask = 16'hCCB8;
defparam \Mux50~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X68_Y38_N8
cycloneive_lcell_comb \Mux50~3 (
// Equation(s):
// \Mux50~3_combout  = (Selector7 & ((\Mux50~2_combout  & ((\register[30][13]~q ))) # (!\Mux50~2_combout  & (\register[26][13]~q )))) # (!Selector7 & (((\Mux50~2_combout ))))

	.dataa(Selector7),
	.datab(\register[26][13]~q ),
	.datac(\register[30][13]~q ),
	.datad(\Mux50~2_combout ),
	.cin(gnd),
	.combout(\Mux50~3_combout ),
	.cout());
// synopsys translate_off
defparam \Mux50~3 .lut_mask = 16'hF588;
defparam \Mux50~3 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X65_Y38_N18
cycloneive_lcell_comb \Mux50~6 (
// Equation(s):
// \Mux50~6_combout  = (Selector10 & (((Selector91)))) # (!Selector10 & ((Selector91 & ((\Mux50~3_combout ))) # (!Selector91 & (\Mux50~5_combout ))))

	.dataa(Selector10),
	.datab(\Mux50~5_combout ),
	.datac(Selector91),
	.datad(\Mux50~3_combout ),
	.cin(gnd),
	.combout(\Mux50~6_combout ),
	.cout());
// synopsys translate_off
defparam \Mux50~6 .lut_mask = 16'hF4A4;
defparam \Mux50~6 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X60_Y36_N7
dffeas \register[12][13] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\register~82_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~52_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\register[12][13]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \register[12][13] .is_wysiwyg = "true";
defparam \register[12][13] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X60_Y36_N6
cycloneive_lcell_comb \Mux50~17 (
// Equation(s):
// \Mux50~17_combout  = (Selector10 & ((\register[13][13]~q ) # ((Selector91)))) # (!Selector10 & (((\register[12][13]~q  & !Selector91))))

	.dataa(\register[13][13]~q ),
	.datab(Selector10),
	.datac(\register[12][13]~q ),
	.datad(Selector91),
	.cin(gnd),
	.combout(\Mux50~17_combout ),
	.cout());
// synopsys translate_off
defparam \Mux50~17 .lut_mask = 16'hCCB8;
defparam \Mux50~17 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X61_Y36_N27
dffeas \register[15][13] (
	.clk(!CLK),
	.d(\register~82_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~53_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\register[15][13]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \register[15][13] .is_wysiwyg = "true";
defparam \register[15][13] .power_up = "low";
// synopsys translate_on

// Location: FF_X60_Y36_N17
dffeas \register[14][13] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\register~82_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~61_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\register[14][13]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \register[14][13] .is_wysiwyg = "true";
defparam \register[14][13] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X65_Y36_N20
cycloneive_lcell_comb \Mux50~18 (
// Equation(s):
// \Mux50~18_combout  = (\Mux50~17_combout  & ((\register[15][13]~q ) # ((!Selector91)))) # (!\Mux50~17_combout  & (((\register[14][13]~q  & Selector91))))

	.dataa(\Mux50~17_combout ),
	.datab(\register[15][13]~q ),
	.datac(\register[14][13]~q ),
	.datad(Selector91),
	.cin(gnd),
	.combout(\Mux50~18_combout ),
	.cout());
// synopsys translate_off
defparam \Mux50~18 .lut_mask = 16'hD8AA;
defparam \Mux50~18 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X68_Y32_N27
dffeas \register[7][13] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\register~82_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~43_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\register[7][13]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \register[7][13] .is_wysiwyg = "true";
defparam \register[7][13] .power_up = "low";
// synopsys translate_on

// Location: FF_X69_Y32_N17
dffeas \register[5][13] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\register~82_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~59_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\register[5][13]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \register[5][13] .is_wysiwyg = "true";
defparam \register[5][13] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X69_Y32_N16
cycloneive_lcell_comb \Mux50~10 (
// Equation(s):
// \Mux50~10_combout  = (Selector91 & (((Selector10)))) # (!Selector91 & ((Selector10 & ((\register[5][13]~q ))) # (!Selector10 & (\register[4][13]~q ))))

	.dataa(\register[4][13]~q ),
	.datab(Selector91),
	.datac(\register[5][13]~q ),
	.datad(Selector10),
	.cin(gnd),
	.combout(\Mux50~10_combout ),
	.cout());
// synopsys translate_off
defparam \Mux50~10 .lut_mask = 16'hFC22;
defparam \Mux50~10 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X68_Y32_N25
dffeas \register[6][13] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\register~82_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~58_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\register[6][13]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \register[6][13] .is_wysiwyg = "true";
defparam \register[6][13] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X68_Y32_N24
cycloneive_lcell_comb \Mux50~11 (
// Equation(s):
// \Mux50~11_combout  = (\Mux50~10_combout  & ((\register[7][13]~q ) # ((!Selector91)))) # (!\Mux50~10_combout  & (((\register[6][13]~q  & Selector91))))

	.dataa(\register[7][13]~q ),
	.datab(\Mux50~10_combout ),
	.datac(\register[6][13]~q ),
	.datad(Selector91),
	.cin(gnd),
	.combout(\Mux50~11_combout ),
	.cout());
// synopsys translate_off
defparam \Mux50~11 .lut_mask = 16'hB8CC;
defparam \Mux50~11 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X66_Y34_N17
dffeas \register[2][13] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\register~82_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~50_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\register[2][13]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \register[2][13] .is_wysiwyg = "true";
defparam \register[2][13] .power_up = "low";
// synopsys translate_on

// Location: FF_X65_Y36_N19
dffeas \register[1][13] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\register~82_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~49_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\register[1][13]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \register[1][13] .is_wysiwyg = "true";
defparam \register[1][13] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X65_Y36_N18
cycloneive_lcell_comb \Mux50~14 (
// Equation(s):
// \Mux50~14_combout  = (Selector10 & ((Selector91 & (\register[3][13]~q )) # (!Selector91 & ((\register[1][13]~q )))))

	.dataa(\register[3][13]~q ),
	.datab(Selector91),
	.datac(\register[1][13]~q ),
	.datad(Selector10),
	.cin(gnd),
	.combout(\Mux50~14_combout ),
	.cout());
// synopsys translate_off
defparam \Mux50~14 .lut_mask = 16'hB800;
defparam \Mux50~14 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X65_Y36_N4
cycloneive_lcell_comb \Mux50~15 (
// Equation(s):
// \Mux50~15_combout  = (\Mux50~14_combout ) # ((Selector91 & (\register[2][13]~q  & !Selector10)))

	.dataa(Selector91),
	.datab(\register[2][13]~q ),
	.datac(\Mux50~14_combout ),
	.datad(Selector10),
	.cin(gnd),
	.combout(\Mux50~15_combout ),
	.cout());
// synopsys translate_off
defparam \Mux50~15 .lut_mask = 16'hF0F8;
defparam \Mux50~15 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X63_Y40_N13
dffeas \register[9][13] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\register~82_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~44_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\register[9][13]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \register[9][13] .is_wysiwyg = "true";
defparam \register[9][13] .power_up = "low";
// synopsys translate_on

// Location: FF_X62_Y40_N25
dffeas \register[10][13] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\register~82_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~45_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\register[10][13]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \register[10][13] .is_wysiwyg = "true";
defparam \register[10][13] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X62_Y40_N24
cycloneive_lcell_comb \Mux50~12 (
// Equation(s):
// \Mux50~12_combout  = (Selector91 & (((\register[10][13]~q ) # (Selector10)))) # (!Selector91 & (\register[8][13]~q  & ((!Selector10))))

	.dataa(\register[8][13]~q ),
	.datab(Selector91),
	.datac(\register[10][13]~q ),
	.datad(Selector10),
	.cin(gnd),
	.combout(\Mux50~12_combout ),
	.cout());
// synopsys translate_off
defparam \Mux50~12 .lut_mask = 16'hCCE2;
defparam \Mux50~12 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X63_Y40_N12
cycloneive_lcell_comb \Mux50~13 (
// Equation(s):
// \Mux50~13_combout  = (Selector10 & ((\Mux50~12_combout  & (\register[11][13]~q )) # (!\Mux50~12_combout  & ((\register[9][13]~q ))))) # (!Selector10 & (((\Mux50~12_combout ))))

	.dataa(\register[11][13]~q ),
	.datab(Selector10),
	.datac(\register[9][13]~q ),
	.datad(\Mux50~12_combout ),
	.cin(gnd),
	.combout(\Mux50~13_combout ),
	.cout());
// synopsys translate_off
defparam \Mux50~13 .lut_mask = 16'hBBC0;
defparam \Mux50~13 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X65_Y36_N2
cycloneive_lcell_comb \Mux50~16 (
// Equation(s):
// \Mux50~16_combout  = (Selector7 & ((Selector8) # ((\Mux50~13_combout )))) # (!Selector7 & (!Selector8 & (\Mux50~15_combout )))

	.dataa(Selector7),
	.datab(Selector8),
	.datac(\Mux50~15_combout ),
	.datad(\Mux50~13_combout ),
	.cin(gnd),
	.combout(\Mux50~16_combout ),
	.cout());
// synopsys translate_off
defparam \Mux50~16 .lut_mask = 16'hBA98;
defparam \Mux50~16 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y35_N28
cycloneive_lcell_comb \register~83 (
// Equation(s):
// \register~83_combout  = (WideOr01 & ((\wdat[12]~38_combout ) # ((plif_memwbregsrc_l_1 & plif_memwbrtnaddr_l_12))))

	.dataa(WideOr0),
	.datab(plif_memwbregsrc_l_1),
	.datac(plif_memwbrtnaddr_l_12),
	.datad(wdat_12),
	.cin(gnd),
	.combout(\register~83_combout ),
	.cout());
// synopsys translate_off
defparam \register~83 .lut_mask = 16'hAA80;
defparam \register~83 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y30_N20
cycloneive_lcell_comb \register[31][12]~feeder (
// Equation(s):
// \register[31][12]~feeder_combout  = \register~83_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(\register~83_combout ),
	.cin(gnd),
	.combout(\register[31][12]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \register[31][12]~feeder .lut_mask = 16'hFF00;
defparam \register[31][12]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X61_Y30_N21
dffeas \register[31][12] (
	.clk(!CLK),
	.d(\register[31][12]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~40_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\register[31][12]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \register[31][12] .is_wysiwyg = "true";
defparam \register[31][12] .power_up = "low";
// synopsys translate_on

// Location: FF_X60_Y37_N15
dffeas \register[19][12] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\register~83_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~39_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\register[19][12]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \register[19][12] .is_wysiwyg = "true";
defparam \register[19][12] .power_up = "low";
// synopsys translate_on

// Location: FF_X62_Y38_N19
dffeas \register[23][12] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\register~83_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~37_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\register[23][12]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \register[23][12] .is_wysiwyg = "true";
defparam \register[23][12] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X62_Y38_N18
cycloneive_lcell_comb \Mux51~7 (
// Equation(s):
// \Mux51~7_combout  = (Selector8 & (((\register[23][12]~q ) # (Selector7)))) # (!Selector8 & (\register[19][12]~q  & ((!Selector7))))

	.dataa(Selector8),
	.datab(\register[19][12]~q ),
	.datac(\register[23][12]~q ),
	.datad(Selector7),
	.cin(gnd),
	.combout(\Mux51~7_combout ),
	.cout());
// synopsys translate_off
defparam \Mux51~7 .lut_mask = 16'hAAE4;
defparam \Mux51~7 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y39_N2
cycloneive_lcell_comb \register[27][12]~feeder (
// Equation(s):
// \register[27][12]~feeder_combout  = \register~83_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(\register~83_combout ),
	.datad(gnd),
	.cin(gnd),
	.combout(\register[27][12]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \register[27][12]~feeder .lut_mask = 16'hF0F0;
defparam \register[27][12]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X62_Y39_N3
dffeas \register[27][12] (
	.clk(!CLK),
	.d(\register[27][12]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~38_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\register[27][12]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \register[27][12] .is_wysiwyg = "true";
defparam \register[27][12] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X61_Y30_N22
cycloneive_lcell_comb \Mux51~8 (
// Equation(s):
// \Mux51~8_combout  = (Selector7 & ((\Mux51~7_combout  & (\register[31][12]~q )) # (!\Mux51~7_combout  & ((\register[27][12]~q ))))) # (!Selector7 & (((\Mux51~7_combout ))))

	.dataa(Selector7),
	.datab(\register[31][12]~q ),
	.datac(\Mux51~7_combout ),
	.datad(\register[27][12]~q ),
	.cin(gnd),
	.combout(\Mux51~8_combout ),
	.cout());
// synopsys translate_off
defparam \Mux51~8 .lut_mask = 16'hDAD0;
defparam \Mux51~8 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X60_Y37_N13
dffeas \register[17][12] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\register~83_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~26_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\register[17][12]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \register[17][12] .is_wysiwyg = "true";
defparam \register[17][12] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X63_Y33_N10
cycloneive_lcell_comb \register[21][12]~feeder (
// Equation(s):
// \register[21][12]~feeder_combout  = \register~83_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(\register~83_combout ),
	.cin(gnd),
	.combout(\register[21][12]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \register[21][12]~feeder .lut_mask = 16'hFF00;
defparam \register[21][12]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X63_Y33_N11
dffeas \register[21][12] (
	.clk(!CLK),
	.d(\register[21][12]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~22_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\register[21][12]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \register[21][12] .is_wysiwyg = "true";
defparam \register[21][12] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X60_Y37_N12
cycloneive_lcell_comb \Mux51~0 (
// Equation(s):
// \Mux51~0_combout  = (Selector8 & ((Selector7) # ((\register[21][12]~q )))) # (!Selector8 & (!Selector7 & (\register[17][12]~q )))

	.dataa(Selector8),
	.datab(Selector7),
	.datac(\register[17][12]~q ),
	.datad(\register[21][12]~q ),
	.cin(gnd),
	.combout(\Mux51~0_combout ),
	.cout());
// synopsys translate_off
defparam \Mux51~0 .lut_mask = 16'hBA98;
defparam \Mux51~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X60_Y34_N31
dffeas \register[25][12] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\register~83_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~24_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\register[25][12]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \register[25][12] .is_wysiwyg = "true";
defparam \register[25][12] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X63_Y33_N28
cycloneive_lcell_comb \register[29][12]~feeder (
// Equation(s):
// \register[29][12]~feeder_combout  = \register~83_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(\register~83_combout ),
	.cin(gnd),
	.combout(\register[29][12]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \register[29][12]~feeder .lut_mask = 16'hFF00;
defparam \register[29][12]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X63_Y33_N29
dffeas \register[29][12] (
	.clk(!CLK),
	.d(\register[29][12]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~28_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\register[29][12]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \register[29][12] .is_wysiwyg = "true";
defparam \register[29][12] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X63_Y33_N18
cycloneive_lcell_comb \Mux51~1 (
// Equation(s):
// \Mux51~1_combout  = (\Mux51~0_combout  & (((\register[29][12]~q )) # (!Selector7))) # (!\Mux51~0_combout  & (Selector7 & (\register[25][12]~q )))

	.dataa(\Mux51~0_combout ),
	.datab(Selector7),
	.datac(\register[25][12]~q ),
	.datad(\register[29][12]~q ),
	.cin(gnd),
	.combout(\Mux51~1_combout ),
	.cout());
// synopsys translate_off
defparam \Mux51~1 .lut_mask = 16'hEA62;
defparam \Mux51~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X69_Y36_N8
cycloneive_lcell_comb \register[30][12]~feeder (
// Equation(s):
// \register[30][12]~feeder_combout  = \register~83_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(\register~83_combout ),
	.cin(gnd),
	.combout(\register[30][12]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \register[30][12]~feeder .lut_mask = 16'hFF00;
defparam \register[30][12]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X69_Y36_N9
dffeas \register[30][12] (
	.clk(!CLK),
	.d(\register[30][12]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~56_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\register[30][12]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \register[30][12] .is_wysiwyg = "true";
defparam \register[30][12] .power_up = "low";
// synopsys translate_on

// Location: FF_X68_Y38_N27
dffeas \register[26][12] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\register~83_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~54_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\register[26][12]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \register[26][12] .is_wysiwyg = "true";
defparam \register[26][12] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X69_Y37_N0
cycloneive_lcell_comb \register[18][12]~feeder (
// Equation(s):
// \register[18][12]~feeder_combout  = \register~83_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(\register~83_combout ),
	.datad(gnd),
	.cin(gnd),
	.combout(\register[18][12]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \register[18][12]~feeder .lut_mask = 16'hF0F0;
defparam \register[18][12]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X69_Y37_N1
dffeas \register[18][12] (
	.clk(!CLK),
	.d(\register[18][12]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~33_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\register[18][12]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \register[18][12] .is_wysiwyg = "true";
defparam \register[18][12] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X68_Y38_N26
cycloneive_lcell_comb \Mux51~2 (
// Equation(s):
// \Mux51~2_combout  = (Selector7 & ((Selector8) # ((\register[26][12]~q )))) # (!Selector7 & (!Selector8 & ((\register[18][12]~q ))))

	.dataa(Selector7),
	.datab(Selector8),
	.datac(\register[26][12]~q ),
	.datad(\register[18][12]~q ),
	.cin(gnd),
	.combout(\Mux51~2_combout ),
	.cout());
// synopsys translate_off
defparam \Mux51~2 .lut_mask = 16'hB9A8;
defparam \Mux51~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X69_Y36_N2
cycloneive_lcell_comb \Mux51~3 (
// Equation(s):
// \Mux51~3_combout  = (Selector8 & ((\Mux51~2_combout  & ((\register[30][12]~q ))) # (!\Mux51~2_combout  & (\register[22][12]~q )))) # (!Selector8 & (((\Mux51~2_combout ))))

	.dataa(\register[22][12]~q ),
	.datab(\register[30][12]~q ),
	.datac(Selector8),
	.datad(\Mux51~2_combout ),
	.cin(gnd),
	.combout(\Mux51~3_combout ),
	.cout());
// synopsys translate_off
defparam \Mux51~3 .lut_mask = 16'hCFA0;
defparam \Mux51~3 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X69_Y36_N24
cycloneive_lcell_comb \register[28][12]~feeder (
// Equation(s):
// \register[28][12]~feeder_combout  = \register~83_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(\register~83_combout ),
	.cin(gnd),
	.combout(\register[28][12]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \register[28][12]~feeder .lut_mask = 16'hFF00;
defparam \register[28][12]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X69_Y36_N25
dffeas \register[28][12] (
	.clk(!CLK),
	.d(\register[28][12]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~57_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\register[28][12]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \register[28][12] .is_wysiwyg = "true";
defparam \register[28][12] .power_up = "low";
// synopsys translate_on

// Location: FF_X69_Y38_N23
dffeas \register[20][12] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\register~83_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~35_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\register[20][12]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \register[20][12] .is_wysiwyg = "true";
defparam \register[20][12] .power_up = "low";
// synopsys translate_on

// Location: FF_X69_Y38_N25
dffeas \register[16][12] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\register~83_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~36_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\register[16][12]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \register[16][12] .is_wysiwyg = "true";
defparam \register[16][12] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X69_Y34_N12
cycloneive_lcell_comb \register[24][12]~feeder (
// Equation(s):
// \register[24][12]~feeder_combout  = \register~83_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(\register~83_combout ),
	.cin(gnd),
	.combout(\register[24][12]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \register[24][12]~feeder .lut_mask = 16'hFF00;
defparam \register[24][12]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X69_Y34_N13
dffeas \register[24][12] (
	.clk(!CLK),
	.d(\register[24][12]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~34_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\register[24][12]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \register[24][12] .is_wysiwyg = "true";
defparam \register[24][12] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X69_Y34_N6
cycloneive_lcell_comb \Mux51~4 (
// Equation(s):
// \Mux51~4_combout  = (Selector7 & ((Selector8) # ((\register[24][12]~q )))) # (!Selector7 & (!Selector8 & (\register[16][12]~q )))

	.dataa(Selector7),
	.datab(Selector8),
	.datac(\register[16][12]~q ),
	.datad(\register[24][12]~q ),
	.cin(gnd),
	.combout(\Mux51~4_combout ),
	.cout());
// synopsys translate_off
defparam \Mux51~4 .lut_mask = 16'hBA98;
defparam \Mux51~4 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X69_Y38_N22
cycloneive_lcell_comb \Mux51~5 (
// Equation(s):
// \Mux51~5_combout  = (Selector8 & ((\Mux51~4_combout  & (\register[28][12]~q )) # (!\Mux51~4_combout  & ((\register[20][12]~q ))))) # (!Selector8 & (((\Mux51~4_combout ))))

	.dataa(Selector8),
	.datab(\register[28][12]~q ),
	.datac(\register[20][12]~q ),
	.datad(\Mux51~4_combout ),
	.cin(gnd),
	.combout(\Mux51~5_combout ),
	.cout());
// synopsys translate_off
defparam \Mux51~5 .lut_mask = 16'hDDA0;
defparam \Mux51~5 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y30_N6
cycloneive_lcell_comb \Mux51~6 (
// Equation(s):
// \Mux51~6_combout  = (Selector10 & (Selector91)) # (!Selector10 & ((Selector91 & (\Mux51~3_combout )) # (!Selector91 & ((\Mux51~5_combout )))))

	.dataa(Selector10),
	.datab(Selector91),
	.datac(\Mux51~3_combout ),
	.datad(\Mux51~5_combout ),
	.cin(gnd),
	.combout(\Mux51~6_combout ),
	.cout());
// synopsys translate_off
defparam \Mux51~6 .lut_mask = 16'hD9C8;
defparam \Mux51~6 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X63_Y40_N17
dffeas \register[9][12] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\register~83_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~44_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\register[9][12]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \register[9][12] .is_wysiwyg = "true";
defparam \register[9][12] .power_up = "low";
// synopsys translate_on

// Location: FF_X63_Y40_N27
dffeas \register[11][12] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\register~83_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~47_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\register[11][12]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \register[11][12] .is_wysiwyg = "true";
defparam \register[11][12] .power_up = "low";
// synopsys translate_on

// Location: FF_X62_Y40_N29
dffeas \register[10][12] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\register~83_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~45_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\register[10][12]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \register[10][12] .is_wysiwyg = "true";
defparam \register[10][12] .power_up = "low";
// synopsys translate_on

// Location: FF_X62_Y40_N19
dffeas \register[8][12] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\register~83_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~46_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\register[8][12]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \register[8][12] .is_wysiwyg = "true";
defparam \register[8][12] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X62_Y40_N18
cycloneive_lcell_comb \Mux51~10 (
// Equation(s):
// \Mux51~10_combout  = (Selector91 & ((\register[10][12]~q ) # ((Selector10)))) # (!Selector91 & (((\register[8][12]~q  & !Selector10))))

	.dataa(Selector91),
	.datab(\register[10][12]~q ),
	.datac(\register[8][12]~q ),
	.datad(Selector10),
	.cin(gnd),
	.combout(\Mux51~10_combout ),
	.cout());
// synopsys translate_off
defparam \Mux51~10 .lut_mask = 16'hAAD8;
defparam \Mux51~10 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X63_Y40_N26
cycloneive_lcell_comb \Mux51~11 (
// Equation(s):
// \Mux51~11_combout  = (Selector10 & ((\Mux51~10_combout  & ((\register[11][12]~q ))) # (!\Mux51~10_combout  & (\register[9][12]~q )))) # (!Selector10 & (((\Mux51~10_combout ))))

	.dataa(Selector10),
	.datab(\register[9][12]~q ),
	.datac(\register[11][12]~q ),
	.datad(\Mux51~10_combout ),
	.cin(gnd),
	.combout(\Mux51~11_combout ),
	.cout());
// synopsys translate_off
defparam \Mux51~11 .lut_mask = 16'hF588;
defparam \Mux51~11 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X60_Y34_N21
dffeas \register[14][12] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\register~83_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~61_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\register[14][12]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \register[14][12] .is_wysiwyg = "true";
defparam \register[14][12] .power_up = "low";
// synopsys translate_on

// Location: FF_X61_Y35_N29
dffeas \register[15][12] (
	.clk(!CLK),
	.d(\register~83_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~53_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\register[15][12]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \register[15][12] .is_wysiwyg = "true";
defparam \register[15][12] .power_up = "low";
// synopsys translate_on

// Location: FF_X60_Y33_N7
dffeas \register[12][12] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\register~83_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~52_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\register[12][12]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \register[12][12] .is_wysiwyg = "true";
defparam \register[12][12] .power_up = "low";
// synopsys translate_on

// Location: FF_X60_Y33_N1
dffeas \register[13][12] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\register~83_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~62_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\register[13][12]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \register[13][12] .is_wysiwyg = "true";
defparam \register[13][12] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X60_Y33_N6
cycloneive_lcell_comb \Mux51~17 (
// Equation(s):
// \Mux51~17_combout  = (Selector10 & ((Selector91) # ((\register[13][12]~q )))) # (!Selector10 & (!Selector91 & (\register[12][12]~q )))

	.dataa(Selector10),
	.datab(Selector91),
	.datac(\register[12][12]~q ),
	.datad(\register[13][12]~q ),
	.cin(gnd),
	.combout(\Mux51~17_combout ),
	.cout());
// synopsys translate_off
defparam \Mux51~17 .lut_mask = 16'hBA98;
defparam \Mux51~17 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y30_N8
cycloneive_lcell_comb \Mux51~18 (
// Equation(s):
// \Mux51~18_combout  = (Selector91 & ((\Mux51~17_combout  & ((\register[15][12]~q ))) # (!\Mux51~17_combout  & (\register[14][12]~q )))) # (!Selector91 & (((\Mux51~17_combout ))))

	.dataa(\register[14][12]~q ),
	.datab(Selector91),
	.datac(\register[15][12]~q ),
	.datad(\Mux51~17_combout ),
	.cin(gnd),
	.combout(\Mux51~18_combout ),
	.cout());
// synopsys translate_off
defparam \Mux51~18 .lut_mask = 16'hF388;
defparam \Mux51~18 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X67_Y33_N22
cycloneive_lcell_comb \register[6][12]~feeder (
// Equation(s):
// \register[6][12]~feeder_combout  = \register~83_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(\register~83_combout ),
	.datad(gnd),
	.cin(gnd),
	.combout(\register[6][12]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \register[6][12]~feeder .lut_mask = 16'hF0F0;
defparam \register[6][12]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X67_Y33_N23
dffeas \register[6][12] (
	.clk(!CLK),
	.d(\register[6][12]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~58_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\register[6][12]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \register[6][12] .is_wysiwyg = "true";
defparam \register[6][12] .power_up = "low";
// synopsys translate_on

// Location: FF_X68_Y33_N25
dffeas \register[7][12] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\register~83_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~43_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\register[7][12]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \register[7][12] .is_wysiwyg = "true";
defparam \register[7][12] .power_up = "low";
// synopsys translate_on

// Location: FF_X69_Y32_N13
dffeas \register[5][12] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\register~83_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~59_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\register[5][12]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \register[5][12] .is_wysiwyg = "true";
defparam \register[5][12] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X69_Y32_N12
cycloneive_lcell_comb \Mux51~12 (
// Equation(s):
// \Mux51~12_combout  = (Selector91 & (((Selector10)))) # (!Selector91 & ((Selector10 & ((\register[5][12]~q ))) # (!Selector10 & (\register[4][12]~q ))))

	.dataa(\register[4][12]~q ),
	.datab(Selector91),
	.datac(\register[5][12]~q ),
	.datad(Selector10),
	.cin(gnd),
	.combout(\Mux51~12_combout ),
	.cout());
// synopsys translate_off
defparam \Mux51~12 .lut_mask = 16'hFC22;
defparam \Mux51~12 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X68_Y33_N24
cycloneive_lcell_comb \Mux51~13 (
// Equation(s):
// \Mux51~13_combout  = (Selector91 & ((\Mux51~12_combout  & ((\register[7][12]~q ))) # (!\Mux51~12_combout  & (\register[6][12]~q )))) # (!Selector91 & (((\Mux51~12_combout ))))

	.dataa(Selector91),
	.datab(\register[6][12]~q ),
	.datac(\register[7][12]~q ),
	.datad(\Mux51~12_combout ),
	.cin(gnd),
	.combout(\Mux51~13_combout ),
	.cout());
// synopsys translate_off
defparam \Mux51~13 .lut_mask = 16'hF588;
defparam \Mux51~13 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X68_Y33_N23
dffeas \register[2][12] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\register~83_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~50_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\register[2][12]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \register[2][12] .is_wysiwyg = "true";
defparam \register[2][12] .power_up = "low";
// synopsys translate_on

// Location: FF_X65_Y33_N29
dffeas \register[3][12] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\register~83_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~48_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\register[3][12]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \register[3][12] .is_wysiwyg = "true";
defparam \register[3][12] .power_up = "low";
// synopsys translate_on

// Location: FF_X65_Y33_N31
dffeas \register[1][12] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\register~83_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~49_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\register[1][12]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \register[1][12] .is_wysiwyg = "true";
defparam \register[1][12] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X65_Y33_N30
cycloneive_lcell_comb \Mux51~14 (
// Equation(s):
// \Mux51~14_combout  = (Selector10 & ((Selector91 & (\register[3][12]~q )) # (!Selector91 & ((\register[1][12]~q )))))

	.dataa(Selector91),
	.datab(\register[3][12]~q ),
	.datac(\register[1][12]~q ),
	.datad(Selector10),
	.cin(gnd),
	.combout(\Mux51~14_combout ),
	.cout());
// synopsys translate_off
defparam \Mux51~14 .lut_mask = 16'hD800;
defparam \Mux51~14 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X68_Y33_N22
cycloneive_lcell_comb \Mux51~15 (
// Equation(s):
// \Mux51~15_combout  = (\Mux51~14_combout ) # ((!Selector10 & (Selector91 & \register[2][12]~q )))

	.dataa(Selector10),
	.datab(Selector91),
	.datac(\register[2][12]~q ),
	.datad(\Mux51~14_combout ),
	.cin(gnd),
	.combout(\Mux51~15_combout ),
	.cout());
// synopsys translate_off
defparam \Mux51~15 .lut_mask = 16'hFF40;
defparam \Mux51~15 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y30_N10
cycloneive_lcell_comb \Mux51~16 (
// Equation(s):
// \Mux51~16_combout  = (Selector7 & (Selector8)) # (!Selector7 & ((Selector8 & (\Mux51~13_combout )) # (!Selector8 & ((\Mux51~15_combout )))))

	.dataa(Selector7),
	.datab(Selector8),
	.datac(\Mux51~13_combout ),
	.datad(\Mux51~15_combout ),
	.cin(gnd),
	.combout(\Mux51~16_combout ),
	.cout());
// synopsys translate_off
defparam \Mux51~16 .lut_mask = 16'hD9C8;
defparam \Mux51~16 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y35_N14
cycloneive_lcell_comb \register~84 (
// Equation(s):
// \register~84_combout  = (WideOr01 & ((\wdat[11]~40_combout ) # ((plif_memwbregsrc_l_1 & plif_memwbrtnaddr_l_11))))

	.dataa(WideOr0),
	.datab(plif_memwbregsrc_l_1),
	.datac(plif_memwbrtnaddr_l_11),
	.datad(wdat_11),
	.cin(gnd),
	.combout(\register~84_combout ),
	.cout());
// synopsys translate_off
defparam \register~84 .lut_mask = 16'hAA80;
defparam \register~84 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y33_N10
cycloneive_lcell_comb \register[21][11]~feeder (
// Equation(s):
// \register[21][11]~feeder_combout  = \register~84_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(\register~84_combout ),
	.cin(gnd),
	.combout(\register[21][11]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \register[21][11]~feeder .lut_mask = 16'hFF00;
defparam \register[21][11]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X62_Y33_N11
dffeas \register[21][11] (
	.clk(!CLK),
	.d(\register[21][11]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~22_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\register[21][11]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \register[21][11] .is_wysiwyg = "true";
defparam \register[21][11] .power_up = "low";
// synopsys translate_on

// Location: FF_X62_Y34_N11
dffeas \register[17][11] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\register~84_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~26_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\register[17][11]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \register[17][11] .is_wysiwyg = "true";
defparam \register[17][11] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X63_Y38_N26
cycloneive_lcell_comb \register[25][11]~feeder (
// Equation(s):
// \register[25][11]~feeder_combout  = \register~84_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(\register~84_combout ),
	.cin(gnd),
	.combout(\register[25][11]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \register[25][11]~feeder .lut_mask = 16'hFF00;
defparam \register[25][11]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X63_Y38_N27
dffeas \register[25][11] (
	.clk(!CLK),
	.d(\register[25][11]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~24_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\register[25][11]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \register[25][11] .is_wysiwyg = "true";
defparam \register[25][11] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X62_Y34_N10
cycloneive_lcell_comb \Mux52~0 (
// Equation(s):
// \Mux52~0_combout  = (Selector7 & ((Selector8) # ((\register[25][11]~q )))) # (!Selector7 & (!Selector8 & (\register[17][11]~q )))

	.dataa(Selector7),
	.datab(Selector8),
	.datac(\register[17][11]~q ),
	.datad(\register[25][11]~q ),
	.cin(gnd),
	.combout(\Mux52~0_combout ),
	.cout());
// synopsys translate_off
defparam \Mux52~0 .lut_mask = 16'hBA98;
defparam \Mux52~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X61_Y38_N5
dffeas \register[29][11] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\register~84_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~28_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\register[29][11]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \register[29][11] .is_wysiwyg = "true";
defparam \register[29][11] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X61_Y38_N4
cycloneive_lcell_comb \Mux52~1 (
// Equation(s):
// \Mux52~1_combout  = (\Mux52~0_combout  & (((\register[29][11]~q ) # (!Selector8)))) # (!\Mux52~0_combout  & (\register[21][11]~q  & ((Selector8))))

	.dataa(\register[21][11]~q ),
	.datab(\Mux52~0_combout ),
	.datac(\register[29][11]~q ),
	.datad(Selector8),
	.cin(gnd),
	.combout(\Mux52~1_combout ),
	.cout());
// synopsys translate_off
defparam \Mux52~1 .lut_mask = 16'hE2CC;
defparam \Mux52~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X60_Y40_N21
dffeas \register[23][11] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\register~84_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~37_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\register[23][11]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \register[23][11] .is_wysiwyg = "true";
defparam \register[23][11] .power_up = "low";
// synopsys translate_on

// Location: FF_X61_Y38_N19
dffeas \register[31][11] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\register~84_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~40_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\register[31][11]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \register[31][11] .is_wysiwyg = "true";
defparam \register[31][11] .power_up = "low";
// synopsys translate_on

// Location: FF_X60_Y38_N13
dffeas \register[19][11] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\register~84_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~39_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\register[19][11]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \register[19][11] .is_wysiwyg = "true";
defparam \register[19][11] .power_up = "low";
// synopsys translate_on

// Location: FF_X60_Y38_N7
dffeas \register[27][11] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\register~84_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~38_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\register[27][11]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \register[27][11] .is_wysiwyg = "true";
defparam \register[27][11] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X60_Y38_N12
cycloneive_lcell_comb \Mux52~7 (
// Equation(s):
// \Mux52~7_combout  = (Selector8 & (Selector7)) # (!Selector8 & ((Selector7 & ((\register[27][11]~q ))) # (!Selector7 & (\register[19][11]~q ))))

	.dataa(Selector8),
	.datab(Selector7),
	.datac(\register[19][11]~q ),
	.datad(\register[27][11]~q ),
	.cin(gnd),
	.combout(\Mux52~7_combout ),
	.cout());
// synopsys translate_off
defparam \Mux52~7 .lut_mask = 16'hDC98;
defparam \Mux52~7 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y38_N18
cycloneive_lcell_comb \Mux52~8 (
// Equation(s):
// \Mux52~8_combout  = (Selector8 & ((\Mux52~7_combout  & ((\register[31][11]~q ))) # (!\Mux52~7_combout  & (\register[23][11]~q )))) # (!Selector8 & (((\Mux52~7_combout ))))

	.dataa(\register[23][11]~q ),
	.datab(Selector8),
	.datac(\register[31][11]~q ),
	.datad(\Mux52~7_combout ),
	.cin(gnd),
	.combout(\Mux52~8_combout ),
	.cout());
// synopsys translate_off
defparam \Mux52~8 .lut_mask = 16'hF388;
defparam \Mux52~8 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X68_Y38_N5
dffeas \register[26][11] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\register~84_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~54_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\register[26][11]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \register[26][11] .is_wysiwyg = "true";
defparam \register[26][11] .power_up = "low";
// synopsys translate_on

// Location: FF_X68_Y39_N5
dffeas \register[30][11] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\register~84_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~56_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\register[30][11]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \register[30][11] .is_wysiwyg = "true";
defparam \register[30][11] .power_up = "low";
// synopsys translate_on

// Location: FF_X68_Y38_N7
dffeas \register[18][11] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\register~84_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~33_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\register[18][11]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \register[18][11] .is_wysiwyg = "true";
defparam \register[18][11] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X68_Y38_N6
cycloneive_lcell_comb \Mux52~2 (
// Equation(s):
// \Mux52~2_combout  = (Selector8 & ((\register[22][11]~q ) # ((Selector7)))) # (!Selector8 & (((\register[18][11]~q  & !Selector7))))

	.dataa(\register[22][11]~q ),
	.datab(Selector8),
	.datac(\register[18][11]~q ),
	.datad(Selector7),
	.cin(gnd),
	.combout(\Mux52~2_combout ),
	.cout());
// synopsys translate_off
defparam \Mux52~2 .lut_mask = 16'hCCB8;
defparam \Mux52~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X68_Y38_N12
cycloneive_lcell_comb \Mux52~3 (
// Equation(s):
// \Mux52~3_combout  = (Selector7 & ((\Mux52~2_combout  & ((\register[30][11]~q ))) # (!\Mux52~2_combout  & (\register[26][11]~q )))) # (!Selector7 & (((\Mux52~2_combout ))))

	.dataa(Selector7),
	.datab(\register[26][11]~q ),
	.datac(\register[30][11]~q ),
	.datad(\Mux52~2_combout ),
	.cin(gnd),
	.combout(\Mux52~3_combout ),
	.cout());
// synopsys translate_off
defparam \Mux52~3 .lut_mask = 16'hF588;
defparam \Mux52~3 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y40_N22
cycloneive_lcell_comb \register[28][11]~feeder (
// Equation(s):
// \register[28][11]~feeder_combout  = \register~84_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(\register~84_combout ),
	.datad(gnd),
	.cin(gnd),
	.combout(\register[28][11]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \register[28][11]~feeder .lut_mask = 16'hF0F0;
defparam \register[28][11]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X61_Y40_N23
dffeas \register[28][11] (
	.clk(!CLK),
	.d(\register[28][11]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~57_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\register[28][11]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \register[28][11] .is_wysiwyg = "true";
defparam \register[28][11] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X69_Y38_N8
cycloneive_lcell_comb \register[16][11]~feeder (
// Equation(s):
// \register[16][11]~feeder_combout  = \register~84_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(\register~84_combout ),
	.datad(gnd),
	.cin(gnd),
	.combout(\register[16][11]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \register[16][11]~feeder .lut_mask = 16'hF0F0;
defparam \register[16][11]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X69_Y38_N9
dffeas \register[16][11] (
	.clk(!CLK),
	.d(\register[16][11]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~36_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\register[16][11]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \register[16][11] .is_wysiwyg = "true";
defparam \register[16][11] .power_up = "low";
// synopsys translate_on

// Location: FF_X69_Y38_N3
dffeas \register[20][11] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\register~84_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~35_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\register[20][11]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \register[20][11] .is_wysiwyg = "true";
defparam \register[20][11] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X69_Y38_N2
cycloneive_lcell_comb \Mux52~4 (
// Equation(s):
// \Mux52~4_combout  = (Selector8 & (((\register[20][11]~q ) # (Selector7)))) # (!Selector8 & (\register[16][11]~q  & ((!Selector7))))

	.dataa(Selector8),
	.datab(\register[16][11]~q ),
	.datac(\register[20][11]~q ),
	.datad(Selector7),
	.cin(gnd),
	.combout(\Mux52~4_combout ),
	.cout());
// synopsys translate_off
defparam \Mux52~4 .lut_mask = 16'hAAE4;
defparam \Mux52~4 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y40_N28
cycloneive_lcell_comb \Mux52~5 (
// Equation(s):
// \Mux52~5_combout  = (Selector7 & ((\Mux52~4_combout  & ((\register[28][11]~q ))) # (!\Mux52~4_combout  & (\register[24][11]~q )))) # (!Selector7 & (((\Mux52~4_combout ))))

	.dataa(\register[24][11]~q ),
	.datab(Selector7),
	.datac(\register[28][11]~q ),
	.datad(\Mux52~4_combout ),
	.cin(gnd),
	.combout(\Mux52~5_combout ),
	.cout());
// synopsys translate_off
defparam \Mux52~5 .lut_mask = 16'hF388;
defparam \Mux52~5 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y40_N18
cycloneive_lcell_comb \Mux52~6 (
// Equation(s):
// \Mux52~6_combout  = (Selector10 & (Selector91)) # (!Selector10 & ((Selector91 & (\Mux52~3_combout )) # (!Selector91 & ((\Mux52~5_combout )))))

	.dataa(Selector10),
	.datab(Selector91),
	.datac(\Mux52~3_combout ),
	.datad(\Mux52~5_combout ),
	.cin(gnd),
	.combout(\Mux52~6_combout ),
	.cout());
// synopsys translate_off
defparam \Mux52~6 .lut_mask = 16'hD9C8;
defparam \Mux52~6 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X68_Y32_N23
dffeas \register[7][11] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\register~84_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~43_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\register[7][11]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \register[7][11] .is_wysiwyg = "true";
defparam \register[7][11] .power_up = "low";
// synopsys translate_on

// Location: FF_X69_Y32_N19
dffeas \register[4][11] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\register~84_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~60_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\register[4][11]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \register[4][11] .is_wysiwyg = "true";
defparam \register[4][11] .power_up = "low";
// synopsys translate_on

// Location: FF_X69_Y32_N9
dffeas \register[5][11] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\register~84_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~59_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\register[5][11]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \register[5][11] .is_wysiwyg = "true";
defparam \register[5][11] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X69_Y32_N8
cycloneive_lcell_comb \Mux52~10 (
// Equation(s):
// \Mux52~10_combout  = (Selector10 & (((\register[5][11]~q ) # (Selector91)))) # (!Selector10 & (\register[4][11]~q  & ((!Selector91))))

	.dataa(Selector10),
	.datab(\register[4][11]~q ),
	.datac(\register[5][11]~q ),
	.datad(Selector91),
	.cin(gnd),
	.combout(\Mux52~10_combout ),
	.cout());
// synopsys translate_off
defparam \Mux52~10 .lut_mask = 16'hAAE4;
defparam \Mux52~10 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X68_Y32_N1
dffeas \register[6][11] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\register~84_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~58_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\register[6][11]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \register[6][11] .is_wysiwyg = "true";
defparam \register[6][11] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X68_Y32_N0
cycloneive_lcell_comb \Mux52~11 (
// Equation(s):
// \Mux52~11_combout  = (\Mux52~10_combout  & ((\register[7][11]~q ) # ((!Selector91)))) # (!\Mux52~10_combout  & (((\register[6][11]~q  & Selector91))))

	.dataa(\register[7][11]~q ),
	.datab(\Mux52~10_combout ),
	.datac(\register[6][11]~q ),
	.datad(Selector91),
	.cin(gnd),
	.combout(\Mux52~11_combout ),
	.cout());
// synopsys translate_off
defparam \Mux52~11 .lut_mask = 16'hB8CC;
defparam \Mux52~11 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y33_N24
cycloneive_lcell_comb \register[14][11]~feeder (
// Equation(s):
// \register[14][11]~feeder_combout  = \register~84_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(\register~84_combout ),
	.cin(gnd),
	.combout(\register[14][11]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \register[14][11]~feeder .lut_mask = 16'hFF00;
defparam \register[14][11]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X62_Y33_N25
dffeas \register[14][11] (
	.clk(!CLK),
	.d(\register[14][11]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~61_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\register[14][11]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \register[14][11] .is_wysiwyg = "true";
defparam \register[14][11] .power_up = "low";
// synopsys translate_on

// Location: FF_X63_Y30_N13
dffeas \register[13][11] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\register~84_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~62_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\register[13][11]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \register[13][11] .is_wysiwyg = "true";
defparam \register[13][11] .power_up = "low";
// synopsys translate_on

// Location: FF_X63_Y30_N11
dffeas \register[12][11] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\register~84_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~52_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\register[12][11]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \register[12][11] .is_wysiwyg = "true";
defparam \register[12][11] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X63_Y30_N12
cycloneive_lcell_comb \Mux52~17 (
// Equation(s):
// \Mux52~17_combout  = (Selector91 & (Selector10)) # (!Selector91 & ((Selector10 & (\register[13][11]~q )) # (!Selector10 & ((\register[12][11]~q )))))

	.dataa(Selector91),
	.datab(Selector10),
	.datac(\register[13][11]~q ),
	.datad(\register[12][11]~q ),
	.cin(gnd),
	.combout(\Mux52~17_combout ),
	.cout());
// synopsys translate_off
defparam \Mux52~17 .lut_mask = 16'hD9C8;
defparam \Mux52~17 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X61_Y35_N15
dffeas \register[15][11] (
	.clk(!CLK),
	.d(\register~84_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~53_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\register[15][11]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \register[15][11] .is_wysiwyg = "true";
defparam \register[15][11] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X66_Y33_N4
cycloneive_lcell_comb \Mux52~18 (
// Equation(s):
// \Mux52~18_combout  = (Selector91 & ((\Mux52~17_combout  & ((\register[15][11]~q ))) # (!\Mux52~17_combout  & (\register[14][11]~q )))) # (!Selector91 & (((\Mux52~17_combout ))))

	.dataa(\register[14][11]~q ),
	.datab(Selector91),
	.datac(\Mux52~17_combout ),
	.datad(\register[15][11]~q ),
	.cin(gnd),
	.combout(\Mux52~18_combout ),
	.cout());
// synopsys translate_off
defparam \Mux52~18 .lut_mask = 16'hF838;
defparam \Mux52~18 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X66_Y34_N31
dffeas \register[2][11] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\register~84_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~50_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\register[2][11]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \register[2][11] .is_wysiwyg = "true";
defparam \register[2][11] .power_up = "low";
// synopsys translate_on

// Location: FF_X65_Y36_N15
dffeas \register[1][11] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\register~84_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~49_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\register[1][11]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \register[1][11] .is_wysiwyg = "true";
defparam \register[1][11] .power_up = "low";
// synopsys translate_on

// Location: FF_X65_Y36_N9
dffeas \register[3][11] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\register~84_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~48_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\register[3][11]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \register[3][11] .is_wysiwyg = "true";
defparam \register[3][11] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X65_Y36_N8
cycloneive_lcell_comb \Mux52~14 (
// Equation(s):
// \Mux52~14_combout  = (Selector10 & ((Selector91 & ((\register[3][11]~q ))) # (!Selector91 & (\register[1][11]~q ))))

	.dataa(Selector91),
	.datab(\register[1][11]~q ),
	.datac(\register[3][11]~q ),
	.datad(Selector10),
	.cin(gnd),
	.combout(\Mux52~14_combout ),
	.cout());
// synopsys translate_off
defparam \Mux52~14 .lut_mask = 16'hE400;
defparam \Mux52~14 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X66_Y33_N8
cycloneive_lcell_comb \Mux52~15 (
// Equation(s):
// \Mux52~15_combout  = (\Mux52~14_combout ) # ((!Selector10 & (Selector91 & \register[2][11]~q )))

	.dataa(Selector10),
	.datab(Selector91),
	.datac(\register[2][11]~q ),
	.datad(\Mux52~14_combout ),
	.cin(gnd),
	.combout(\Mux52~15_combout ),
	.cout());
// synopsys translate_off
defparam \Mux52~15 .lut_mask = 16'hFF40;
defparam \Mux52~15 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X63_Y40_N21
dffeas \register[9][11] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\register~84_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~44_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\register[9][11]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \register[9][11] .is_wysiwyg = "true";
defparam \register[9][11] .power_up = "low";
// synopsys translate_on

// Location: FF_X62_Y40_N13
dffeas \register[10][11] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\register~84_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~45_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\register[10][11]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \register[10][11] .is_wysiwyg = "true";
defparam \register[10][11] .power_up = "low";
// synopsys translate_on

// Location: FF_X62_Y40_N7
dffeas \register[8][11] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\register~84_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~46_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\register[8][11]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \register[8][11] .is_wysiwyg = "true";
defparam \register[8][11] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X62_Y40_N12
cycloneive_lcell_comb \Mux52~12 (
// Equation(s):
// \Mux52~12_combout  = (Selector10 & (Selector91)) # (!Selector10 & ((Selector91 & (\register[10][11]~q )) # (!Selector91 & ((\register[8][11]~q )))))

	.dataa(Selector10),
	.datab(Selector91),
	.datac(\register[10][11]~q ),
	.datad(\register[8][11]~q ),
	.cin(gnd),
	.combout(\Mux52~12_combout ),
	.cout());
// synopsys translate_off
defparam \Mux52~12 .lut_mask = 16'hD9C8;
defparam \Mux52~12 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X63_Y40_N20
cycloneive_lcell_comb \Mux52~13 (
// Equation(s):
// \Mux52~13_combout  = (Selector10 & ((\Mux52~12_combout  & (\register[11][11]~q )) # (!\Mux52~12_combout  & ((\register[9][11]~q ))))) # (!Selector10 & (((\Mux52~12_combout ))))

	.dataa(\register[11][11]~q ),
	.datab(Selector10),
	.datac(\register[9][11]~q ),
	.datad(\Mux52~12_combout ),
	.cin(gnd),
	.combout(\Mux52~13_combout ),
	.cout());
// synopsys translate_off
defparam \Mux52~13 .lut_mask = 16'hBBC0;
defparam \Mux52~13 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X66_Y33_N18
cycloneive_lcell_comb \Mux52~16 (
// Equation(s):
// \Mux52~16_combout  = (Selector7 & ((Selector8) # ((\Mux52~13_combout )))) # (!Selector7 & (!Selector8 & (\Mux52~15_combout )))

	.dataa(Selector7),
	.datab(Selector8),
	.datac(\Mux52~15_combout ),
	.datad(\Mux52~13_combout ),
	.cin(gnd),
	.combout(\Mux52~16_combout ),
	.cout());
// synopsys translate_off
defparam \Mux52~16 .lut_mask = 16'hBA98;
defparam \Mux52~16 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y36_N12
cycloneive_lcell_comb \register~85 (
// Equation(s):
// \register~85_combout  = (WideOr01 & ((\wdat[10]~42_combout ) # ((plif_memwbrtnaddr_l_10 & plif_memwbregsrc_l_1))))

	.dataa(plif_memwbrtnaddr_l_10),
	.datab(plif_memwbregsrc_l_1),
	.datac(wdat_10),
	.datad(WideOr0),
	.cin(gnd),
	.combout(\register~85_combout ),
	.cout());
// synopsys translate_off
defparam \register~85 .lut_mask = 16'hF800;
defparam \register~85 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X65_Y38_N8
cycloneive_lcell_comb \register[28][10]~feeder (
// Equation(s):
// \register[28][10]~feeder_combout  = \register~85_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(\register~85_combout ),
	.cin(gnd),
	.combout(\register[28][10]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \register[28][10]~feeder .lut_mask = 16'hFF00;
defparam \register[28][10]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X65_Y38_N9
dffeas \register[28][10] (
	.clk(!CLK),
	.d(\register[28][10]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~57_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\register[28][10]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \register[28][10] .is_wysiwyg = "true";
defparam \register[28][10] .power_up = "low";
// synopsys translate_on

// Location: FF_X65_Y38_N7
dffeas \register[24][10] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\register~85_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~34_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\register[24][10]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \register[24][10] .is_wysiwyg = "true";
defparam \register[24][10] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X66_Y36_N0
cycloneive_lcell_comb \register[16][10]~feeder (
// Equation(s):
// \register[16][10]~feeder_combout  = \register~85_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(\register~85_combout ),
	.datad(gnd),
	.cin(gnd),
	.combout(\register[16][10]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \register[16][10]~feeder .lut_mask = 16'hF0F0;
defparam \register[16][10]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X66_Y36_N1
dffeas \register[16][10] (
	.clk(!CLK),
	.d(\register[16][10]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~36_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\register[16][10]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \register[16][10] .is_wysiwyg = "true";
defparam \register[16][10] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X65_Y38_N6
cycloneive_lcell_comb \Mux53~4 (
// Equation(s):
// \Mux53~4_combout  = (Selector8 & (Selector7)) # (!Selector8 & ((Selector7 & (\register[24][10]~q )) # (!Selector7 & ((\register[16][10]~q )))))

	.dataa(Selector8),
	.datab(Selector7),
	.datac(\register[24][10]~q ),
	.datad(\register[16][10]~q ),
	.cin(gnd),
	.combout(\Mux53~4_combout ),
	.cout());
// synopsys translate_off
defparam \Mux53~4 .lut_mask = 16'hD9C8;
defparam \Mux53~4 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X65_Y38_N26
cycloneive_lcell_comb \Mux53~5 (
// Equation(s):
// \Mux53~5_combout  = (Selector8 & ((\Mux53~4_combout  & ((\register[28][10]~q ))) # (!\Mux53~4_combout  & (\register[20][10]~q )))) # (!Selector8 & (((\Mux53~4_combout ))))

	.dataa(\register[20][10]~q ),
	.datab(Selector8),
	.datac(\register[28][10]~q ),
	.datad(\Mux53~4_combout ),
	.cin(gnd),
	.combout(\Mux53~5_combout ),
	.cout());
// synopsys translate_off
defparam \Mux53~5 .lut_mask = 16'hF388;
defparam \Mux53~5 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X68_Y35_N10
cycloneive_lcell_comb \register[26][10]~feeder (
// Equation(s):
// \register[26][10]~feeder_combout  = \register~85_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(\register~85_combout ),
	.cin(gnd),
	.combout(\register[26][10]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \register[26][10]~feeder .lut_mask = 16'hFF00;
defparam \register[26][10]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X68_Y35_N11
dffeas \register[26][10] (
	.clk(!CLK),
	.d(\register[26][10]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~54_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\register[26][10]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \register[26][10] .is_wysiwyg = "true";
defparam \register[26][10] .power_up = "low";
// synopsys translate_on

// Location: FF_X69_Y35_N31
dffeas \register[18][10] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\register~85_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~33_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\register[18][10]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \register[18][10] .is_wysiwyg = "true";
defparam \register[18][10] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X69_Y35_N30
cycloneive_lcell_comb \Mux53~2 (
// Equation(s):
// \Mux53~2_combout  = (Selector8 & (((Selector7)))) # (!Selector8 & ((Selector7 & (\register[26][10]~q )) # (!Selector7 & ((\register[18][10]~q )))))

	.dataa(Selector8),
	.datab(\register[26][10]~q ),
	.datac(\register[18][10]~q ),
	.datad(Selector7),
	.cin(gnd),
	.combout(\Mux53~2_combout ),
	.cout());
// synopsys translate_off
defparam \Mux53~2 .lut_mask = 16'hEE50;
defparam \Mux53~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X68_Y39_N7
dffeas \register[30][10] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\register~85_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~56_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\register[30][10]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \register[30][10] .is_wysiwyg = "true";
defparam \register[30][10] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X68_Y40_N16
cycloneive_lcell_comb \Mux53~3 (
// Equation(s):
// \Mux53~3_combout  = (Selector8 & ((\Mux53~2_combout  & ((\register[30][10]~q ))) # (!\Mux53~2_combout  & (\register[22][10]~q )))) # (!Selector8 & (((\Mux53~2_combout ))))

	.dataa(\register[22][10]~q ),
	.datab(Selector8),
	.datac(\Mux53~2_combout ),
	.datad(\register[30][10]~q ),
	.cin(gnd),
	.combout(\Mux53~3_combout ),
	.cout());
// synopsys translate_off
defparam \Mux53~3 .lut_mask = 16'hF838;
defparam \Mux53~3 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X68_Y40_N14
cycloneive_lcell_comb \Mux53~6 (
// Equation(s):
// \Mux53~6_combout  = (Selector10 & (Selector91)) # (!Selector10 & ((Selector91 & ((\Mux53~3_combout ))) # (!Selector91 & (\Mux53~5_combout ))))

	.dataa(Selector10),
	.datab(Selector91),
	.datac(\Mux53~5_combout ),
	.datad(\Mux53~3_combout ),
	.cin(gnd),
	.combout(\Mux53~6_combout ),
	.cout());
// synopsys translate_off
defparam \Mux53~6 .lut_mask = 16'hDC98;
defparam \Mux53~6 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X68_Y40_N0
cycloneive_lcell_comb \register[31][10]~feeder (
// Equation(s):
// \register[31][10]~feeder_combout  = \register~85_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(\register~85_combout ),
	.cin(gnd),
	.combout(\register[31][10]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \register[31][10]~feeder .lut_mask = 16'hFF00;
defparam \register[31][10]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X68_Y40_N1
dffeas \register[31][10] (
	.clk(!CLK),
	.d(\register[31][10]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~40_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\register[31][10]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \register[31][10] .is_wysiwyg = "true";
defparam \register[31][10] .power_up = "low";
// synopsys translate_on

// Location: FF_X62_Y38_N29
dffeas \register[23][10] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\register~85_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~37_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\register[23][10]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \register[23][10] .is_wysiwyg = "true";
defparam \register[23][10] .power_up = "low";
// synopsys translate_on

// Location: FF_X62_Y38_N11
dffeas \register[19][10] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\register~85_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~39_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\register[19][10]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \register[19][10] .is_wysiwyg = "true";
defparam \register[19][10] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X62_Y38_N10
cycloneive_lcell_comb \Mux53~7 (
// Equation(s):
// \Mux53~7_combout  = (Selector8 & ((\register[23][10]~q ) # ((Selector7)))) # (!Selector8 & (((\register[19][10]~q  & !Selector7))))

	.dataa(Selector8),
	.datab(\register[23][10]~q ),
	.datac(\register[19][10]~q ),
	.datad(Selector7),
	.cin(gnd),
	.combout(\Mux53~7_combout ),
	.cout());
// synopsys translate_off
defparam \Mux53~7 .lut_mask = 16'hAAD8;
defparam \Mux53~7 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X62_Y39_N9
dffeas \register[27][10] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\register~85_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~38_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\register[27][10]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \register[27][10] .is_wysiwyg = "true";
defparam \register[27][10] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X68_Y40_N26
cycloneive_lcell_comb \Mux53~8 (
// Equation(s):
// \Mux53~8_combout  = (Selector7 & ((\Mux53~7_combout  & (\register[31][10]~q )) # (!\Mux53~7_combout  & ((\register[27][10]~q ))))) # (!Selector7 & (((\Mux53~7_combout ))))

	.dataa(Selector7),
	.datab(\register[31][10]~q ),
	.datac(\Mux53~7_combout ),
	.datad(\register[27][10]~q ),
	.cin(gnd),
	.combout(\Mux53~8_combout ),
	.cout());
// synopsys translate_off
defparam \Mux53~8 .lut_mask = 16'hDAD0;
defparam \Mux53~8 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X61_Y34_N19
dffeas \register[29][10] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\register~85_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~28_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\register[29][10]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \register[29][10] .is_wysiwyg = "true";
defparam \register[29][10] .power_up = "low";
// synopsys translate_on

// Location: FF_X61_Y37_N9
dffeas \register[25][10] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\register~85_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~24_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\register[25][10]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \register[25][10] .is_wysiwyg = "true";
defparam \register[25][10] .power_up = "low";
// synopsys translate_on

// Location: FF_X62_Y33_N23
dffeas \register[21][10] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\register~85_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~22_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\register[21][10]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \register[21][10] .is_wysiwyg = "true";
defparam \register[21][10] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X62_Y33_N22
cycloneive_lcell_comb \Mux53~0 (
// Equation(s):
// \Mux53~0_combout  = (Selector8 & (((\register[21][10]~q ) # (Selector7)))) # (!Selector8 & (\register[17][10]~q  & ((!Selector7))))

	.dataa(\register[17][10]~q ),
	.datab(Selector8),
	.datac(\register[21][10]~q ),
	.datad(Selector7),
	.cin(gnd),
	.combout(\Mux53~0_combout ),
	.cout());
// synopsys translate_off
defparam \Mux53~0 .lut_mask = 16'hCCE2;
defparam \Mux53~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y37_N8
cycloneive_lcell_comb \Mux53~1 (
// Equation(s):
// \Mux53~1_combout  = (Selector7 & ((\Mux53~0_combout  & (\register[29][10]~q )) # (!\Mux53~0_combout  & ((\register[25][10]~q ))))) # (!Selector7 & (((\Mux53~0_combout ))))

	.dataa(Selector7),
	.datab(\register[29][10]~q ),
	.datac(\register[25][10]~q ),
	.datad(\Mux53~0_combout ),
	.cin(gnd),
	.combout(\Mux53~1_combout ),
	.cout());
// synopsys translate_off
defparam \Mux53~1 .lut_mask = 16'hDDA0;
defparam \Mux53~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X63_Y40_N3
dffeas \register[11][10] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\register~85_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~47_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\register[11][10]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \register[11][10] .is_wysiwyg = "true";
defparam \register[11][10] .power_up = "low";
// synopsys translate_on

// Location: FF_X63_Y40_N5
dffeas \register[9][10] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\register~85_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~44_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\register[9][10]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \register[9][10] .is_wysiwyg = "true";
defparam \register[9][10] .power_up = "low";
// synopsys translate_on

// Location: FF_X62_Y41_N15
dffeas \register[8][10] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\register~85_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~46_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\register[8][10]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \register[8][10] .is_wysiwyg = "true";
defparam \register[8][10] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X62_Y41_N14
cycloneive_lcell_comb \Mux53~10 (
// Equation(s):
// \Mux53~10_combout  = (Selector91 & ((\register[10][10]~q ) # ((Selector10)))) # (!Selector91 & (((\register[8][10]~q  & !Selector10))))

	.dataa(\register[10][10]~q ),
	.datab(Selector91),
	.datac(\register[8][10]~q ),
	.datad(Selector10),
	.cin(gnd),
	.combout(\Mux53~10_combout ),
	.cout());
// synopsys translate_off
defparam \Mux53~10 .lut_mask = 16'hCCB8;
defparam \Mux53~10 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X63_Y40_N4
cycloneive_lcell_comb \Mux53~11 (
// Equation(s):
// \Mux53~11_combout  = (Selector10 & ((\Mux53~10_combout  & (\register[11][10]~q )) # (!\Mux53~10_combout  & ((\register[9][10]~q ))))) # (!Selector10 & (((\Mux53~10_combout ))))

	.dataa(Selector10),
	.datab(\register[11][10]~q ),
	.datac(\register[9][10]~q ),
	.datad(\Mux53~10_combout ),
	.cin(gnd),
	.combout(\Mux53~11_combout ),
	.cout());
// synopsys translate_off
defparam \Mux53~11 .lut_mask = 16'hDDA0;
defparam \Mux53~11 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X62_Y36_N13
dffeas \register[15][10] (
	.clk(!CLK),
	.d(\register~85_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~53_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\register[15][10]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \register[15][10] .is_wysiwyg = "true";
defparam \register[15][10] .power_up = "low";
// synopsys translate_on

// Location: FF_X62_Y33_N5
dffeas \register[14][10] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\register~85_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~61_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\register[14][10]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \register[14][10] .is_wysiwyg = "true";
defparam \register[14][10] .power_up = "low";
// synopsys translate_on

// Location: FF_X60_Y33_N31
dffeas \register[12][10] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\register~85_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~52_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\register[12][10]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \register[12][10] .is_wysiwyg = "true";
defparam \register[12][10] .power_up = "low";
// synopsys translate_on

// Location: FF_X60_Y33_N29
dffeas \register[13][10] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\register~85_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~62_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\register[13][10]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \register[13][10] .is_wysiwyg = "true";
defparam \register[13][10] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X60_Y33_N30
cycloneive_lcell_comb \Mux53~17 (
// Equation(s):
// \Mux53~17_combout  = (Selector10 & ((Selector91) # ((\register[13][10]~q )))) # (!Selector10 & (!Selector91 & (\register[12][10]~q )))

	.dataa(Selector10),
	.datab(Selector91),
	.datac(\register[12][10]~q ),
	.datad(\register[13][10]~q ),
	.cin(gnd),
	.combout(\Mux53~17_combout ),
	.cout());
// synopsys translate_off
defparam \Mux53~17 .lut_mask = 16'hBA98;
defparam \Mux53~17 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y33_N4
cycloneive_lcell_comb \Mux53~18 (
// Equation(s):
// \Mux53~18_combout  = (Selector91 & ((\Mux53~17_combout  & (\register[15][10]~q )) # (!\Mux53~17_combout  & ((\register[14][10]~q ))))) # (!Selector91 & (((\Mux53~17_combout ))))

	.dataa(Selector91),
	.datab(\register[15][10]~q ),
	.datac(\register[14][10]~q ),
	.datad(\Mux53~17_combout ),
	.cin(gnd),
	.combout(\Mux53~18_combout ),
	.cout());
// synopsys translate_off
defparam \Mux53~18 .lut_mask = 16'hDDA0;
defparam \Mux53~18 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X65_Y33_N19
dffeas \register[1][10] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\register~85_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~49_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\register[1][10]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \register[1][10] .is_wysiwyg = "true";
defparam \register[1][10] .power_up = "low";
// synopsys translate_on

// Location: FF_X65_Y33_N25
dffeas \register[3][10] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\register~85_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~48_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\register[3][10]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \register[3][10] .is_wysiwyg = "true";
defparam \register[3][10] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X65_Y33_N24
cycloneive_lcell_comb \Mux53~14 (
// Equation(s):
// \Mux53~14_combout  = (Selector10 & ((Selector91 & ((\register[3][10]~q ))) # (!Selector91 & (\register[1][10]~q ))))

	.dataa(Selector91),
	.datab(\register[1][10]~q ),
	.datac(\register[3][10]~q ),
	.datad(Selector10),
	.cin(gnd),
	.combout(\Mux53~14_combout ),
	.cout());
// synopsys translate_off
defparam \Mux53~14 .lut_mask = 16'hE400;
defparam \Mux53~14 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X68_Y33_N21
dffeas \register[2][10] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\register~85_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~50_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\register[2][10]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \register[2][10] .is_wysiwyg = "true";
defparam \register[2][10] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X68_Y33_N20
cycloneive_lcell_comb \Mux53~15 (
// Equation(s):
// \Mux53~15_combout  = (\Mux53~14_combout ) # ((Selector91 & (\register[2][10]~q  & !Selector10)))

	.dataa(Selector91),
	.datab(\Mux53~14_combout ),
	.datac(\register[2][10]~q ),
	.datad(Selector10),
	.cin(gnd),
	.combout(\Mux53~15_combout ),
	.cout());
// synopsys translate_off
defparam \Mux53~15 .lut_mask = 16'hCCEC;
defparam \Mux53~15 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X67_Y32_N3
dffeas \register[4][10] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\register~85_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~60_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\register[4][10]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \register[4][10] .is_wysiwyg = "true";
defparam \register[4][10] .power_up = "low";
// synopsys translate_on

// Location: FF_X67_Y32_N1
dffeas \register[5][10] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\register~85_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~59_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\register[5][10]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \register[5][10] .is_wysiwyg = "true";
defparam \register[5][10] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X67_Y32_N2
cycloneive_lcell_comb \Mux53~12 (
// Equation(s):
// \Mux53~12_combout  = (Selector10 & ((Selector91) # ((\register[5][10]~q )))) # (!Selector10 & (!Selector91 & (\register[4][10]~q )))

	.dataa(Selector10),
	.datab(Selector91),
	.datac(\register[4][10]~q ),
	.datad(\register[5][10]~q ),
	.cin(gnd),
	.combout(\Mux53~12_combout ),
	.cout());
// synopsys translate_off
defparam \Mux53~12 .lut_mask = 16'hBA98;
defparam \Mux53~12 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X68_Y33_N28
cycloneive_lcell_comb \register[7][10]~feeder (
// Equation(s):
// \register[7][10]~feeder_combout  = \register~85_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(\register~85_combout ),
	.datad(gnd),
	.cin(gnd),
	.combout(\register[7][10]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \register[7][10]~feeder .lut_mask = 16'hF0F0;
defparam \register[7][10]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X68_Y33_N29
dffeas \register[7][10] (
	.clk(!CLK),
	.d(\register[7][10]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~43_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\register[7][10]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \register[7][10] .is_wysiwyg = "true";
defparam \register[7][10] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X68_Y33_N2
cycloneive_lcell_comb \Mux53~13 (
// Equation(s):
// \Mux53~13_combout  = (\Mux53~12_combout  & (((\register[7][10]~q ) # (!Selector91)))) # (!\Mux53~12_combout  & (\register[6][10]~q  & (Selector91)))

	.dataa(\register[6][10]~q ),
	.datab(\Mux53~12_combout ),
	.datac(Selector91),
	.datad(\register[7][10]~q ),
	.cin(gnd),
	.combout(\Mux53~13_combout ),
	.cout());
// synopsys translate_off
defparam \Mux53~13 .lut_mask = 16'hEC2C;
defparam \Mux53~13 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X68_Y40_N6
cycloneive_lcell_comb \Mux53~16 (
// Equation(s):
// \Mux53~16_combout  = (Selector7 & (Selector8)) # (!Selector7 & ((Selector8 & ((\Mux53~13_combout ))) # (!Selector8 & (\Mux53~15_combout ))))

	.dataa(Selector7),
	.datab(Selector8),
	.datac(\Mux53~15_combout ),
	.datad(\Mux53~13_combout ),
	.cin(gnd),
	.combout(\Mux53~16_combout ),
	.cout());
// synopsys translate_off
defparam \Mux53~16 .lut_mask = 16'hDC98;
defparam \Mux53~16 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y35_N4
cycloneive_lcell_comb \register~86 (
// Equation(s):
// \register~86_combout  = (WideOr01 & ((\wdat[9]~44_combout ) # ((plif_memwbregsrc_l_1 & plif_memwbrtnaddr_l_9))))

	.dataa(WideOr0),
	.datab(plif_memwbregsrc_l_1),
	.datac(plif_memwbrtnaddr_l_9),
	.datad(wdat_9),
	.cin(gnd),
	.combout(\register~86_combout ),
	.cout());
// synopsys translate_off
defparam \register~86 .lut_mask = 16'hAA80;
defparam \register~86 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X69_Y36_N18
cycloneive_lcell_comb \register[28][9]~feeder (
// Equation(s):
// \register[28][9]~feeder_combout  = \register~86_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(\register~86_combout ),
	.cin(gnd),
	.combout(\register[28][9]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \register[28][9]~feeder .lut_mask = 16'hFF00;
defparam \register[28][9]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X69_Y36_N19
dffeas \register[28][9] (
	.clk(!CLK),
	.d(\register[28][9]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~57_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\register[28][9]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \register[28][9] .is_wysiwyg = "true";
defparam \register[28][9] .power_up = "low";
// synopsys translate_on

// Location: FF_X65_Y39_N19
dffeas \register[20][9] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\register~86_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~35_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\register[20][9]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \register[20][9] .is_wysiwyg = "true";
defparam \register[20][9] .power_up = "low";
// synopsys translate_on

// Location: FF_X65_Y39_N13
dffeas \register[16][9] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\register~86_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~36_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\register[16][9]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \register[16][9] .is_wysiwyg = "true";
defparam \register[16][9] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X65_Y39_N18
cycloneive_lcell_comb \Mux54~4 (
// Equation(s):
// \Mux54~4_combout  = (Selector7 & (Selector8)) # (!Selector7 & ((Selector8 & (\register[20][9]~q )) # (!Selector8 & ((\register[16][9]~q )))))

	.dataa(Selector7),
	.datab(Selector8),
	.datac(\register[20][9]~q ),
	.datad(\register[16][9]~q ),
	.cin(gnd),
	.combout(\Mux54~4_combout ),
	.cout());
// synopsys translate_off
defparam \Mux54~4 .lut_mask = 16'hD9C8;
defparam \Mux54~4 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X69_Y36_N0
cycloneive_lcell_comb \Mux54~5 (
// Equation(s):
// \Mux54~5_combout  = (\Mux54~4_combout  & (((\register[28][9]~q ) # (!Selector7)))) # (!\Mux54~4_combout  & (\register[24][9]~q  & ((Selector7))))

	.dataa(\register[24][9]~q ),
	.datab(\register[28][9]~q ),
	.datac(\Mux54~4_combout ),
	.datad(Selector7),
	.cin(gnd),
	.combout(\Mux54~5_combout ),
	.cout());
// synopsys translate_off
defparam \Mux54~5 .lut_mask = 16'hCAF0;
defparam \Mux54~5 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X69_Y37_N5
dffeas \register[18][9] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\register~86_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~33_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\register[18][9]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \register[18][9] .is_wysiwyg = "true";
defparam \register[18][9] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X69_Y37_N4
cycloneive_lcell_comb \Mux54~2 (
// Equation(s):
// \Mux54~2_combout  = (Selector8 & ((\register[22][9]~q ) # ((Selector7)))) # (!Selector8 & (((\register[18][9]~q  & !Selector7))))

	.dataa(\register[22][9]~q ),
	.datab(Selector8),
	.datac(\register[18][9]~q ),
	.datad(Selector7),
	.cin(gnd),
	.combout(\Mux54~2_combout ),
	.cout());
// synopsys translate_off
defparam \Mux54~2 .lut_mask = 16'hCCB8;
defparam \Mux54~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X68_Y37_N17
dffeas \register[26][9] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\register~86_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~54_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\register[26][9]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \register[26][9] .is_wysiwyg = "true";
defparam \register[26][9] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X69_Y36_N16
cycloneive_lcell_comb \Mux54~3 (
// Equation(s):
// \Mux54~3_combout  = (\Mux54~2_combout  & ((\register[30][9]~q ) # ((!Selector7)))) # (!\Mux54~2_combout  & (((\register[26][9]~q  & Selector7))))

	.dataa(\register[30][9]~q ),
	.datab(\Mux54~2_combout ),
	.datac(\register[26][9]~q ),
	.datad(Selector7),
	.cin(gnd),
	.combout(\Mux54~3_combout ),
	.cout());
// synopsys translate_off
defparam \Mux54~3 .lut_mask = 16'hB8CC;
defparam \Mux54~3 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X69_Y36_N14
cycloneive_lcell_comb \Mux54~6 (
// Equation(s):
// \Mux54~6_combout  = (Selector10 & (((Selector91)))) # (!Selector10 & ((Selector91 & ((\Mux54~3_combout ))) # (!Selector91 & (\Mux54~5_combout ))))

	.dataa(Selector10),
	.datab(\Mux54~5_combout ),
	.datac(Selector91),
	.datad(\Mux54~3_combout ),
	.cin(gnd),
	.combout(\Mux54~6_combout ),
	.cout());
// synopsys translate_off
defparam \Mux54~6 .lut_mask = 16'hF4A4;
defparam \Mux54~6 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X60_Y35_N27
dffeas \register[23][9] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\register~86_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~37_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\register[23][9]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \register[23][9] .is_wysiwyg = "true";
defparam \register[23][9] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X68_Y40_N18
cycloneive_lcell_comb \register[31][9]~feeder (
// Equation(s):
// \register[31][9]~feeder_combout  = \register~86_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(\register~86_combout ),
	.cin(gnd),
	.combout(\register[31][9]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \register[31][9]~feeder .lut_mask = 16'hFF00;
defparam \register[31][9]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X68_Y40_N19
dffeas \register[31][9] (
	.clk(!CLK),
	.d(\register[31][9]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~40_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\register[31][9]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \register[31][9] .is_wysiwyg = "true";
defparam \register[31][9] .power_up = "low";
// synopsys translate_on

// Location: FF_X60_Y35_N17
dffeas \register[19][9] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\register~86_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~39_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\register[19][9]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \register[19][9] .is_wysiwyg = "true";
defparam \register[19][9] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X57_Y41_N8
cycloneive_lcell_comb \register[27][9]~feeder (
// Equation(s):
// \register[27][9]~feeder_combout  = \register~86_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(\register~86_combout ),
	.cin(gnd),
	.combout(\register[27][9]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \register[27][9]~feeder .lut_mask = 16'hFF00;
defparam \register[27][9]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X57_Y41_N9
dffeas \register[27][9] (
	.clk(!CLK),
	.d(\register[27][9]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~38_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\register[27][9]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \register[27][9] .is_wysiwyg = "true";
defparam \register[27][9] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X60_Y35_N16
cycloneive_lcell_comb \Mux54~7 (
// Equation(s):
// \Mux54~7_combout  = (Selector7 & ((Selector8) # ((\register[27][9]~q )))) # (!Selector7 & (!Selector8 & (\register[19][9]~q )))

	.dataa(Selector7),
	.datab(Selector8),
	.datac(\register[19][9]~q ),
	.datad(\register[27][9]~q ),
	.cin(gnd),
	.combout(\Mux54~7_combout ),
	.cout());
// synopsys translate_off
defparam \Mux54~7 .lut_mask = 16'hBA98;
defparam \Mux54~7 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X68_Y40_N4
cycloneive_lcell_comb \Mux54~8 (
// Equation(s):
// \Mux54~8_combout  = (Selector8 & ((\Mux54~7_combout  & ((\register[31][9]~q ))) # (!\Mux54~7_combout  & (\register[23][9]~q )))) # (!Selector8 & (((\Mux54~7_combout ))))

	.dataa(\register[23][9]~q ),
	.datab(\register[31][9]~q ),
	.datac(Selector8),
	.datad(\Mux54~7_combout ),
	.cin(gnd),
	.combout(\Mux54~8_combout ),
	.cout());
// synopsys translate_off
defparam \Mux54~8 .lut_mask = 16'hCFA0;
defparam \Mux54~8 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X61_Y34_N31
dffeas \register[29][9] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\register~86_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~28_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\register[29][9]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \register[29][9] .is_wysiwyg = "true";
defparam \register[29][9] .power_up = "low";
// synopsys translate_on

// Location: FF_X61_Y37_N19
dffeas \register[25][9] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\register~86_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~24_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\register[25][9]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \register[25][9] .is_wysiwyg = "true";
defparam \register[25][9] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X61_Y37_N18
cycloneive_lcell_comb \Mux54~0 (
// Equation(s):
// \Mux54~0_combout  = (Selector8 & (((Selector7)))) # (!Selector8 & ((Selector7 & ((\register[25][9]~q ))) # (!Selector7 & (\register[17][9]~q ))))

	.dataa(\register[17][9]~q ),
	.datab(Selector8),
	.datac(\register[25][9]~q ),
	.datad(Selector7),
	.cin(gnd),
	.combout(\Mux54~0_combout ),
	.cout());
// synopsys translate_off
defparam \Mux54~0 .lut_mask = 16'hFC22;
defparam \Mux54~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y34_N16
cycloneive_lcell_comb \register[21][9]~feeder (
// Equation(s):
// \register[21][9]~feeder_combout  = \register~86_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(\register~86_combout ),
	.datad(gnd),
	.cin(gnd),
	.combout(\register[21][9]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \register[21][9]~feeder .lut_mask = 16'hF0F0;
defparam \register[21][9]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X61_Y34_N17
dffeas \register[21][9] (
	.clk(!CLK),
	.d(\register[21][9]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~22_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\register[21][9]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \register[21][9] .is_wysiwyg = "true";
defparam \register[21][9] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X61_Y34_N24
cycloneive_lcell_comb \Mux54~1 (
// Equation(s):
// \Mux54~1_combout  = (Selector8 & ((\Mux54~0_combout  & (\register[29][9]~q )) # (!\Mux54~0_combout  & ((\register[21][9]~q ))))) # (!Selector8 & (((\Mux54~0_combout ))))

	.dataa(\register[29][9]~q ),
	.datab(Selector8),
	.datac(\Mux54~0_combout ),
	.datad(\register[21][9]~q ),
	.cin(gnd),
	.combout(\Mux54~1_combout ),
	.cout());
// synopsys translate_off
defparam \Mux54~1 .lut_mask = 16'hBCB0;
defparam \Mux54~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X61_Y35_N5
dffeas \register[15][9] (
	.clk(!CLK),
	.d(\register~86_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~53_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\register[15][9]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \register[15][9] .is_wysiwyg = "true";
defparam \register[15][9] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X67_Y33_N20
cycloneive_lcell_comb \register[14][9]~feeder (
// Equation(s):
// \register[14][9]~feeder_combout  = \register~86_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(\register~86_combout ),
	.cin(gnd),
	.combout(\register[14][9]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \register[14][9]~feeder .lut_mask = 16'hFF00;
defparam \register[14][9]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X67_Y33_N21
dffeas \register[14][9] (
	.clk(!CLK),
	.d(\register[14][9]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~61_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\register[14][9]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \register[14][9] .is_wysiwyg = "true";
defparam \register[14][9] .power_up = "low";
// synopsys translate_on

// Location: FF_X60_Y33_N15
dffeas \register[12][9] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\register~86_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~52_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\register[12][9]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \register[12][9] .is_wysiwyg = "true";
defparam \register[12][9] .power_up = "low";
// synopsys translate_on

// Location: FF_X60_Y33_N25
dffeas \register[13][9] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\register~86_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~62_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\register[13][9]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \register[13][9] .is_wysiwyg = "true";
defparam \register[13][9] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X60_Y33_N14
cycloneive_lcell_comb \Mux54~17 (
// Equation(s):
// \Mux54~17_combout  = (Selector10 & ((Selector91) # ((\register[13][9]~q )))) # (!Selector10 & (!Selector91 & (\register[12][9]~q )))

	.dataa(Selector10),
	.datab(Selector91),
	.datac(\register[12][9]~q ),
	.datad(\register[13][9]~q ),
	.cin(gnd),
	.combout(\Mux54~17_combout ),
	.cout());
// synopsys translate_off
defparam \Mux54~17 .lut_mask = 16'hBA98;
defparam \Mux54~17 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X67_Y33_N14
cycloneive_lcell_comb \Mux54~18 (
// Equation(s):
// \Mux54~18_combout  = (\Mux54~17_combout  & ((\register[15][9]~q ) # ((!Selector91)))) # (!\Mux54~17_combout  & (((\register[14][9]~q  & Selector91))))

	.dataa(\register[15][9]~q ),
	.datab(\register[14][9]~q ),
	.datac(\Mux54~17_combout ),
	.datad(Selector91),
	.cin(gnd),
	.combout(\Mux54~18_combout ),
	.cout());
// synopsys translate_off
defparam \Mux54~18 .lut_mask = 16'hACF0;
defparam \Mux54~18 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X67_Y33_N30
cycloneive_lcell_comb \register[6][9]~feeder (
// Equation(s):
// \register[6][9]~feeder_combout  = \register~86_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(\register~86_combout ),
	.cin(gnd),
	.combout(\register[6][9]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \register[6][9]~feeder .lut_mask = 16'hFF00;
defparam \register[6][9]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X67_Y33_N31
dffeas \register[6][9] (
	.clk(!CLK),
	.d(\register[6][9]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~58_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\register[6][9]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \register[6][9] .is_wysiwyg = "true";
defparam \register[6][9] .power_up = "low";
// synopsys translate_on

// Location: FF_X67_Y32_N27
dffeas \register[4][9] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\register~86_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~60_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\register[4][9]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \register[4][9] .is_wysiwyg = "true";
defparam \register[4][9] .power_up = "low";
// synopsys translate_on

// Location: FF_X67_Y32_N25
dffeas \register[5][9] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\register~86_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~59_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\register[5][9]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \register[5][9] .is_wysiwyg = "true";
defparam \register[5][9] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X67_Y32_N26
cycloneive_lcell_comb \Mux54~10 (
// Equation(s):
// \Mux54~10_combout  = (Selector10 & ((Selector91) # ((\register[5][9]~q )))) # (!Selector10 & (!Selector91 & (\register[4][9]~q )))

	.dataa(Selector10),
	.datab(Selector91),
	.datac(\register[4][9]~q ),
	.datad(\register[5][9]~q ),
	.cin(gnd),
	.combout(\Mux54~10_combout ),
	.cout());
// synopsys translate_off
defparam \Mux54~10 .lut_mask = 16'hBA98;
defparam \Mux54~10 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X68_Y33_N19
dffeas \register[7][9] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\register~86_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~43_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\register[7][9]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \register[7][9] .is_wysiwyg = "true";
defparam \register[7][9] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X68_Y33_N16
cycloneive_lcell_comb \Mux54~11 (
// Equation(s):
// \Mux54~11_combout  = (Selector91 & ((\Mux54~10_combout  & ((\register[7][9]~q ))) # (!\Mux54~10_combout  & (\register[6][9]~q )))) # (!Selector91 & (((\Mux54~10_combout ))))

	.dataa(Selector91),
	.datab(\register[6][9]~q ),
	.datac(\Mux54~10_combout ),
	.datad(\register[7][9]~q ),
	.cin(gnd),
	.combout(\Mux54~11_combout ),
	.cout());
// synopsys translate_off
defparam \Mux54~11 .lut_mask = 16'hF858;
defparam \Mux54~11 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X66_Y38_N6
cycloneive_lcell_comb \register[11][9]~feeder (
// Equation(s):
// \register[11][9]~feeder_combout  = \register~86_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(\register~86_combout ),
	.cin(gnd),
	.combout(\register[11][9]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \register[11][9]~feeder .lut_mask = 16'hFF00;
defparam \register[11][9]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X66_Y38_N7
dffeas \register[11][9] (
	.clk(!CLK),
	.d(\register[11][9]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~47_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\register[11][9]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \register[11][9] .is_wysiwyg = "true";
defparam \register[11][9] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X66_Y38_N12
cycloneive_lcell_comb \register[9][9]~feeder (
// Equation(s):
// \register[9][9]~feeder_combout  = \register~86_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(\register~86_combout ),
	.cin(gnd),
	.combout(\register[9][9]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \register[9][9]~feeder .lut_mask = 16'hFF00;
defparam \register[9][9]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X66_Y38_N13
dffeas \register[9][9] (
	.clk(!CLK),
	.d(\register[9][9]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~44_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\register[9][9]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \register[9][9] .is_wysiwyg = "true";
defparam \register[9][9] .power_up = "low";
// synopsys translate_on

// Location: FF_X62_Y41_N7
dffeas \register[8][9] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\register~86_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~46_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\register[8][9]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \register[8][9] .is_wysiwyg = "true";
defparam \register[8][9] .power_up = "low";
// synopsys translate_on

// Location: FF_X62_Y41_N29
dffeas \register[10][9] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\register~86_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~45_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\register[10][9]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \register[10][9] .is_wysiwyg = "true";
defparam \register[10][9] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X62_Y41_N6
cycloneive_lcell_comb \Mux54~12 (
// Equation(s):
// \Mux54~12_combout  = (Selector10 & (Selector91)) # (!Selector10 & ((Selector91 & ((\register[10][9]~q ))) # (!Selector91 & (\register[8][9]~q ))))

	.dataa(Selector10),
	.datab(Selector91),
	.datac(\register[8][9]~q ),
	.datad(\register[10][9]~q ),
	.cin(gnd),
	.combout(\Mux54~12_combout ),
	.cout());
// synopsys translate_off
defparam \Mux54~12 .lut_mask = 16'hDC98;
defparam \Mux54~12 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X67_Y41_N12
cycloneive_lcell_comb \Mux54~13 (
// Equation(s):
// \Mux54~13_combout  = (Selector10 & ((\Mux54~12_combout  & (\register[11][9]~q )) # (!\Mux54~12_combout  & ((\register[9][9]~q ))))) # (!Selector10 & (((\Mux54~12_combout ))))

	.dataa(Selector10),
	.datab(\register[11][9]~q ),
	.datac(\register[9][9]~q ),
	.datad(\Mux54~12_combout ),
	.cin(gnd),
	.combout(\Mux54~13_combout ),
	.cout());
// synopsys translate_off
defparam \Mux54~13 .lut_mask = 16'hDDA0;
defparam \Mux54~13 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X69_Y33_N11
dffeas \register[1][9] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\register~86_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~49_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\register[1][9]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \register[1][9] .is_wysiwyg = "true";
defparam \register[1][9] .power_up = "low";
// synopsys translate_on

// Location: FF_X69_Y33_N29
dffeas \register[3][9] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\register~86_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~48_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\register[3][9]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \register[3][9] .is_wysiwyg = "true";
defparam \register[3][9] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X69_Y33_N10
cycloneive_lcell_comb \Mux54~14 (
// Equation(s):
// \Mux54~14_combout  = (Selector9 & ((plif_ifidinstr_l_17 & ((\register[3][9]~q ))) # (!plif_ifidinstr_l_17 & (\register[1][9]~q )))) # (!Selector9 & (((\register[1][9]~q ))))

	.dataa(Selector9),
	.datab(plif_ifidinstr_l_17),
	.datac(\register[1][9]~q ),
	.datad(\register[3][9]~q ),
	.cin(gnd),
	.combout(\Mux54~14_combout ),
	.cout());
// synopsys translate_off
defparam \Mux54~14 .lut_mask = 16'hF870;
defparam \Mux54~14 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X68_Y33_N7
dffeas \register[2][9] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\register~86_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~50_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\register[2][9]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \register[2][9] .is_wysiwyg = "true";
defparam \register[2][9] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X68_Y33_N6
cycloneive_lcell_comb \Mux54~15 (
// Equation(s):
// \Mux54~15_combout  = (Selector10 & (((\Mux54~14_combout )))) # (!Selector10 & (Selector91 & ((\register[2][9]~q ))))

	.dataa(Selector91),
	.datab(\Mux54~14_combout ),
	.datac(\register[2][9]~q ),
	.datad(Selector10),
	.cin(gnd),
	.combout(\Mux54~15_combout ),
	.cout());
// synopsys translate_off
defparam \Mux54~15 .lut_mask = 16'hCCA0;
defparam \Mux54~15 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X68_Y40_N24
cycloneive_lcell_comb \Mux54~16 (
// Equation(s):
// \Mux54~16_combout  = (Selector7 & ((\Mux54~13_combout ) # ((Selector8)))) # (!Selector7 & (((!Selector8 & \Mux54~15_combout ))))

	.dataa(Selector7),
	.datab(\Mux54~13_combout ),
	.datac(Selector8),
	.datad(\Mux54~15_combout ),
	.cin(gnd),
	.combout(\Mux54~16_combout ),
	.cout());
// synopsys translate_off
defparam \Mux54~16 .lut_mask = 16'hADA8;
defparam \Mux54~16 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X63_Y37_N2
cycloneive_lcell_comb \register~87 (
// Equation(s):
// \register~87_combout  = (WideOr01 & ((\wdat[8]~46_combout ) # ((plif_memwbrtnaddr_l_8 & plif_memwbregsrc_l_1))))

	.dataa(WideOr0),
	.datab(plif_memwbrtnaddr_l_8),
	.datac(wdat_8),
	.datad(plif_memwbregsrc_l_1),
	.cin(gnd),
	.combout(\register~87_combout ),
	.cout());
// synopsys translate_off
defparam \register~87 .lut_mask = 16'hA8A0;
defparam \register~87 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X63_Y33_N8
cycloneive_lcell_comb \register[29][8]~feeder (
// Equation(s):
// \register[29][8]~feeder_combout  = \register~87_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(\register~87_combout ),
	.datad(gnd),
	.cin(gnd),
	.combout(\register[29][8]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \register[29][8]~feeder .lut_mask = 16'hF0F0;
defparam \register[29][8]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X63_Y33_N9
dffeas \register[29][8] (
	.clk(!CLK),
	.d(\register[29][8]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~28_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\register[29][8]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \register[29][8] .is_wysiwyg = "true";
defparam \register[29][8] .power_up = "low";
// synopsys translate_on

// Location: FF_X62_Y36_N31
dffeas \register[25][8] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\register~87_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~24_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\register[25][8]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \register[25][8] .is_wysiwyg = "true";
defparam \register[25][8] .power_up = "low";
// synopsys translate_on

// Location: FF_X63_Y35_N13
dffeas \register[21][8] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\register~87_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~22_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\register[21][8]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \register[21][8] .is_wysiwyg = "true";
defparam \register[21][8] .power_up = "low";
// synopsys translate_on

// Location: FF_X62_Y35_N1
dffeas \register[17][8] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\register~87_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~26_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\register[17][8]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \register[17][8] .is_wysiwyg = "true";
defparam \register[17][8] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X63_Y35_N12
cycloneive_lcell_comb \Mux55~0 (
// Equation(s):
// \Mux55~0_combout  = (Selector7 & (Selector8)) # (!Selector7 & ((Selector8 & (\register[21][8]~q )) # (!Selector8 & ((\register[17][8]~q )))))

	.dataa(Selector7),
	.datab(Selector8),
	.datac(\register[21][8]~q ),
	.datad(\register[17][8]~q ),
	.cin(gnd),
	.combout(\Mux55~0_combout ),
	.cout());
// synopsys translate_off
defparam \Mux55~0 .lut_mask = 16'hD9C8;
defparam \Mux55~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y36_N30
cycloneive_lcell_comb \Mux55~1 (
// Equation(s):
// \Mux55~1_combout  = (Selector7 & ((\Mux55~0_combout  & (\register[29][8]~q )) # (!\Mux55~0_combout  & ((\register[25][8]~q ))))) # (!Selector7 & (((\Mux55~0_combout ))))

	.dataa(\register[29][8]~q ),
	.datab(Selector7),
	.datac(\register[25][8]~q ),
	.datad(\Mux55~0_combout ),
	.cin(gnd),
	.combout(\Mux55~1_combout ),
	.cout());
// synopsys translate_off
defparam \Mux55~1 .lut_mask = 16'hBBC0;
defparam \Mux55~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X69_Y37_N26
cycloneive_lcell_comb \register[22][8]~feeder (
// Equation(s):
// \register[22][8]~feeder_combout  = \register~87_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(\register~87_combout ),
	.cin(gnd),
	.combout(\register[22][8]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \register[22][8]~feeder .lut_mask = 16'hFF00;
defparam \register[22][8]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X69_Y37_N27
dffeas \register[22][8] (
	.clk(!CLK),
	.d(\register[22][8]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~55_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\register[22][8]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \register[22][8] .is_wysiwyg = "true";
defparam \register[22][8] .power_up = "low";
// synopsys translate_on

// Location: FF_X68_Y37_N5
dffeas \register[30][8] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\register~87_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~56_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\register[30][8]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \register[30][8] .is_wysiwyg = "true";
defparam \register[30][8] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X68_Y37_N4
cycloneive_lcell_comb \Mux55~3 (
// Equation(s):
// \Mux55~3_combout  = (\Mux55~2_combout  & (((\register[30][8]~q ) # (!Selector8)))) # (!\Mux55~2_combout  & (\register[22][8]~q  & ((Selector8))))

	.dataa(\Mux55~2_combout ),
	.datab(\register[22][8]~q ),
	.datac(\register[30][8]~q ),
	.datad(Selector8),
	.cin(gnd),
	.combout(\Mux55~3_combout ),
	.cout());
// synopsys translate_off
defparam \Mux55~3 .lut_mask = 16'hE4AA;
defparam \Mux55~3 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X69_Y36_N13
dffeas \register[28][8] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\register~87_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~57_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\register[28][8]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \register[28][8] .is_wysiwyg = "true";
defparam \register[28][8] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X70_Y38_N4
cycloneive_lcell_comb \register[24][8]~feeder (
// Equation(s):
// \register[24][8]~feeder_combout  = \register~87_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(\register~87_combout ),
	.cin(gnd),
	.combout(\register[24][8]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \register[24][8]~feeder .lut_mask = 16'hFF00;
defparam \register[24][8]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X70_Y38_N5
dffeas \register[24][8] (
	.clk(!CLK),
	.d(\register[24][8]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~34_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\register[24][8]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \register[24][8] .is_wysiwyg = "true";
defparam \register[24][8] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X70_Y39_N20
cycloneive_lcell_comb \register[16][8]~feeder (
// Equation(s):
// \register[16][8]~feeder_combout  = \register~87_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(\register~87_combout ),
	.cin(gnd),
	.combout(\register[16][8]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \register[16][8]~feeder .lut_mask = 16'hFF00;
defparam \register[16][8]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X70_Y39_N21
dffeas \register[16][8] (
	.clk(!CLK),
	.d(\register[16][8]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~36_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\register[16][8]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \register[16][8] .is_wysiwyg = "true";
defparam \register[16][8] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X70_Y38_N10
cycloneive_lcell_comb \Mux55~4 (
// Equation(s):
// \Mux55~4_combout  = (Selector7 & ((Selector8) # ((\register[24][8]~q )))) # (!Selector7 & (!Selector8 & ((\register[16][8]~q ))))

	.dataa(Selector7),
	.datab(Selector8),
	.datac(\register[24][8]~q ),
	.datad(\register[16][8]~q ),
	.cin(gnd),
	.combout(\Mux55~4_combout ),
	.cout());
// synopsys translate_off
defparam \Mux55~4 .lut_mask = 16'hB9A8;
defparam \Mux55~4 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X69_Y36_N12
cycloneive_lcell_comb \Mux55~5 (
// Equation(s):
// \Mux55~5_combout  = (Selector8 & ((\Mux55~4_combout  & ((\register[28][8]~q ))) # (!\Mux55~4_combout  & (\register[20][8]~q )))) # (!Selector8 & (((\Mux55~4_combout ))))

	.dataa(\register[20][8]~q ),
	.datab(Selector8),
	.datac(\register[28][8]~q ),
	.datad(\Mux55~4_combout ),
	.cin(gnd),
	.combout(\Mux55~5_combout ),
	.cout());
// synopsys translate_off
defparam \Mux55~5 .lut_mask = 16'hF388;
defparam \Mux55~5 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X69_Y36_N26
cycloneive_lcell_comb \Mux55~6 (
// Equation(s):
// \Mux55~6_combout  = (Selector10 & (Selector91)) # (!Selector10 & ((Selector91 & (\Mux55~3_combout )) # (!Selector91 & ((\Mux55~5_combout )))))

	.dataa(Selector10),
	.datab(Selector91),
	.datac(\Mux55~3_combout ),
	.datad(\Mux55~5_combout ),
	.cin(gnd),
	.combout(\Mux55~6_combout ),
	.cout());
// synopsys translate_off
defparam \Mux55~6 .lut_mask = 16'hD9C8;
defparam \Mux55~6 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X62_Y39_N31
dffeas \register[27][8] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\register~87_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~38_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\register[27][8]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \register[27][8] .is_wysiwyg = "true";
defparam \register[27][8] .power_up = "low";
// synopsys translate_on

// Location: FF_X62_Y39_N13
dffeas \register[31][8] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\register~87_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~40_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\register[31][8]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \register[31][8] .is_wysiwyg = "true";
defparam \register[31][8] .power_up = "low";
// synopsys translate_on

// Location: FF_X62_Y38_N27
dffeas \register[19][8] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\register~87_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~39_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\register[19][8]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \register[19][8] .is_wysiwyg = "true";
defparam \register[19][8] .power_up = "low";
// synopsys translate_on

// Location: FF_X62_Y38_N13
dffeas \register[23][8] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\register~87_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~37_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\register[23][8]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \register[23][8] .is_wysiwyg = "true";
defparam \register[23][8] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X62_Y38_N26
cycloneive_lcell_comb \Mux55~7 (
// Equation(s):
// \Mux55~7_combout  = (Selector7 & (Selector8)) # (!Selector7 & ((Selector8 & ((\register[23][8]~q ))) # (!Selector8 & (\register[19][8]~q ))))

	.dataa(Selector7),
	.datab(Selector8),
	.datac(\register[19][8]~q ),
	.datad(\register[23][8]~q ),
	.cin(gnd),
	.combout(\Mux55~7_combout ),
	.cout());
// synopsys translate_off
defparam \Mux55~7 .lut_mask = 16'hDC98;
defparam \Mux55~7 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y39_N12
cycloneive_lcell_comb \Mux55~8 (
// Equation(s):
// \Mux55~8_combout  = (Selector7 & ((\Mux55~7_combout  & ((\register[31][8]~q ))) # (!\Mux55~7_combout  & (\register[27][8]~q )))) # (!Selector7 & (((\Mux55~7_combout ))))

	.dataa(\register[27][8]~q ),
	.datab(Selector7),
	.datac(\register[31][8]~q ),
	.datad(\Mux55~7_combout ),
	.cin(gnd),
	.combout(\Mux55~8_combout ),
	.cout());
// synopsys translate_off
defparam \Mux55~8 .lut_mask = 16'hF388;
defparam \Mux55~8 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X60_Y33_N9
dffeas \register[13][8] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\register~87_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~62_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\register[13][8]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \register[13][8] .is_wysiwyg = "true";
defparam \register[13][8] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X60_Y33_N8
cycloneive_lcell_comb \Mux55~17 (
// Equation(s):
// \Mux55~17_combout  = (Selector10 & (((\register[13][8]~q ) # (Selector91)))) # (!Selector10 & (\register[12][8]~q  & ((!Selector91))))

	.dataa(\register[12][8]~q ),
	.datab(Selector10),
	.datac(\register[13][8]~q ),
	.datad(Selector91),
	.cin(gnd),
	.combout(\Mux55~17_combout ),
	.cout());
// synopsys translate_off
defparam \Mux55~17 .lut_mask = 16'hCCE2;
defparam \Mux55~17 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X67_Y33_N8
cycloneive_lcell_comb \register[14][8]~feeder (
// Equation(s):
// \register[14][8]~feeder_combout  = \register~87_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(\register~87_combout ),
	.datad(gnd),
	.cin(gnd),
	.combout(\register[14][8]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \register[14][8]~feeder .lut_mask = 16'hF0F0;
defparam \register[14][8]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X67_Y33_N9
dffeas \register[14][8] (
	.clk(!CLK),
	.d(\register[14][8]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~61_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\register[14][8]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \register[14][8] .is_wysiwyg = "true";
defparam \register[14][8] .power_up = "low";
// synopsys translate_on

// Location: FF_X63_Y37_N3
dffeas \register[15][8] (
	.clk(!CLK),
	.d(\register~87_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~53_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\register[15][8]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \register[15][8] .is_wysiwyg = "true";
defparam \register[15][8] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X66_Y33_N16
cycloneive_lcell_comb \Mux55~18 (
// Equation(s):
// \Mux55~18_combout  = (\Mux55~17_combout  & (((\register[15][8]~q ) # (!Selector91)))) # (!\Mux55~17_combout  & (\register[14][8]~q  & ((Selector91))))

	.dataa(\Mux55~17_combout ),
	.datab(\register[14][8]~q ),
	.datac(\register[15][8]~q ),
	.datad(Selector91),
	.cin(gnd),
	.combout(\Mux55~18_combout ),
	.cout());
// synopsys translate_off
defparam \Mux55~18 .lut_mask = 16'hE4AA;
defparam \Mux55~18 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X67_Y38_N5
dffeas \register[10][8] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\register~87_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~45_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\register[10][8]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \register[10][8] .is_wysiwyg = "true";
defparam \register[10][8] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X67_Y38_N4
cycloneive_lcell_comb \Mux55~10 (
// Equation(s):
// \Mux55~10_combout  = (Selector91 & (((\register[10][8]~q ) # (Selector10)))) # (!Selector91 & (\register[8][8]~q  & ((!Selector10))))

	.dataa(\register[8][8]~q ),
	.datab(Selector91),
	.datac(\register[10][8]~q ),
	.datad(Selector10),
	.cin(gnd),
	.combout(\Mux55~10_combout ),
	.cout());
// synopsys translate_off
defparam \Mux55~10 .lut_mask = 16'hCCE2;
defparam \Mux55~10 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X66_Y38_N3
dffeas \register[11][8] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\register~87_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~47_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\register[11][8]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \register[11][8] .is_wysiwyg = "true";
defparam \register[11][8] .power_up = "low";
// synopsys translate_on

// Location: FF_X66_Y38_N5
dffeas \register[9][8] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\register~87_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~44_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\register[9][8]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \register[9][8] .is_wysiwyg = "true";
defparam \register[9][8] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X66_Y38_N4
cycloneive_lcell_comb \Mux55~11 (
// Equation(s):
// \Mux55~11_combout  = (\Mux55~10_combout  & ((\register[11][8]~q ) # ((!Selector10)))) # (!\Mux55~10_combout  & (((\register[9][8]~q  & Selector10))))

	.dataa(\Mux55~10_combout ),
	.datab(\register[11][8]~q ),
	.datac(\register[9][8]~q ),
	.datad(Selector10),
	.cin(gnd),
	.combout(\Mux55~11_combout ),
	.cout());
// synopsys translate_off
defparam \Mux55~11 .lut_mask = 16'hD8AA;
defparam \Mux55~11 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X67_Y33_N17
dffeas \register[6][8] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\register~87_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~58_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\register[6][8]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \register[6][8] .is_wysiwyg = "true";
defparam \register[6][8] .power_up = "low";
// synopsys translate_on

// Location: FF_X67_Y31_N1
dffeas \register[5][8] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\register~87_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~59_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\register[5][8]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \register[5][8] .is_wysiwyg = "true";
defparam \register[5][8] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X67_Y31_N0
cycloneive_lcell_comb \Mux55~12 (
// Equation(s):
// \Mux55~12_combout  = (Selector91 & (((Selector10)))) # (!Selector91 & ((Selector10 & ((\register[5][8]~q ))) # (!Selector10 & (\register[4][8]~q ))))

	.dataa(\register[4][8]~q ),
	.datab(Selector91),
	.datac(\register[5][8]~q ),
	.datad(Selector10),
	.cin(gnd),
	.combout(\Mux55~12_combout ),
	.cout());
// synopsys translate_off
defparam \Mux55~12 .lut_mask = 16'hFC22;
defparam \Mux55~12 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X67_Y33_N16
cycloneive_lcell_comb \Mux55~13 (
// Equation(s):
// \Mux55~13_combout  = (Selector91 & ((\Mux55~12_combout  & (\register[7][8]~q )) # (!\Mux55~12_combout  & ((\register[6][8]~q ))))) # (!Selector91 & (((\Mux55~12_combout ))))

	.dataa(\register[7][8]~q ),
	.datab(Selector91),
	.datac(\register[6][8]~q ),
	.datad(\Mux55~12_combout ),
	.cin(gnd),
	.combout(\Mux55~13_combout ),
	.cout());
// synopsys translate_off
defparam \Mux55~13 .lut_mask = 16'hBBC0;
defparam \Mux55~13 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X68_Y33_N27
dffeas \register[2][8] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\register~87_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~50_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\register[2][8]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \register[2][8] .is_wysiwyg = "true";
defparam \register[2][8] .power_up = "low";
// synopsys translate_on

// Location: FF_X70_Y34_N25
dffeas \register[3][8] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\register~87_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~48_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\register[3][8]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \register[3][8] .is_wysiwyg = "true";
defparam \register[3][8] .power_up = "low";
// synopsys translate_on

// Location: FF_X70_Y34_N11
dffeas \register[1][8] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\register~87_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~49_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\register[1][8]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \register[1][8] .is_wysiwyg = "true";
defparam \register[1][8] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X70_Y34_N24
cycloneive_lcell_comb \Mux55~14 (
// Equation(s):
// \Mux55~14_combout  = (Selector10 & ((Selector91 & (\register[3][8]~q )) # (!Selector91 & ((\register[1][8]~q )))))

	.dataa(Selector10),
	.datab(Selector91),
	.datac(\register[3][8]~q ),
	.datad(\register[1][8]~q ),
	.cin(gnd),
	.combout(\Mux55~14_combout ),
	.cout());
// synopsys translate_off
defparam \Mux55~14 .lut_mask = 16'hA280;
defparam \Mux55~14 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X68_Y33_N26
cycloneive_lcell_comb \Mux55~15 (
// Equation(s):
// \Mux55~15_combout  = (\Mux55~14_combout ) # ((!Selector10 & (Selector91 & \register[2][8]~q )))

	.dataa(Selector10),
	.datab(Selector91),
	.datac(\register[2][8]~q ),
	.datad(\Mux55~14_combout ),
	.cin(gnd),
	.combout(\Mux55~15_combout ),
	.cout());
// synopsys translate_off
defparam \Mux55~15 .lut_mask = 16'hFF40;
defparam \Mux55~15 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X67_Y33_N18
cycloneive_lcell_comb \Mux55~16 (
// Equation(s):
// \Mux55~16_combout  = (Selector8 & ((\Mux55~13_combout ) # ((Selector7)))) # (!Selector8 & (((!Selector7 & \Mux55~15_combout ))))

	.dataa(Selector8),
	.datab(\Mux55~13_combout ),
	.datac(Selector7),
	.datad(\Mux55~15_combout ),
	.cin(gnd),
	.combout(\Mux55~16_combout ),
	.cout());
// synopsys translate_off
defparam \Mux55~16 .lut_mask = 16'hADA8;
defparam \Mux55~16 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y36_N6
cycloneive_lcell_comb \register~88 (
// Equation(s):
// \register~88_combout  = (WideOr01 & ((\wdat[7]~48_combout ) # ((plif_memwbregsrc_l_1 & plif_memwbrtnaddr_l_7))))

	.dataa(plif_memwbregsrc_l_1),
	.datab(WideOr0),
	.datac(plif_memwbrtnaddr_l_7),
	.datad(wdat_7),
	.cin(gnd),
	.combout(\register~88_combout ),
	.cout());
// synopsys translate_off
defparam \register~88 .lut_mask = 16'hCC80;
defparam \register~88 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X62_Y31_N13
dffeas \register[23][7] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\register~88_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~37_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\register[23][7]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \register[23][7] .is_wysiwyg = "true";
defparam \register[23][7] .power_up = "low";
// synopsys translate_on

// Location: FF_X62_Y35_N9
dffeas \register[31][7] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\register~88_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~40_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\register[31][7]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \register[31][7] .is_wysiwyg = "true";
defparam \register[31][7] .power_up = "low";
// synopsys translate_on

// Location: FF_X62_Y31_N19
dffeas \register[19][7] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\register~88_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~39_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\register[19][7]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \register[19][7] .is_wysiwyg = "true";
defparam \register[19][7] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X61_Y31_N28
cycloneive_lcell_comb \register[27][7]~feeder (
// Equation(s):
// \register[27][7]~feeder_combout  = \register~88_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(\register~88_combout ),
	.cin(gnd),
	.combout(\register[27][7]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \register[27][7]~feeder .lut_mask = 16'hFF00;
defparam \register[27][7]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X61_Y31_N29
dffeas \register[27][7] (
	.clk(!CLK),
	.d(\register[27][7]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~38_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\register[27][7]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \register[27][7] .is_wysiwyg = "true";
defparam \register[27][7] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X62_Y31_N18
cycloneive_lcell_comb \Mux56~7 (
// Equation(s):
// \Mux56~7_combout  = (Selector8 & (Selector7)) # (!Selector8 & ((Selector7 & ((\register[27][7]~q ))) # (!Selector7 & (\register[19][7]~q ))))

	.dataa(Selector8),
	.datab(Selector7),
	.datac(\register[19][7]~q ),
	.datad(\register[27][7]~q ),
	.cin(gnd),
	.combout(\Mux56~7_combout ),
	.cout());
// synopsys translate_off
defparam \Mux56~7 .lut_mask = 16'hDC98;
defparam \Mux56~7 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y35_N8
cycloneive_lcell_comb \Mux56~8 (
// Equation(s):
// \Mux56~8_combout  = (Selector8 & ((\Mux56~7_combout  & ((\register[31][7]~q ))) # (!\Mux56~7_combout  & (\register[23][7]~q )))) # (!Selector8 & (((\Mux56~7_combout ))))

	.dataa(Selector8),
	.datab(\register[23][7]~q ),
	.datac(\register[31][7]~q ),
	.datad(\Mux56~7_combout ),
	.cin(gnd),
	.combout(\Mux56~8_combout ),
	.cout());
// synopsys translate_off
defparam \Mux56~8 .lut_mask = 16'hF588;
defparam \Mux56~8 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X63_Y33_N22
cycloneive_lcell_comb \register[29][7]~feeder (
// Equation(s):
// \register[29][7]~feeder_combout  = \register~88_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(\register~88_combout ),
	.datad(gnd),
	.cin(gnd),
	.combout(\register[29][7]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \register[29][7]~feeder .lut_mask = 16'hF0F0;
defparam \register[29][7]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X63_Y33_N23
dffeas \register[29][7] (
	.clk(!CLK),
	.d(\register[29][7]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~28_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\register[29][7]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \register[29][7] .is_wysiwyg = "true";
defparam \register[29][7] .power_up = "low";
// synopsys translate_on

// Location: FF_X63_Y35_N7
dffeas \register[21][7] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\register~88_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~22_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\register[21][7]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \register[21][7] .is_wysiwyg = "true";
defparam \register[21][7] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X62_Y36_N0
cycloneive_lcell_comb \register[25][7]~feeder (
// Equation(s):
// \register[25][7]~feeder_combout  = \register~88_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(\register~88_combout ),
	.cin(gnd),
	.combout(\register[25][7]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \register[25][7]~feeder .lut_mask = 16'hFF00;
defparam \register[25][7]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X62_Y36_N1
dffeas \register[25][7] (
	.clk(!CLK),
	.d(\register[25][7]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~24_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\register[25][7]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \register[25][7] .is_wysiwyg = "true";
defparam \register[25][7] .power_up = "low";
// synopsys translate_on

// Location: FF_X62_Y35_N11
dffeas \register[17][7] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\register~88_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~26_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\register[17][7]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \register[17][7] .is_wysiwyg = "true";
defparam \register[17][7] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X62_Y36_N14
cycloneive_lcell_comb \Mux56~0 (
// Equation(s):
// \Mux56~0_combout  = (Selector8 & (((Selector7)))) # (!Selector8 & ((Selector7 & (\register[25][7]~q )) # (!Selector7 & ((\register[17][7]~q )))))

	.dataa(Selector8),
	.datab(\register[25][7]~q ),
	.datac(\register[17][7]~q ),
	.datad(Selector7),
	.cin(gnd),
	.combout(\Mux56~0_combout ),
	.cout());
// synopsys translate_off
defparam \Mux56~0 .lut_mask = 16'hEE50;
defparam \Mux56~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X63_Y35_N6
cycloneive_lcell_comb \Mux56~1 (
// Equation(s):
// \Mux56~1_combout  = (Selector8 & ((\Mux56~0_combout  & (\register[29][7]~q )) # (!\Mux56~0_combout  & ((\register[21][7]~q ))))) # (!Selector8 & (((\Mux56~0_combout ))))

	.dataa(\register[29][7]~q ),
	.datab(Selector8),
	.datac(\register[21][7]~q ),
	.datad(\Mux56~0_combout ),
	.cin(gnd),
	.combout(\Mux56~1_combout ),
	.cout());
// synopsys translate_off
defparam \Mux56~1 .lut_mask = 16'hBBC0;
defparam \Mux56~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X70_Y38_N16
cycloneive_lcell_comb \register[24][7]~feeder (
// Equation(s):
// \register[24][7]~feeder_combout  = \register~88_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(\register~88_combout ),
	.cin(gnd),
	.combout(\register[24][7]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \register[24][7]~feeder .lut_mask = 16'hFF00;
defparam \register[24][7]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X70_Y38_N17
dffeas \register[24][7] (
	.clk(!CLK),
	.d(\register[24][7]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~34_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\register[24][7]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \register[24][7] .is_wysiwyg = "true";
defparam \register[24][7] .power_up = "low";
// synopsys translate_on

// Location: FF_X66_Y35_N3
dffeas \register[28][7] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\register~88_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~57_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\register[28][7]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \register[28][7] .is_wysiwyg = "true";
defparam \register[28][7] .power_up = "low";
// synopsys translate_on

// Location: FF_X69_Y38_N13
dffeas \register[16][7] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\register~88_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~36_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\register[16][7]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \register[16][7] .is_wysiwyg = "true";
defparam \register[16][7] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X69_Y38_N12
cycloneive_lcell_comb \Mux56~4 (
// Equation(s):
// \Mux56~4_combout  = (Selector8 & ((\register[20][7]~q ) # ((Selector7)))) # (!Selector8 & (((\register[16][7]~q  & !Selector7))))

	.dataa(\register[20][7]~q ),
	.datab(Selector8),
	.datac(\register[16][7]~q ),
	.datad(Selector7),
	.cin(gnd),
	.combout(\Mux56~4_combout ),
	.cout());
// synopsys translate_off
defparam \Mux56~4 .lut_mask = 16'hCCB8;
defparam \Mux56~4 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X66_Y35_N2
cycloneive_lcell_comb \Mux56~5 (
// Equation(s):
// \Mux56~5_combout  = (Selector7 & ((\Mux56~4_combout  & ((\register[28][7]~q ))) # (!\Mux56~4_combout  & (\register[24][7]~q )))) # (!Selector7 & (((\Mux56~4_combout ))))

	.dataa(Selector7),
	.datab(\register[24][7]~q ),
	.datac(\register[28][7]~q ),
	.datad(\Mux56~4_combout ),
	.cin(gnd),
	.combout(\Mux56~5_combout ),
	.cout());
// synopsys translate_off
defparam \Mux56~5 .lut_mask = 16'hF588;
defparam \Mux56~5 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X68_Y38_N19
dffeas \register[26][7] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\register~88_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~54_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\register[26][7]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \register[26][7] .is_wysiwyg = "true";
defparam \register[26][7] .power_up = "low";
// synopsys translate_on

// Location: FF_X66_Y35_N17
dffeas \register[30][7] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\register~88_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~56_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\register[30][7]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \register[30][7] .is_wysiwyg = "true";
defparam \register[30][7] .power_up = "low";
// synopsys translate_on

// Location: FF_X68_Y38_N29
dffeas \register[18][7] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\register~88_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~33_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\register[18][7]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \register[18][7] .is_wysiwyg = "true";
defparam \register[18][7] .power_up = "low";
// synopsys translate_on

// Location: FF_X67_Y37_N1
dffeas \register[22][7] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\register~88_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~55_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\register[22][7]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \register[22][7] .is_wysiwyg = "true";
defparam \register[22][7] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X68_Y38_N28
cycloneive_lcell_comb \Mux56~2 (
// Equation(s):
// \Mux56~2_combout  = (Selector7 & (Selector8)) # (!Selector7 & ((Selector8 & ((\register[22][7]~q ))) # (!Selector8 & (\register[18][7]~q ))))

	.dataa(Selector7),
	.datab(Selector8),
	.datac(\register[18][7]~q ),
	.datad(\register[22][7]~q ),
	.cin(gnd),
	.combout(\Mux56~2_combout ),
	.cout());
// synopsys translate_off
defparam \Mux56~2 .lut_mask = 16'hDC98;
defparam \Mux56~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X66_Y35_N16
cycloneive_lcell_comb \Mux56~3 (
// Equation(s):
// \Mux56~3_combout  = (Selector7 & ((\Mux56~2_combout  & ((\register[30][7]~q ))) # (!\Mux56~2_combout  & (\register[26][7]~q )))) # (!Selector7 & (((\Mux56~2_combout ))))

	.dataa(Selector7),
	.datab(\register[26][7]~q ),
	.datac(\register[30][7]~q ),
	.datad(\Mux56~2_combout ),
	.cin(gnd),
	.combout(\Mux56~3_combout ),
	.cout());
// synopsys translate_off
defparam \Mux56~3 .lut_mask = 16'hF588;
defparam \Mux56~3 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X66_Y35_N24
cycloneive_lcell_comb \Mux56~6 (
// Equation(s):
// \Mux56~6_combout  = (Selector91 & (((Selector10) # (\Mux56~3_combout )))) # (!Selector91 & (\Mux56~5_combout  & (!Selector10)))

	.dataa(Selector91),
	.datab(\Mux56~5_combout ),
	.datac(Selector10),
	.datad(\Mux56~3_combout ),
	.cin(gnd),
	.combout(\Mux56~6_combout ),
	.cout());
// synopsys translate_off
defparam \Mux56~6 .lut_mask = 16'hAEA4;
defparam \Mux56~6 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X66_Y38_N27
dffeas \register[11][7] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\register~88_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~47_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\register[11][7]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \register[11][7] .is_wysiwyg = "true";
defparam \register[11][7] .power_up = "low";
// synopsys translate_on

// Location: FF_X66_Y38_N17
dffeas \register[9][7] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\register~88_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~44_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\register[9][7]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \register[9][7] .is_wysiwyg = "true";
defparam \register[9][7] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X66_Y38_N26
cycloneive_lcell_comb \Mux56~13 (
// Equation(s):
// \Mux56~13_combout  = (\Mux56~12_combout  & (((\register[11][7]~q )) # (!Selector10))) # (!\Mux56~12_combout  & (Selector10 & ((\register[9][7]~q ))))

	.dataa(\Mux56~12_combout ),
	.datab(Selector10),
	.datac(\register[11][7]~q ),
	.datad(\register[9][7]~q ),
	.cin(gnd),
	.combout(\Mux56~13_combout ),
	.cout());
// synopsys translate_off
defparam \Mux56~13 .lut_mask = 16'hE6A2;
defparam \Mux56~13 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X68_Y33_N9
dffeas \register[2][7] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\register~88_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~50_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\register[2][7]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \register[2][7] .is_wysiwyg = "true";
defparam \register[2][7] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X70_Y33_N24
cycloneive_lcell_comb \register[3][7]~feeder (
// Equation(s):
// \register[3][7]~feeder_combout  = \register~88_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(\register~88_combout ),
	.cin(gnd),
	.combout(\register[3][7]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \register[3][7]~feeder .lut_mask = 16'hFF00;
defparam \register[3][7]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X70_Y33_N25
dffeas \register[3][7] (
	.clk(!CLK),
	.d(\register[3][7]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~48_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\register[3][7]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \register[3][7] .is_wysiwyg = "true";
defparam \register[3][7] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X70_Y33_N10
cycloneive_lcell_comb \register[1][7]~feeder (
// Equation(s):
// \register[1][7]~feeder_combout  = \register~88_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(\register~88_combout ),
	.cin(gnd),
	.combout(\register[1][7]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \register[1][7]~feeder .lut_mask = 16'hFF00;
defparam \register[1][7]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X70_Y33_N11
dffeas \register[1][7] (
	.clk(!CLK),
	.d(\register[1][7]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~49_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\register[1][7]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \register[1][7] .is_wysiwyg = "true";
defparam \register[1][7] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X70_Y33_N12
cycloneive_lcell_comb \Mux56~14 (
// Equation(s):
// \Mux56~14_combout  = (plif_ifidinstr_l_17 & ((Selector9 & (\register[3][7]~q )) # (!Selector9 & ((\register[1][7]~q ))))) # (!plif_ifidinstr_l_17 & (((\register[1][7]~q ))))

	.dataa(plif_ifidinstr_l_17),
	.datab(\register[3][7]~q ),
	.datac(Selector9),
	.datad(\register[1][7]~q ),
	.cin(gnd),
	.combout(\Mux56~14_combout ),
	.cout());
// synopsys translate_off
defparam \Mux56~14 .lut_mask = 16'hDF80;
defparam \Mux56~14 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X68_Y33_N8
cycloneive_lcell_comb \Mux56~15 (
// Equation(s):
// \Mux56~15_combout  = (Selector10 & (((\Mux56~14_combout )))) # (!Selector10 & (Selector91 & (\register[2][7]~q )))

	.dataa(Selector10),
	.datab(Selector91),
	.datac(\register[2][7]~q ),
	.datad(\Mux56~14_combout ),
	.cin(gnd),
	.combout(\Mux56~15_combout ),
	.cout());
// synopsys translate_off
defparam \Mux56~15 .lut_mask = 16'hEA40;
defparam \Mux56~15 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X67_Y39_N14
cycloneive_lcell_comb \Mux56~16 (
// Equation(s):
// \Mux56~16_combout  = (Selector7 & ((\Mux56~13_combout ) # ((Selector8)))) # (!Selector7 & (((!Selector8 & \Mux56~15_combout ))))

	.dataa(Selector7),
	.datab(\Mux56~13_combout ),
	.datac(Selector8),
	.datad(\Mux56~15_combout ),
	.cin(gnd),
	.combout(\Mux56~16_combout ),
	.cout());
// synopsys translate_off
defparam \Mux56~16 .lut_mask = 16'hADA8;
defparam \Mux56~16 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X68_Y32_N11
dffeas \register[7][7] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\register~88_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~43_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\register[7][7]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \register[7][7] .is_wysiwyg = "true";
defparam \register[7][7] .power_up = "low";
// synopsys translate_on

// Location: FF_X68_Y32_N5
dffeas \register[6][7] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\register~88_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~58_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\register[6][7]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \register[6][7] .is_wysiwyg = "true";
defparam \register[6][7] .power_up = "low";
// synopsys translate_on

// Location: FF_X67_Y31_N15
dffeas \register[4][7] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\register~88_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~60_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\register[4][7]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \register[4][7] .is_wysiwyg = "true";
defparam \register[4][7] .power_up = "low";
// synopsys translate_on

// Location: FF_X67_Y31_N25
dffeas \register[5][7] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\register~88_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~59_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\register[5][7]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \register[5][7] .is_wysiwyg = "true";
defparam \register[5][7] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X67_Y31_N24
cycloneive_lcell_comb \Mux56~10 (
// Equation(s):
// \Mux56~10_combout  = (Selector10 & (((\register[5][7]~q ) # (Selector91)))) # (!Selector10 & (\register[4][7]~q  & ((!Selector91))))

	.dataa(Selector10),
	.datab(\register[4][7]~q ),
	.datac(\register[5][7]~q ),
	.datad(Selector91),
	.cin(gnd),
	.combout(\Mux56~10_combout ),
	.cout());
// synopsys translate_off
defparam \Mux56~10 .lut_mask = 16'hAAE4;
defparam \Mux56~10 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X68_Y32_N4
cycloneive_lcell_comb \Mux56~11 (
// Equation(s):
// \Mux56~11_combout  = (Selector91 & ((\Mux56~10_combout  & (\register[7][7]~q )) # (!\Mux56~10_combout  & ((\register[6][7]~q ))))) # (!Selector91 & (((\Mux56~10_combout ))))

	.dataa(\register[7][7]~q ),
	.datab(Selector91),
	.datac(\register[6][7]~q ),
	.datad(\Mux56~10_combout ),
	.cin(gnd),
	.combout(\Mux56~11_combout ),
	.cout());
// synopsys translate_off
defparam \Mux56~11 .lut_mask = 16'hBBC0;
defparam \Mux56~11 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y36_N28
cycloneive_lcell_comb \register[15][7]~feeder (
// Equation(s):
// \register[15][7]~feeder_combout  = \register~88_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(\register~88_combout ),
	.cin(gnd),
	.combout(\register[15][7]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \register[15][7]~feeder .lut_mask = 16'hFF00;
defparam \register[15][7]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X62_Y36_N29
dffeas \register[15][7] (
	.clk(!CLK),
	.d(\register[15][7]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~53_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\register[15][7]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \register[15][7] .is_wysiwyg = "true";
defparam \register[15][7] .power_up = "low";
// synopsys translate_on

// Location: FF_X67_Y33_N7
dffeas \register[14][7] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\register~88_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~61_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\register[14][7]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \register[14][7] .is_wysiwyg = "true";
defparam \register[14][7] .power_up = "low";
// synopsys translate_on

// Location: FF_X63_Y30_N25
dffeas \register[13][7] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\register~88_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~62_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\register[13][7]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \register[13][7] .is_wysiwyg = "true";
defparam \register[13][7] .power_up = "low";
// synopsys translate_on

// Location: FF_X63_Y30_N7
dffeas \register[12][7] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\register~88_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~52_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\register[12][7]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \register[12][7] .is_wysiwyg = "true";
defparam \register[12][7] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X63_Y30_N24
cycloneive_lcell_comb \Mux56~17 (
// Equation(s):
// \Mux56~17_combout  = (Selector91 & (Selector10)) # (!Selector91 & ((Selector10 & (\register[13][7]~q )) # (!Selector10 & ((\register[12][7]~q )))))

	.dataa(Selector91),
	.datab(Selector10),
	.datac(\register[13][7]~q ),
	.datad(\register[12][7]~q ),
	.cin(gnd),
	.combout(\Mux56~17_combout ),
	.cout());
// synopsys translate_off
defparam \Mux56~17 .lut_mask = 16'hD9C8;
defparam \Mux56~17 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X67_Y33_N6
cycloneive_lcell_comb \Mux56~18 (
// Equation(s):
// \Mux56~18_combout  = (Selector91 & ((\Mux56~17_combout  & (\register[15][7]~q )) # (!\Mux56~17_combout  & ((\register[14][7]~q ))))) # (!Selector91 & (((\Mux56~17_combout ))))

	.dataa(\register[15][7]~q ),
	.datab(Selector91),
	.datac(\register[14][7]~q ),
	.datad(\Mux56~17_combout ),
	.cin(gnd),
	.combout(\Mux56~18_combout ),
	.cout());
// synopsys translate_off
defparam \Mux56~18 .lut_mask = 16'hBBC0;
defparam \Mux56~18 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X63_Y37_N8
cycloneive_lcell_comb \register~89 (
// Equation(s):
// \register~89_combout  = (WideOr01 & ((\wdat[6]~50_combout ) # ((plif_memwbregsrc_l_1 & plif_memwbrtnaddr_l_6))))

	.dataa(plif_memwbregsrc_l_1),
	.datab(plif_memwbrtnaddr_l_6),
	.datac(WideOr0),
	.datad(wdat_6),
	.cin(gnd),
	.combout(\register~89_combout ),
	.cout());
// synopsys translate_off
defparam \register~89 .lut_mask = 16'hF080;
defparam \register~89 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X62_Y38_N5
dffeas \register[23][6] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\register~89_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~37_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\register[23][6]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \register[23][6] .is_wysiwyg = "true";
defparam \register[23][6] .power_up = "low";
// synopsys translate_on

// Location: FF_X62_Y38_N15
dffeas \register[19][6] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\register~89_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~39_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\register[19][6]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \register[19][6] .is_wysiwyg = "true";
defparam \register[19][6] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X62_Y38_N14
cycloneive_lcell_comb \Mux57~7 (
// Equation(s):
// \Mux57~7_combout  = (Selector7 & (((Selector8)))) # (!Selector7 & ((Selector8 & (\register[23][6]~q )) # (!Selector8 & ((\register[19][6]~q )))))

	.dataa(Selector7),
	.datab(\register[23][6]~q ),
	.datac(\register[19][6]~q ),
	.datad(Selector8),
	.cin(gnd),
	.combout(\Mux57~7_combout ),
	.cout());
// synopsys translate_off
defparam \Mux57~7 .lut_mask = 16'hEE50;
defparam \Mux57~7 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X65_Y30_N18
cycloneive_lcell_comb \register[31][6]~feeder (
// Equation(s):
// \register[31][6]~feeder_combout  = \register~89_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(\register~89_combout ),
	.cin(gnd),
	.combout(\register[31][6]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \register[31][6]~feeder .lut_mask = 16'hFF00;
defparam \register[31][6]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X65_Y30_N19
dffeas \register[31][6] (
	.clk(!CLK),
	.d(\register[31][6]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~40_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\register[31][6]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \register[31][6] .is_wysiwyg = "true";
defparam \register[31][6] .power_up = "low";
// synopsys translate_on

// Location: FF_X62_Y39_N27
dffeas \register[27][6] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\register~89_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~38_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\register[27][6]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \register[27][6] .is_wysiwyg = "true";
defparam \register[27][6] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X65_Y30_N8
cycloneive_lcell_comb \Mux57~8 (
// Equation(s):
// \Mux57~8_combout  = (Selector7 & ((\Mux57~7_combout  & (\register[31][6]~q )) # (!\Mux57~7_combout  & ((\register[27][6]~q ))))) # (!Selector7 & (\Mux57~7_combout ))

	.dataa(Selector7),
	.datab(\Mux57~7_combout ),
	.datac(\register[31][6]~q ),
	.datad(\register[27][6]~q ),
	.cin(gnd),
	.combout(\Mux57~8_combout ),
	.cout());
// synopsys translate_off
defparam \Mux57~8 .lut_mask = 16'hE6C4;
defparam \Mux57~8 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X69_Y37_N31
dffeas \register[22][6] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\register~89_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~55_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\register[22][6]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \register[22][6] .is_wysiwyg = "true";
defparam \register[22][6] .power_up = "low";
// synopsys translate_on

// Location: FF_X68_Y37_N1
dffeas \register[30][6] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\register~89_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~56_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\register[30][6]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \register[30][6] .is_wysiwyg = "true";
defparam \register[30][6] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X68_Y37_N0
cycloneive_lcell_comb \Mux57~3 (
// Equation(s):
// \Mux57~3_combout  = (\Mux57~2_combout  & (((\register[30][6]~q ) # (!Selector8)))) # (!\Mux57~2_combout  & (\register[22][6]~q  & ((Selector8))))

	.dataa(\Mux57~2_combout ),
	.datab(\register[22][6]~q ),
	.datac(\register[30][6]~q ),
	.datad(Selector8),
	.cin(gnd),
	.combout(\Mux57~3_combout ),
	.cout());
// synopsys translate_off
defparam \Mux57~3 .lut_mask = 16'hE4AA;
defparam \Mux57~3 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X65_Y37_N27
dffeas \register[20][6] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\register~89_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~35_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\register[20][6]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \register[20][6] .is_wysiwyg = "true";
defparam \register[20][6] .power_up = "low";
// synopsys translate_on

// Location: FF_X65_Y38_N15
dffeas \register[28][6] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\register~89_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~57_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\register[28][6]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \register[28][6] .is_wysiwyg = "true";
defparam \register[28][6] .power_up = "low";
// synopsys translate_on

// Location: FF_X65_Y38_N1
dffeas \register[24][6] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\register~89_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~34_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\register[24][6]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \register[24][6] .is_wysiwyg = "true";
defparam \register[24][6] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X65_Y38_N0
cycloneive_lcell_comb \Mux57~4 (
// Equation(s):
// \Mux57~4_combout  = (Selector8 & (((Selector7)))) # (!Selector8 & ((Selector7 & ((\register[24][6]~q ))) # (!Selector7 & (\register[16][6]~q ))))

	.dataa(\register[16][6]~q ),
	.datab(Selector8),
	.datac(\register[24][6]~q ),
	.datad(Selector7),
	.cin(gnd),
	.combout(\Mux57~4_combout ),
	.cout());
// synopsys translate_off
defparam \Mux57~4 .lut_mask = 16'hFC22;
defparam \Mux57~4 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X65_Y38_N14
cycloneive_lcell_comb \Mux57~5 (
// Equation(s):
// \Mux57~5_combout  = (Selector8 & ((\Mux57~4_combout  & ((\register[28][6]~q ))) # (!\Mux57~4_combout  & (\register[20][6]~q )))) # (!Selector8 & (((\Mux57~4_combout ))))

	.dataa(Selector8),
	.datab(\register[20][6]~q ),
	.datac(\register[28][6]~q ),
	.datad(\Mux57~4_combout ),
	.cin(gnd),
	.combout(\Mux57~5_combout ),
	.cout());
// synopsys translate_off
defparam \Mux57~5 .lut_mask = 16'hF588;
defparam \Mux57~5 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X65_Y30_N4
cycloneive_lcell_comb \Mux57~6 (
// Equation(s):
// \Mux57~6_combout  = (Selector10 & (((Selector91)))) # (!Selector10 & ((Selector91 & (\Mux57~3_combout )) # (!Selector91 & ((\Mux57~5_combout )))))

	.dataa(\Mux57~3_combout ),
	.datab(Selector10),
	.datac(\Mux57~5_combout ),
	.datad(Selector91),
	.cin(gnd),
	.combout(\Mux57~6_combout ),
	.cout());
// synopsys translate_off
defparam \Mux57~6 .lut_mask = 16'hEE30;
defparam \Mux57~6 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X63_Y33_N26
cycloneive_lcell_comb \register[29][6]~feeder (
// Equation(s):
// \register[29][6]~feeder_combout  = \register~89_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(\register~89_combout ),
	.datad(gnd),
	.cin(gnd),
	.combout(\register[29][6]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \register[29][6]~feeder .lut_mask = 16'hF0F0;
defparam \register[29][6]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X63_Y33_N27
dffeas \register[29][6] (
	.clk(!CLK),
	.d(\register[29][6]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~28_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\register[29][6]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \register[29][6] .is_wysiwyg = "true";
defparam \register[29][6] .power_up = "low";
// synopsys translate_on

// Location: FF_X63_Y33_N25
dffeas \register[21][6] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\register~89_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~22_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\register[21][6]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \register[21][6] .is_wysiwyg = "true";
defparam \register[21][6] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X63_Y33_N24
cycloneive_lcell_comb \Mux57~0 (
// Equation(s):
// \Mux57~0_combout  = (Selector8 & (((\register[21][6]~q ) # (Selector7)))) # (!Selector8 & (\register[17][6]~q  & ((!Selector7))))

	.dataa(\register[17][6]~q ),
	.datab(Selector8),
	.datac(\register[21][6]~q ),
	.datad(Selector7),
	.cin(gnd),
	.combout(\Mux57~0_combout ),
	.cout());
// synopsys translate_off
defparam \Mux57~0 .lut_mask = 16'hCCE2;
defparam \Mux57~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X63_Y31_N0
cycloneive_lcell_comb \register[25][6]~feeder (
// Equation(s):
// \register[25][6]~feeder_combout  = \register~89_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(\register~89_combout ),
	.datad(gnd),
	.cin(gnd),
	.combout(\register[25][6]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \register[25][6]~feeder .lut_mask = 16'hF0F0;
defparam \register[25][6]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X63_Y31_N1
dffeas \register[25][6] (
	.clk(!CLK),
	.d(\register[25][6]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~24_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\register[25][6]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \register[25][6] .is_wysiwyg = "true";
defparam \register[25][6] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X63_Y31_N30
cycloneive_lcell_comb \Mux57~1 (
// Equation(s):
// \Mux57~1_combout  = (Selector7 & ((\Mux57~0_combout  & (\register[29][6]~q )) # (!\Mux57~0_combout  & ((\register[25][6]~q ))))) # (!Selector7 & (((\Mux57~0_combout ))))

	.dataa(\register[29][6]~q ),
	.datab(Selector7),
	.datac(\Mux57~0_combout ),
	.datad(\register[25][6]~q ),
	.cin(gnd),
	.combout(\Mux57~1_combout ),
	.cout());
// synopsys translate_off
defparam \Mux57~1 .lut_mask = 16'hBCB0;
defparam \Mux57~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X66_Y34_N25
dffeas \register[11][6] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\register~89_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~47_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\register[11][6]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \register[11][6] .is_wysiwyg = "true";
defparam \register[11][6] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X63_Y34_N2
cycloneive_lcell_comb \register[9][6]~feeder (
// Equation(s):
// \register[9][6]~feeder_combout  = \register~89_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(\register~89_combout ),
	.datad(gnd),
	.cin(gnd),
	.combout(\register[9][6]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \register[9][6]~feeder .lut_mask = 16'hF0F0;
defparam \register[9][6]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X63_Y34_N3
dffeas \register[9][6] (
	.clk(!CLK),
	.d(\register[9][6]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~44_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\register[9][6]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \register[9][6] .is_wysiwyg = "true";
defparam \register[9][6] .power_up = "low";
// synopsys translate_on

// Location: FF_X67_Y38_N19
dffeas \register[8][6] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\register~89_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~46_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\register[8][6]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \register[8][6] .is_wysiwyg = "true";
defparam \register[8][6] .power_up = "low";
// synopsys translate_on

// Location: FF_X67_Y38_N1
dffeas \register[10][6] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\register~89_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~45_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\register[10][6]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \register[10][6] .is_wysiwyg = "true";
defparam \register[10][6] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X67_Y38_N0
cycloneive_lcell_comb \Mux57~10 (
// Equation(s):
// \Mux57~10_combout  = (Selector10 & (((Selector91)))) # (!Selector10 & ((Selector91 & ((\register[10][6]~q ))) # (!Selector91 & (\register[8][6]~q ))))

	.dataa(Selector10),
	.datab(\register[8][6]~q ),
	.datac(\register[10][6]~q ),
	.datad(Selector91),
	.cin(gnd),
	.combout(\Mux57~10_combout ),
	.cout());
// synopsys translate_off
defparam \Mux57~10 .lut_mask = 16'hFA44;
defparam \Mux57~10 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X63_Y34_N16
cycloneive_lcell_comb \Mux57~11 (
// Equation(s):
// \Mux57~11_combout  = (Selector10 & ((\Mux57~10_combout  & (\register[11][6]~q )) # (!\Mux57~10_combout  & ((\register[9][6]~q ))))) # (!Selector10 & (((\Mux57~10_combout ))))

	.dataa(\register[11][6]~q ),
	.datab(\register[9][6]~q ),
	.datac(Selector10),
	.datad(\Mux57~10_combout ),
	.cin(gnd),
	.combout(\Mux57~11_combout ),
	.cout());
// synopsys translate_off
defparam \Mux57~11 .lut_mask = 16'hAFC0;
defparam \Mux57~11 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X66_Y34_N23
dffeas \register[2][6] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\register~89_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~50_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\register[2][6]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \register[2][6] .is_wysiwyg = "true";
defparam \register[2][6] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X70_Y33_N28
cycloneive_lcell_comb \register[1][6]~feeder (
// Equation(s):
// \register[1][6]~feeder_combout  = \register~89_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(\register~89_combout ),
	.cin(gnd),
	.combout(\register[1][6]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \register[1][6]~feeder .lut_mask = 16'hFF00;
defparam \register[1][6]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X70_Y33_N29
dffeas \register[1][6] (
	.clk(!CLK),
	.d(\register[1][6]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~49_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\register[1][6]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \register[1][6] .is_wysiwyg = "true";
defparam \register[1][6] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X70_Y33_N18
cycloneive_lcell_comb \register[3][6]~feeder (
// Equation(s):
// \register[3][6]~feeder_combout  = \register~89_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(\register~89_combout ),
	.cin(gnd),
	.combout(\register[3][6]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \register[3][6]~feeder .lut_mask = 16'hFF00;
defparam \register[3][6]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X70_Y33_N19
dffeas \register[3][6] (
	.clk(!CLK),
	.d(\register[3][6]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~48_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\register[3][6]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \register[3][6] .is_wysiwyg = "true";
defparam \register[3][6] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X70_Y33_N26
cycloneive_lcell_comb \Mux57~14 (
// Equation(s):
// \Mux57~14_combout  = (plif_ifidinstr_l_17 & ((Selector9 & ((\register[3][6]~q ))) # (!Selector9 & (\register[1][6]~q )))) # (!plif_ifidinstr_l_17 & (\register[1][6]~q ))

	.dataa(plif_ifidinstr_l_17),
	.datab(\register[1][6]~q ),
	.datac(Selector9),
	.datad(\register[3][6]~q ),
	.cin(gnd),
	.combout(\Mux57~14_combout ),
	.cout());
// synopsys translate_off
defparam \Mux57~14 .lut_mask = 16'hEC4C;
defparam \Mux57~14 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X65_Y30_N24
cycloneive_lcell_comb \Mux57~15 (
// Equation(s):
// \Mux57~15_combout  = (Selector10 & (((\Mux57~14_combout )))) # (!Selector10 & (Selector91 & (\register[2][6]~q )))

	.dataa(Selector10),
	.datab(Selector91),
	.datac(\register[2][6]~q ),
	.datad(\Mux57~14_combout ),
	.cin(gnd),
	.combout(\Mux57~15_combout ),
	.cout());
// synopsys translate_off
defparam \Mux57~15 .lut_mask = 16'hEA40;
defparam \Mux57~15 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X66_Y32_N11
dffeas \register[7][6] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\register~89_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~43_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\register[7][6]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \register[7][6] .is_wysiwyg = "true";
defparam \register[7][6] .power_up = "low";
// synopsys translate_on

// Location: FF_X67_Y31_N11
dffeas \register[4][6] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\register~89_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~60_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\register[4][6]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \register[4][6] .is_wysiwyg = "true";
defparam \register[4][6] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X67_Y31_N10
cycloneive_lcell_comb \Mux57~12 (
// Equation(s):
// \Mux57~12_combout  = (Selector91 & (((Selector10)))) # (!Selector91 & ((Selector10 & (\register[5][6]~q )) # (!Selector10 & ((\register[4][6]~q )))))

	.dataa(\register[5][6]~q ),
	.datab(Selector91),
	.datac(\register[4][6]~q ),
	.datad(Selector10),
	.cin(gnd),
	.combout(\Mux57~12_combout ),
	.cout());
// synopsys translate_off
defparam \Mux57~12 .lut_mask = 16'hEE30;
defparam \Mux57~12 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X66_Y32_N10
cycloneive_lcell_comb \Mux57~13 (
// Equation(s):
// \Mux57~13_combout  = (Selector91 & ((\Mux57~12_combout  & ((\register[7][6]~q ))) # (!\Mux57~12_combout  & (\register[6][6]~q )))) # (!Selector91 & (((\Mux57~12_combout ))))

	.dataa(\register[6][6]~q ),
	.datab(Selector91),
	.datac(\register[7][6]~q ),
	.datad(\Mux57~12_combout ),
	.cin(gnd),
	.combout(\Mux57~13_combout ),
	.cout());
// synopsys translate_off
defparam \Mux57~13 .lut_mask = 16'hF388;
defparam \Mux57~13 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X65_Y30_N26
cycloneive_lcell_comb \Mux57~16 (
// Equation(s):
// \Mux57~16_combout  = (Selector7 & (((Selector8)))) # (!Selector7 & ((Selector8 & ((\Mux57~13_combout ))) # (!Selector8 & (\Mux57~15_combout ))))

	.dataa(Selector7),
	.datab(\Mux57~15_combout ),
	.datac(Selector8),
	.datad(\Mux57~13_combout ),
	.cin(gnd),
	.combout(\Mux57~16_combout ),
	.cout());
// synopsys translate_off
defparam \Mux57~16 .lut_mask = 16'hF4A4;
defparam \Mux57~16 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X63_Y37_N9
dffeas \register[15][6] (
	.clk(!CLK),
	.d(\register~89_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~53_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\register[15][6]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \register[15][6] .is_wysiwyg = "true";
defparam \register[15][6] .power_up = "low";
// synopsys translate_on

// Location: FF_X63_Y30_N19
dffeas \register[12][6] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\register~89_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~52_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\register[12][6]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \register[12][6] .is_wysiwyg = "true";
defparam \register[12][6] .power_up = "low";
// synopsys translate_on

// Location: FF_X63_Y30_N9
dffeas \register[13][6] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\register~89_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~62_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\register[13][6]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \register[13][6] .is_wysiwyg = "true";
defparam \register[13][6] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X63_Y30_N8
cycloneive_lcell_comb \Mux57~17 (
// Equation(s):
// \Mux57~17_combout  = (Selector91 & (((Selector10)))) # (!Selector91 & ((Selector10 & ((\register[13][6]~q ))) # (!Selector10 & (\register[12][6]~q ))))

	.dataa(Selector91),
	.datab(\register[12][6]~q ),
	.datac(\register[13][6]~q ),
	.datad(Selector10),
	.cin(gnd),
	.combout(\Mux57~17_combout ),
	.cout());
// synopsys translate_off
defparam \Mux57~17 .lut_mask = 16'hFA44;
defparam \Mux57~17 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X67_Y33_N4
cycloneive_lcell_comb \register[14][6]~feeder (
// Equation(s):
// \register[14][6]~feeder_combout  = \register~89_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(\register~89_combout ),
	.datad(gnd),
	.cin(gnd),
	.combout(\register[14][6]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \register[14][6]~feeder .lut_mask = 16'hF0F0;
defparam \register[14][6]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X67_Y33_N5
dffeas \register[14][6] (
	.clk(!CLK),
	.d(\register[14][6]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~61_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\register[14][6]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \register[14][6] .is_wysiwyg = "true";
defparam \register[14][6] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X65_Y30_N12
cycloneive_lcell_comb \Mux57~18 (
// Equation(s):
// \Mux57~18_combout  = (Selector91 & ((\Mux57~17_combout  & (\register[15][6]~q )) # (!\Mux57~17_combout  & ((\register[14][6]~q ))))) # (!Selector91 & (((\Mux57~17_combout ))))

	.dataa(\register[15][6]~q ),
	.datab(Selector91),
	.datac(\Mux57~17_combout ),
	.datad(\register[14][6]~q ),
	.cin(gnd),
	.combout(\Mux57~18_combout ),
	.cout());
// synopsys translate_off
defparam \Mux57~18 .lut_mask = 16'hBCB0;
defparam \Mux57~18 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X63_Y37_N14
cycloneive_lcell_comb \register~90 (
// Equation(s):
// \register~90_combout  = (WideOr01 & ((\wdat[5]~52_combout ) # ((plif_memwbrtnaddr_l_5 & plif_memwbregsrc_l_1))))

	.dataa(WideOr0),
	.datab(plif_memwbrtnaddr_l_5),
	.datac(wdat_5),
	.datad(plif_memwbregsrc_l_1),
	.cin(gnd),
	.combout(\register~90_combout ),
	.cout());
// synopsys translate_off
defparam \register~90 .lut_mask = 16'hA8A0;
defparam \register~90 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X62_Y31_N9
dffeas \register[23][5] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\register~90_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~37_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\register[23][5]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \register[23][5] .is_wysiwyg = "true";
defparam \register[23][5] .power_up = "low";
// synopsys translate_on

// Location: FF_X65_Y30_N3
dffeas \register[31][5] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\register~90_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~40_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\register[31][5]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \register[31][5] .is_wysiwyg = "true";
defparam \register[31][5] .power_up = "low";
// synopsys translate_on

// Location: FF_X62_Y31_N11
dffeas \register[19][5] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\register~90_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~39_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\register[19][5]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \register[19][5] .is_wysiwyg = "true";
defparam \register[19][5] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X63_Y31_N24
cycloneive_lcell_comb \register[27][5]~feeder (
// Equation(s):
// \register[27][5]~feeder_combout  = \register~90_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(\register~90_combout ),
	.cin(gnd),
	.combout(\register[27][5]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \register[27][5]~feeder .lut_mask = 16'hFF00;
defparam \register[27][5]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X63_Y31_N25
dffeas \register[27][5] (
	.clk(!CLK),
	.d(\register[27][5]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~38_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\register[27][5]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \register[27][5] .is_wysiwyg = "true";
defparam \register[27][5] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X62_Y31_N10
cycloneive_lcell_comb \Mux58~7 (
// Equation(s):
// \Mux58~7_combout  = (Selector8 & (Selector7)) # (!Selector8 & ((Selector7 & ((\register[27][5]~q ))) # (!Selector7 & (\register[19][5]~q ))))

	.dataa(Selector8),
	.datab(Selector7),
	.datac(\register[19][5]~q ),
	.datad(\register[27][5]~q ),
	.cin(gnd),
	.combout(\Mux58~7_combout ),
	.cout());
// synopsys translate_off
defparam \Mux58~7 .lut_mask = 16'hDC98;
defparam \Mux58~7 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X65_Y30_N2
cycloneive_lcell_comb \Mux58~8 (
// Equation(s):
// \Mux58~8_combout  = (Selector8 & ((\Mux58~7_combout  & ((\register[31][5]~q ))) # (!\Mux58~7_combout  & (\register[23][5]~q )))) # (!Selector8 & (((\Mux58~7_combout ))))

	.dataa(\register[23][5]~q ),
	.datab(Selector8),
	.datac(\register[31][5]~q ),
	.datad(\Mux58~7_combout ),
	.cin(gnd),
	.combout(\Mux58~8_combout ),
	.cout());
// synopsys translate_off
defparam \Mux58~8 .lut_mask = 16'hF388;
defparam \Mux58~8 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y38_N0
cycloneive_lcell_comb \register[29][5]~feeder (
// Equation(s):
// \register[29][5]~feeder_combout  = \register~90_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(\register~90_combout ),
	.cin(gnd),
	.combout(\register[29][5]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \register[29][5]~feeder .lut_mask = 16'hFF00;
defparam \register[29][5]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X61_Y38_N1
dffeas \register[29][5] (
	.clk(!CLK),
	.d(\register[29][5]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~28_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\register[29][5]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \register[29][5] .is_wysiwyg = "true";
defparam \register[29][5] .power_up = "low";
// synopsys translate_on

// Location: FF_X63_Y35_N25
dffeas \register[21][5] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\register~90_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~22_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\register[21][5]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \register[21][5] .is_wysiwyg = "true";
defparam \register[21][5] .power_up = "low";
// synopsys translate_on

// Location: FF_X62_Y35_N19
dffeas \register[17][5] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\register~90_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~26_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\register[17][5]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \register[17][5] .is_wysiwyg = "true";
defparam \register[17][5] .power_up = "low";
// synopsys translate_on

// Location: FF_X62_Y36_N19
dffeas \register[25][5] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\register~90_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~24_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\register[25][5]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \register[25][5] .is_wysiwyg = "true";
defparam \register[25][5] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X62_Y36_N18
cycloneive_lcell_comb \Mux58~0 (
// Equation(s):
// \Mux58~0_combout  = (Selector8 & (((Selector7)))) # (!Selector8 & ((Selector7 & ((\register[25][5]~q ))) # (!Selector7 & (\register[17][5]~q ))))

	.dataa(Selector8),
	.datab(\register[17][5]~q ),
	.datac(\register[25][5]~q ),
	.datad(Selector7),
	.cin(gnd),
	.combout(\Mux58~0_combout ),
	.cout());
// synopsys translate_off
defparam \Mux58~0 .lut_mask = 16'hFA44;
defparam \Mux58~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X63_Y35_N24
cycloneive_lcell_comb \Mux58~1 (
// Equation(s):
// \Mux58~1_combout  = (Selector8 & ((\Mux58~0_combout  & (\register[29][5]~q )) # (!\Mux58~0_combout  & ((\register[21][5]~q ))))) # (!Selector8 & (((\Mux58~0_combout ))))

	.dataa(Selector8),
	.datab(\register[29][5]~q ),
	.datac(\register[21][5]~q ),
	.datad(\Mux58~0_combout ),
	.cin(gnd),
	.combout(\Mux58~1_combout ),
	.cout());
// synopsys translate_off
defparam \Mux58~1 .lut_mask = 16'hDDA0;
defparam \Mux58~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X68_Y38_N31
dffeas \register[26][5] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\register~90_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~54_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\register[26][5]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \register[26][5] .is_wysiwyg = "true";
defparam \register[26][5] .power_up = "low";
// synopsys translate_on

// Location: FF_X67_Y39_N31
dffeas \register[30][5] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\register~90_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~56_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\register[30][5]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \register[30][5] .is_wysiwyg = "true";
defparam \register[30][5] .power_up = "low";
// synopsys translate_on

// Location: FF_X68_Y38_N21
dffeas \register[18][5] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\register~90_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~33_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\register[18][5]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \register[18][5] .is_wysiwyg = "true";
defparam \register[18][5] .power_up = "low";
// synopsys translate_on

// Location: FF_X69_Y37_N11
dffeas \register[22][5] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\register~90_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~55_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\register[22][5]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \register[22][5] .is_wysiwyg = "true";
defparam \register[22][5] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X68_Y38_N20
cycloneive_lcell_comb \Mux58~2 (
// Equation(s):
// \Mux58~2_combout  = (Selector7 & (Selector8)) # (!Selector7 & ((Selector8 & ((\register[22][5]~q ))) # (!Selector8 & (\register[18][5]~q ))))

	.dataa(Selector7),
	.datab(Selector8),
	.datac(\register[18][5]~q ),
	.datad(\register[22][5]~q ),
	.cin(gnd),
	.combout(\Mux58~2_combout ),
	.cout());
// synopsys translate_off
defparam \Mux58~2 .lut_mask = 16'hDC98;
defparam \Mux58~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X67_Y39_N30
cycloneive_lcell_comb \Mux58~3 (
// Equation(s):
// \Mux58~3_combout  = (Selector7 & ((\Mux58~2_combout  & ((\register[30][5]~q ))) # (!\Mux58~2_combout  & (\register[26][5]~q )))) # (!Selector7 & (((\Mux58~2_combout ))))

	.dataa(Selector7),
	.datab(\register[26][5]~q ),
	.datac(\register[30][5]~q ),
	.datad(\Mux58~2_combout ),
	.cin(gnd),
	.combout(\Mux58~3_combout ),
	.cout());
// synopsys translate_off
defparam \Mux58~3 .lut_mask = 16'hF588;
defparam \Mux58~3 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X69_Y38_N30
cycloneive_lcell_comb \register[20][5]~feeder (
// Equation(s):
// \register[20][5]~feeder_combout  = \register~90_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(\register~90_combout ),
	.cin(gnd),
	.combout(\register[20][5]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \register[20][5]~feeder .lut_mask = 16'hFF00;
defparam \register[20][5]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X69_Y38_N31
dffeas \register[20][5] (
	.clk(!CLK),
	.d(\register[20][5]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~35_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\register[20][5]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \register[20][5] .is_wysiwyg = "true";
defparam \register[20][5] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X70_Y38_N14
cycloneive_lcell_comb \Mux58~4 (
// Equation(s):
// \Mux58~4_combout  = (Selector8 & (((\register[20][5]~q ) # (Selector7)))) # (!Selector8 & (\register[16][5]~q  & ((!Selector7))))

	.dataa(\register[16][5]~q ),
	.datab(\register[20][5]~q ),
	.datac(Selector8),
	.datad(Selector7),
	.cin(gnd),
	.combout(\Mux58~4_combout ),
	.cout());
// synopsys translate_off
defparam \Mux58~4 .lut_mask = 16'hF0CA;
defparam \Mux58~4 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X70_Y38_N18
cycloneive_lcell_comb \register[24][5]~feeder (
// Equation(s):
// \register[24][5]~feeder_combout  = \register~90_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(\register~90_combout ),
	.datad(gnd),
	.cin(gnd),
	.combout(\register[24][5]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \register[24][5]~feeder .lut_mask = 16'hF0F0;
defparam \register[24][5]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X70_Y38_N19
dffeas \register[24][5] (
	.clk(!CLK),
	.d(\register[24][5]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~34_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\register[24][5]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \register[24][5] .is_wysiwyg = "true";
defparam \register[24][5] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X66_Y36_N26
cycloneive_lcell_comb \Mux58~5 (
// Equation(s):
// \Mux58~5_combout  = (Selector7 & ((\Mux58~4_combout  & (\register[28][5]~q )) # (!\Mux58~4_combout  & ((\register[24][5]~q ))))) # (!Selector7 & (((\Mux58~4_combout ))))

	.dataa(\register[28][5]~q ),
	.datab(Selector7),
	.datac(\Mux58~4_combout ),
	.datad(\register[24][5]~q ),
	.cin(gnd),
	.combout(\Mux58~5_combout ),
	.cout());
// synopsys translate_off
defparam \Mux58~5 .lut_mask = 16'hBCB0;
defparam \Mux58~5 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X65_Y30_N16
cycloneive_lcell_comb \Mux58~6 (
// Equation(s):
// \Mux58~6_combout  = (Selector10 & (Selector91)) # (!Selector10 & ((Selector91 & (\Mux58~3_combout )) # (!Selector91 & ((\Mux58~5_combout )))))

	.dataa(Selector10),
	.datab(Selector91),
	.datac(\Mux58~3_combout ),
	.datad(\Mux58~5_combout ),
	.cin(gnd),
	.combout(\Mux58~6_combout ),
	.cout());
// synopsys translate_off
defparam \Mux58~6 .lut_mask = 16'hD9C8;
defparam \Mux58~6 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X66_Y31_N31
dffeas \register[7][5] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\register~90_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~43_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\register[7][5]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \register[7][5] .is_wysiwyg = "true";
defparam \register[7][5] .power_up = "low";
// synopsys translate_on

// Location: FF_X69_Y32_N1
dffeas \register[5][5] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\register~90_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~59_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\register[5][5]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \register[5][5] .is_wysiwyg = "true";
defparam \register[5][5] .power_up = "low";
// synopsys translate_on

// Location: FF_X69_Y32_N31
dffeas \register[4][5] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\register~90_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~60_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\register[4][5]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \register[4][5] .is_wysiwyg = "true";
defparam \register[4][5] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X69_Y32_N30
cycloneive_lcell_comb \Mux58~10 (
// Equation(s):
// \Mux58~10_combout  = (Selector10 & ((\register[5][5]~q ) # ((Selector91)))) # (!Selector10 & (((\register[4][5]~q  & !Selector91))))

	.dataa(Selector10),
	.datab(\register[5][5]~q ),
	.datac(\register[4][5]~q ),
	.datad(Selector91),
	.cin(gnd),
	.combout(\Mux58~10_combout ),
	.cout());
// synopsys translate_off
defparam \Mux58~10 .lut_mask = 16'hAAD8;
defparam \Mux58~10 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X66_Y31_N29
dffeas \register[6][5] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\register~90_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~58_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\register[6][5]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \register[6][5] .is_wysiwyg = "true";
defparam \register[6][5] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X66_Y31_N28
cycloneive_lcell_comb \Mux58~11 (
// Equation(s):
// \Mux58~11_combout  = (\Mux58~10_combout  & ((\register[7][5]~q ) # ((!Selector91)))) # (!\Mux58~10_combout  & (((\register[6][5]~q  & Selector91))))

	.dataa(\register[7][5]~q ),
	.datab(\Mux58~10_combout ),
	.datac(\register[6][5]~q ),
	.datad(Selector91),
	.cin(gnd),
	.combout(\Mux58~11_combout ),
	.cout());
// synopsys translate_off
defparam \Mux58~11 .lut_mask = 16'hB8CC;
defparam \Mux58~11 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X63_Y37_N15
dffeas \register[15][5] (
	.clk(!CLK),
	.d(\register~90_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~53_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\register[15][5]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \register[15][5] .is_wysiwyg = "true";
defparam \register[15][5] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X67_Y33_N2
cycloneive_lcell_comb \register[14][5]~feeder (
// Equation(s):
// \register[14][5]~feeder_combout  = \register~90_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(\register~90_combout ),
	.cin(gnd),
	.combout(\register[14][5]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \register[14][5]~feeder .lut_mask = 16'hFF00;
defparam \register[14][5]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X67_Y33_N3
dffeas \register[14][5] (
	.clk(!CLK),
	.d(\register[14][5]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~61_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\register[14][5]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \register[14][5] .is_wysiwyg = "true";
defparam \register[14][5] .power_up = "low";
// synopsys translate_on

// Location: FF_X63_Y30_N15
dffeas \register[12][5] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\register~90_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~52_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\register[12][5]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \register[12][5] .is_wysiwyg = "true";
defparam \register[12][5] .power_up = "low";
// synopsys translate_on

// Location: FF_X63_Y30_N17
dffeas \register[13][5] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\register~90_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~62_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\register[13][5]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \register[13][5] .is_wysiwyg = "true";
defparam \register[13][5] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X63_Y30_N16
cycloneive_lcell_comb \Mux58~17 (
// Equation(s):
// \Mux58~17_combout  = (Selector91 & (((Selector10)))) # (!Selector91 & ((Selector10 & ((\register[13][5]~q ))) # (!Selector10 & (\register[12][5]~q ))))

	.dataa(Selector91),
	.datab(\register[12][5]~q ),
	.datac(\register[13][5]~q ),
	.datad(Selector10),
	.cin(gnd),
	.combout(\Mux58~17_combout ),
	.cout());
// synopsys translate_off
defparam \Mux58~17 .lut_mask = 16'hFA44;
defparam \Mux58~17 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X67_Y33_N24
cycloneive_lcell_comb \Mux58~18 (
// Equation(s):
// \Mux58~18_combout  = (\Mux58~17_combout  & ((\register[15][5]~q ) # ((!Selector91)))) # (!\Mux58~17_combout  & (((\register[14][5]~q  & Selector91))))

	.dataa(\register[15][5]~q ),
	.datab(\register[14][5]~q ),
	.datac(\Mux58~17_combout ),
	.datad(Selector91),
	.cin(gnd),
	.combout(\Mux58~18_combout ),
	.cout());
// synopsys translate_off
defparam \Mux58~18 .lut_mask = 16'hACF0;
defparam \Mux58~18 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X66_Y34_N1
dffeas \register[2][5] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\register~90_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~50_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\register[2][5]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \register[2][5] .is_wysiwyg = "true";
defparam \register[2][5] .power_up = "low";
// synopsys translate_on

// Location: FF_X70_Y34_N27
dffeas \register[1][5] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\register~90_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~49_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\register[1][5]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \register[1][5] .is_wysiwyg = "true";
defparam \register[1][5] .power_up = "low";
// synopsys translate_on

// Location: FF_X70_Y34_N29
dffeas \register[3][5] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\register~90_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~48_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\register[3][5]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \register[3][5] .is_wysiwyg = "true";
defparam \register[3][5] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X70_Y34_N26
cycloneive_lcell_comb \Mux58~14 (
// Equation(s):
// \Mux58~14_combout  = (Selector9 & ((plif_ifidinstr_l_17 & ((\register[3][5]~q ))) # (!plif_ifidinstr_l_17 & (\register[1][5]~q )))) # (!Selector9 & (((\register[1][5]~q ))))

	.dataa(Selector9),
	.datab(plif_ifidinstr_l_17),
	.datac(\register[1][5]~q ),
	.datad(\register[3][5]~q ),
	.cin(gnd),
	.combout(\Mux58~14_combout ),
	.cout());
// synopsys translate_off
defparam \Mux58~14 .lut_mask = 16'hF870;
defparam \Mux58~14 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X65_Y30_N14
cycloneive_lcell_comb \Mux58~15 (
// Equation(s):
// \Mux58~15_combout  = (Selector10 & (((\Mux58~14_combout )))) # (!Selector10 & (\register[2][5]~q  & ((Selector91))))

	.dataa(Selector10),
	.datab(\register[2][5]~q ),
	.datac(\Mux58~14_combout ),
	.datad(Selector91),
	.cin(gnd),
	.combout(\Mux58~15_combout ),
	.cout());
// synopsys translate_off
defparam \Mux58~15 .lut_mask = 16'hE4A0;
defparam \Mux58~15 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X66_Y38_N21
dffeas \register[9][5] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\register~90_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~44_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\register[9][5]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \register[9][5] .is_wysiwyg = "true";
defparam \register[9][5] .power_up = "low";
// synopsys translate_on

// Location: FF_X66_Y38_N19
dffeas \register[11][5] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\register~90_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~47_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\register[11][5]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \register[11][5] .is_wysiwyg = "true";
defparam \register[11][5] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X66_Y38_N18
cycloneive_lcell_comb \Mux58~13 (
// Equation(s):
// \Mux58~13_combout  = (\Mux58~12_combout  & (((\register[11][5]~q ) # (!Selector10)))) # (!\Mux58~12_combout  & (\register[9][5]~q  & ((Selector10))))

	.dataa(\Mux58~12_combout ),
	.datab(\register[9][5]~q ),
	.datac(\register[11][5]~q ),
	.datad(Selector10),
	.cin(gnd),
	.combout(\Mux58~13_combout ),
	.cout());
// synopsys translate_off
defparam \Mux58~13 .lut_mask = 16'hE4AA;
defparam \Mux58~13 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X65_Y30_N28
cycloneive_lcell_comb \Mux58~16 (
// Equation(s):
// \Mux58~16_combout  = (Selector7 & ((Selector8) # ((\Mux58~13_combout )))) # (!Selector7 & (!Selector8 & (\Mux58~15_combout )))

	.dataa(Selector7),
	.datab(Selector8),
	.datac(\Mux58~15_combout ),
	.datad(\Mux58~13_combout ),
	.cin(gnd),
	.combout(\Mux58~16_combout ),
	.cout());
// synopsys translate_off
defparam \Mux58~16 .lut_mask = 16'hBA98;
defparam \Mux58~16 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X63_Y37_N28
cycloneive_lcell_comb \register~91 (
// Equation(s):
// \register~91_combout  = (WideOr01 & ((\wdat[2]~54_combout ) # ((plif_memwbregsrc_l_1 & plif_memwbrtnaddr_l_2))))

	.dataa(plif_memwbregsrc_l_1),
	.datab(plif_memwbrtnaddr_l_2),
	.datac(WideOr0),
	.datad(wdat_2),
	.cin(gnd),
	.combout(\register~91_combout ),
	.cout());
// synopsys translate_off
defparam \register~91 .lut_mask = 16'hF080;
defparam \register~91 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X62_Y31_N17
dffeas \register[23][2] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\register~91_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~37_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\register[23][2]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \register[23][2] .is_wysiwyg = "true";
defparam \register[23][2] .power_up = "low";
// synopsys translate_on

// Location: FF_X63_Y32_N31
dffeas \register[31][2] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\register~91_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~40_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\register[31][2]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \register[31][2] .is_wysiwyg = "true";
defparam \register[31][2] .power_up = "low";
// synopsys translate_on

// Location: FF_X62_Y31_N31
dffeas \register[19][2] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\register~91_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~39_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\register[19][2]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \register[19][2] .is_wysiwyg = "true";
defparam \register[19][2] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X61_Y31_N30
cycloneive_lcell_comb \register[27][2]~feeder (
// Equation(s):
// \register[27][2]~feeder_combout  = \register~91_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(\register~91_combout ),
	.cin(gnd),
	.combout(\register[27][2]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \register[27][2]~feeder .lut_mask = 16'hFF00;
defparam \register[27][2]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X61_Y31_N31
dffeas \register[27][2] (
	.clk(!CLK),
	.d(\register[27][2]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~38_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\register[27][2]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \register[27][2] .is_wysiwyg = "true";
defparam \register[27][2] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X62_Y31_N30
cycloneive_lcell_comb \Mux29~7 (
// Equation(s):
// \Mux29~7_combout  = (Selector3 & (Selector2)) # (!Selector3 & ((Selector2 & ((\register[27][2]~q ))) # (!Selector2 & (\register[19][2]~q ))))

	.dataa(Selector3),
	.datab(Selector2),
	.datac(\register[19][2]~q ),
	.datad(\register[27][2]~q ),
	.cin(gnd),
	.combout(\Mux29~7_combout ),
	.cout());
// synopsys translate_off
defparam \Mux29~7 .lut_mask = 16'hDC98;
defparam \Mux29~7 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X63_Y32_N30
cycloneive_lcell_comb \Mux29~8 (
// Equation(s):
// \Mux29~8_combout  = (Selector3 & ((\Mux29~7_combout  & ((\register[31][2]~q ))) # (!\Mux29~7_combout  & (\register[23][2]~q )))) # (!Selector3 & (((\Mux29~7_combout ))))

	.dataa(\register[23][2]~q ),
	.datab(Selector3),
	.datac(\register[31][2]~q ),
	.datad(\Mux29~7_combout ),
	.cin(gnd),
	.combout(\Mux29~8_combout ),
	.cout());
// synopsys translate_off
defparam \Mux29~8 .lut_mask = 16'hF388;
defparam \Mux29~8 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X63_Y33_N31
dffeas \register[29][2] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\register~91_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~28_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\register[29][2]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \register[29][2] .is_wysiwyg = "true";
defparam \register[29][2] .power_up = "low";
// synopsys translate_on

// Location: FF_X63_Y33_N5
dffeas \register[21][2] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\register~91_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~22_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\register[21][2]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \register[21][2] .is_wysiwyg = "true";
defparam \register[21][2] .power_up = "low";
// synopsys translate_on

// Location: FF_X60_Y34_N15
dffeas \register[25][2] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\register~91_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~24_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\register[25][2]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \register[25][2] .is_wysiwyg = "true";
defparam \register[25][2] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X60_Y34_N14
cycloneive_lcell_comb \Mux29~0 (
// Equation(s):
// \Mux29~0_combout  = (Selector3 & (((Selector2)))) # (!Selector3 & ((Selector2 & ((\register[25][2]~q ))) # (!Selector2 & (\register[17][2]~q ))))

	.dataa(\register[17][2]~q ),
	.datab(Selector3),
	.datac(\register[25][2]~q ),
	.datad(Selector2),
	.cin(gnd),
	.combout(\Mux29~0_combout ),
	.cout());
// synopsys translate_off
defparam \Mux29~0 .lut_mask = 16'hFC22;
defparam \Mux29~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X63_Y33_N4
cycloneive_lcell_comb \Mux29~1 (
// Equation(s):
// \Mux29~1_combout  = (Selector3 & ((\Mux29~0_combout  & (\register[29][2]~q )) # (!\Mux29~0_combout  & ((\register[21][2]~q ))))) # (!Selector3 & (((\Mux29~0_combout ))))

	.dataa(Selector3),
	.datab(\register[29][2]~q ),
	.datac(\register[21][2]~q ),
	.datad(\Mux29~0_combout ),
	.cin(gnd),
	.combout(\Mux29~1_combout ),
	.cout());
// synopsys translate_off
defparam \Mux29~1 .lut_mask = 16'hDDA0;
defparam \Mux29~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X65_Y38_N28
cycloneive_lcell_comb \register[24][2]~feeder (
// Equation(s):
// \register[24][2]~feeder_combout  = \register~91_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(\register~91_combout ),
	.datad(gnd),
	.cin(gnd),
	.combout(\register[24][2]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \register[24][2]~feeder .lut_mask = 16'hF0F0;
defparam \register[24][2]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X65_Y38_N29
dffeas \register[24][2] (
	.clk(!CLK),
	.d(\register[24][2]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~34_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\register[24][2]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \register[24][2] .is_wysiwyg = "true";
defparam \register[24][2] .power_up = "low";
// synopsys translate_on

// Location: FF_X65_Y38_N23
dffeas \register[28][2] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\register~91_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~57_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\register[28][2]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \register[28][2] .is_wysiwyg = "true";
defparam \register[28][2] .power_up = "low";
// synopsys translate_on

// Location: FF_X65_Y34_N23
dffeas \register[20][2] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\register~91_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~35_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\register[20][2]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \register[20][2] .is_wysiwyg = "true";
defparam \register[20][2] .power_up = "low";
// synopsys translate_on

// Location: FF_X65_Y34_N21
dffeas \register[16][2] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\register~91_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~36_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\register[16][2]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \register[16][2] .is_wysiwyg = "true";
defparam \register[16][2] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X65_Y34_N22
cycloneive_lcell_comb \Mux29~4 (
// Equation(s):
// \Mux29~4_combout  = (Selector2 & (Selector3)) # (!Selector2 & ((Selector3 & (\register[20][2]~q )) # (!Selector3 & ((\register[16][2]~q )))))

	.dataa(Selector2),
	.datab(Selector3),
	.datac(\register[20][2]~q ),
	.datad(\register[16][2]~q ),
	.cin(gnd),
	.combout(\Mux29~4_combout ),
	.cout());
// synopsys translate_off
defparam \Mux29~4 .lut_mask = 16'hD9C8;
defparam \Mux29~4 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X65_Y38_N22
cycloneive_lcell_comb \Mux29~5 (
// Equation(s):
// \Mux29~5_combout  = (Selector2 & ((\Mux29~4_combout  & ((\register[28][2]~q ))) # (!\Mux29~4_combout  & (\register[24][2]~q )))) # (!Selector2 & (((\Mux29~4_combout ))))

	.dataa(Selector2),
	.datab(\register[24][2]~q ),
	.datac(\register[28][2]~q ),
	.datad(\Mux29~4_combout ),
	.cin(gnd),
	.combout(\Mux29~5_combout ),
	.cout());
// synopsys translate_off
defparam \Mux29~5 .lut_mask = 16'hF588;
defparam \Mux29~5 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X68_Y37_N13
dffeas \register[30][2] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\register~91_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~56_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\register[30][2]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \register[30][2] .is_wysiwyg = "true";
defparam \register[30][2] .power_up = "low";
// synopsys translate_on

// Location: FF_X69_Y37_N25
dffeas \register[22][2] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\register~91_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~55_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\register[22][2]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \register[22][2] .is_wysiwyg = "true";
defparam \register[22][2] .power_up = "low";
// synopsys translate_on

// Location: FF_X69_Y37_N15
dffeas \register[18][2] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\register~91_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~33_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\register[18][2]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \register[18][2] .is_wysiwyg = "true";
defparam \register[18][2] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X69_Y37_N14
cycloneive_lcell_comb \Mux29~2 (
// Equation(s):
// \Mux29~2_combout  = (Selector2 & (((Selector3)))) # (!Selector2 & ((Selector3 & (\register[22][2]~q )) # (!Selector3 & ((\register[18][2]~q )))))

	.dataa(Selector2),
	.datab(\register[22][2]~q ),
	.datac(\register[18][2]~q ),
	.datad(Selector3),
	.cin(gnd),
	.combout(\Mux29~2_combout ),
	.cout());
// synopsys translate_off
defparam \Mux29~2 .lut_mask = 16'hEE50;
defparam \Mux29~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X68_Y37_N12
cycloneive_lcell_comb \Mux29~3 (
// Equation(s):
// \Mux29~3_combout  = (Selector2 & ((\Mux29~2_combout  & ((\register[30][2]~q ))) # (!\Mux29~2_combout  & (\register[26][2]~q )))) # (!Selector2 & (((\Mux29~2_combout ))))

	.dataa(\register[26][2]~q ),
	.datab(Selector2),
	.datac(\register[30][2]~q ),
	.datad(\Mux29~2_combout ),
	.cin(gnd),
	.combout(\Mux29~3_combout ),
	.cout());
// synopsys translate_off
defparam \Mux29~3 .lut_mask = 16'hF388;
defparam \Mux29~3 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X63_Y32_N16
cycloneive_lcell_comb \Mux29~6 (
// Equation(s):
// \Mux29~6_combout  = (Selector5 & (((Selector41)))) # (!Selector5 & ((Selector41 & ((\Mux29~3_combout ))) # (!Selector41 & (\Mux29~5_combout ))))

	.dataa(\Mux29~5_combout ),
	.datab(Selector5),
	.datac(Selector41),
	.datad(\Mux29~3_combout ),
	.cin(gnd),
	.combout(\Mux29~6_combout ),
	.cout());
// synopsys translate_off
defparam \Mux29~6 .lut_mask = 16'hF2C2;
defparam \Mux29~6 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X66_Y31_N19
dffeas \register[7][2] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\register~91_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~43_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\register[7][2]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \register[7][2] .is_wysiwyg = "true";
defparam \register[7][2] .power_up = "low";
// synopsys translate_on

// Location: FF_X66_Y31_N25
dffeas \register[6][2] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\register~91_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~58_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\register[6][2]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \register[6][2] .is_wysiwyg = "true";
defparam \register[6][2] .power_up = "low";
// synopsys translate_on

// Location: FF_X67_Y31_N3
dffeas \register[4][2] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\register~91_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~60_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\register[4][2]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \register[4][2] .is_wysiwyg = "true";
defparam \register[4][2] .power_up = "low";
// synopsys translate_on

// Location: FF_X67_Y31_N29
dffeas \register[5][2] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\register~91_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~59_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\register[5][2]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \register[5][2] .is_wysiwyg = "true";
defparam \register[5][2] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X67_Y31_N28
cycloneive_lcell_comb \Mux29~10 (
// Equation(s):
// \Mux29~10_combout  = (Selector41 & (((Selector5)))) # (!Selector41 & ((Selector5 & ((\register[5][2]~q ))) # (!Selector5 & (\register[4][2]~q ))))

	.dataa(Selector41),
	.datab(\register[4][2]~q ),
	.datac(\register[5][2]~q ),
	.datad(Selector5),
	.cin(gnd),
	.combout(\Mux29~10_combout ),
	.cout());
// synopsys translate_off
defparam \Mux29~10 .lut_mask = 16'hFA44;
defparam \Mux29~10 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X66_Y31_N24
cycloneive_lcell_comb \Mux29~11 (
// Equation(s):
// \Mux29~11_combout  = (Selector41 & ((\Mux29~10_combout  & (\register[7][2]~q )) # (!\Mux29~10_combout  & ((\register[6][2]~q ))))) # (!Selector41 & (((\Mux29~10_combout ))))

	.dataa(Selector41),
	.datab(\register[7][2]~q ),
	.datac(\register[6][2]~q ),
	.datad(\Mux29~10_combout ),
	.cin(gnd),
	.combout(\Mux29~11_combout ),
	.cout());
// synopsys translate_off
defparam \Mux29~11 .lut_mask = 16'hDDA0;
defparam \Mux29~11 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X63_Y37_N29
dffeas \register[15][2] (
	.clk(!CLK),
	.d(\register~91_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~53_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\register[15][2]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \register[15][2] .is_wysiwyg = "true";
defparam \register[15][2] .power_up = "low";
// synopsys translate_on

// Location: FF_X60_Y33_N19
dffeas \register[12][2] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\register~91_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~52_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\register[12][2]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \register[12][2] .is_wysiwyg = "true";
defparam \register[12][2] .power_up = "low";
// synopsys translate_on

// Location: FF_X60_Y33_N5
dffeas \register[13][2] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\register~91_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~62_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\register[13][2]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \register[13][2] .is_wysiwyg = "true";
defparam \register[13][2] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X60_Y33_N4
cycloneive_lcell_comb \Mux29~17 (
// Equation(s):
// \Mux29~17_combout  = (Selector5 & (((\register[13][2]~q ) # (Selector41)))) # (!Selector5 & (\register[12][2]~q  & ((!Selector41))))

	.dataa(Selector5),
	.datab(\register[12][2]~q ),
	.datac(\register[13][2]~q ),
	.datad(Selector41),
	.cin(gnd),
	.combout(\Mux29~17_combout ),
	.cout());
// synopsys translate_off
defparam \Mux29~17 .lut_mask = 16'hAAE4;
defparam \Mux29~17 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y34_N24
cycloneive_lcell_comb \register[14][2]~feeder (
// Equation(s):
// \register[14][2]~feeder_combout  = \register~91_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(\register~91_combout ),
	.datad(gnd),
	.cin(gnd),
	.combout(\register[14][2]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \register[14][2]~feeder .lut_mask = 16'hF0F0;
defparam \register[14][2]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X60_Y34_N25
dffeas \register[14][2] (
	.clk(!CLK),
	.d(\register[14][2]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~61_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\register[14][2]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \register[14][2] .is_wysiwyg = "true";
defparam \register[14][2] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X60_Y34_N18
cycloneive_lcell_comb \Mux29~18 (
// Equation(s):
// \Mux29~18_combout  = (Selector41 & ((\Mux29~17_combout  & (\register[15][2]~q )) # (!\Mux29~17_combout  & ((\register[14][2]~q ))))) # (!Selector41 & (((\Mux29~17_combout ))))

	.dataa(\register[15][2]~q ),
	.datab(Selector41),
	.datac(\Mux29~17_combout ),
	.datad(\register[14][2]~q ),
	.cin(gnd),
	.combout(\Mux29~18_combout ),
	.cout());
// synopsys translate_off
defparam \Mux29~18 .lut_mask = 16'hBCB0;
defparam \Mux29~18 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X68_Y33_N11
dffeas \register[2][2] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\register~91_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~50_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\register[2][2]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \register[2][2] .is_wysiwyg = "true";
defparam \register[2][2] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X63_Y32_N22
cycloneive_lcell_comb \Mux29~15 (
// Equation(s):
// \Mux29~15_combout  = (Selector5 & (\Mux29~14_combout )) # (!Selector5 & (((Selector41 & \register[2][2]~q ))))

	.dataa(\Mux29~14_combout ),
	.datab(Selector5),
	.datac(Selector41),
	.datad(\register[2][2]~q ),
	.cin(gnd),
	.combout(\Mux29~15_combout ),
	.cout());
// synopsys translate_off
defparam \Mux29~15 .lut_mask = 16'hB888;
defparam \Mux29~15 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X66_Y38_N9
dffeas \register[9][2] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\register~91_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~44_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\register[9][2]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \register[9][2] .is_wysiwyg = "true";
defparam \register[9][2] .power_up = "low";
// synopsys translate_on

// Location: FF_X66_Y38_N15
dffeas \register[11][2] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\register~91_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~47_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\register[11][2]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \register[11][2] .is_wysiwyg = "true";
defparam \register[11][2] .power_up = "low";
// synopsys translate_on

// Location: FF_X67_Y38_N23
dffeas \register[8][2] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\register~91_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~46_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\register[8][2]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \register[8][2] .is_wysiwyg = "true";
defparam \register[8][2] .power_up = "low";
// synopsys translate_on

// Location: FF_X67_Y38_N29
dffeas \register[10][2] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\register~91_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~45_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\register[10][2]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \register[10][2] .is_wysiwyg = "true";
defparam \register[10][2] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X67_Y38_N22
cycloneive_lcell_comb \Mux29~12 (
// Equation(s):
// \Mux29~12_combout  = (Selector5 & (Selector41)) # (!Selector5 & ((Selector41 & ((\register[10][2]~q ))) # (!Selector41 & (\register[8][2]~q ))))

	.dataa(Selector5),
	.datab(Selector41),
	.datac(\register[8][2]~q ),
	.datad(\register[10][2]~q ),
	.cin(gnd),
	.combout(\Mux29~12_combout ),
	.cout());
// synopsys translate_off
defparam \Mux29~12 .lut_mask = 16'hDC98;
defparam \Mux29~12 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X66_Y38_N14
cycloneive_lcell_comb \Mux29~13 (
// Equation(s):
// \Mux29~13_combout  = (Selector5 & ((\Mux29~12_combout  & ((\register[11][2]~q ))) # (!\Mux29~12_combout  & (\register[9][2]~q )))) # (!Selector5 & (((\Mux29~12_combout ))))

	.dataa(Selector5),
	.datab(\register[9][2]~q ),
	.datac(\register[11][2]~q ),
	.datad(\Mux29~12_combout ),
	.cin(gnd),
	.combout(\Mux29~13_combout ),
	.cout());
// synopsys translate_off
defparam \Mux29~13 .lut_mask = 16'hF588;
defparam \Mux29~13 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X63_Y32_N20
cycloneive_lcell_comb \Mux29~16 (
// Equation(s):
// \Mux29~16_combout  = (Selector2 & (((Selector3) # (\Mux29~13_combout )))) # (!Selector2 & (\Mux29~15_combout  & (!Selector3)))

	.dataa(\Mux29~15_combout ),
	.datab(Selector2),
	.datac(Selector3),
	.datad(\Mux29~13_combout ),
	.cin(gnd),
	.combout(\Mux29~16_combout ),
	.cout());
// synopsys translate_off
defparam \Mux29~16 .lut_mask = 16'hCEC2;
defparam \Mux29~16 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X63_Y37_N18
cycloneive_lcell_comb \register~92 (
// Equation(s):
// \register~92_combout  = (WideOr01 & ((\wdat[1]~56_combout ) # ((plif_memwbregsrc_l_1 & plif_memwbrtnaddr_l_1))))

	.dataa(plif_memwbregsrc_l_1),
	.datab(plif_memwbrtnaddr_l_1),
	.datac(WideOr0),
	.datad(wdat_1),
	.cin(gnd),
	.combout(\register~92_combout ),
	.cout());
// synopsys translate_off
defparam \register~92 .lut_mask = 16'hF080;
defparam \register~92 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X63_Y33_N13
dffeas \register[29][1] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\register~92_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~28_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\register[29][1]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \register[29][1] .is_wysiwyg = "true";
defparam \register[29][1] .power_up = "low";
// synopsys translate_on

// Location: FF_X62_Y33_N15
dffeas \register[21][1] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\register~92_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~22_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\register[21][1]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \register[21][1] .is_wysiwyg = "true";
defparam \register[21][1] .power_up = "low";
// synopsys translate_on

// Location: FF_X62_Y34_N15
dffeas \register[17][1] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\register~92_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~26_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\register[17][1]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \register[17][1] .is_wysiwyg = "true";
defparam \register[17][1] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X62_Y33_N14
cycloneive_lcell_comb \Mux30~0 (
// Equation(s):
// \Mux30~0_combout  = (Selector2 & (Selector3)) # (!Selector2 & ((Selector3 & (\register[21][1]~q )) # (!Selector3 & ((\register[17][1]~q )))))

	.dataa(Selector2),
	.datab(Selector3),
	.datac(\register[21][1]~q ),
	.datad(\register[17][1]~q ),
	.cin(gnd),
	.combout(\Mux30~0_combout ),
	.cout());
// synopsys translate_off
defparam \Mux30~0 .lut_mask = 16'hD9C8;
defparam \Mux30~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X63_Y31_N6
cycloneive_lcell_comb \register[25][1]~feeder (
// Equation(s):
// \register[25][1]~feeder_combout  = \register~92_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(\register~92_combout ),
	.datad(gnd),
	.cin(gnd),
	.combout(\register[25][1]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \register[25][1]~feeder .lut_mask = 16'hF0F0;
defparam \register[25][1]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X63_Y31_N7
dffeas \register[25][1] (
	.clk(!CLK),
	.d(\register[25][1]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~24_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\register[25][1]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \register[25][1] .is_wysiwyg = "true";
defparam \register[25][1] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X63_Y31_N12
cycloneive_lcell_comb \Mux30~1 (
// Equation(s):
// \Mux30~1_combout  = (Selector2 & ((\Mux30~0_combout  & (\register[29][1]~q )) # (!\Mux30~0_combout  & ((\register[25][1]~q ))))) # (!Selector2 & (((\Mux30~0_combout ))))

	.dataa(\register[29][1]~q ),
	.datab(Selector2),
	.datac(\Mux30~0_combout ),
	.datad(\register[25][1]~q ),
	.cin(gnd),
	.combout(\Mux30~1_combout ),
	.cout());
// synopsys translate_off
defparam \Mux30~1 .lut_mask = 16'hBCB0;
defparam \Mux30~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X66_Y35_N4
cycloneive_lcell_comb \register[30][1]~feeder (
// Equation(s):
// \register[30][1]~feeder_combout  = \register~92_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(\register~92_combout ),
	.cin(gnd),
	.combout(\register[30][1]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \register[30][1]~feeder .lut_mask = 16'hFF00;
defparam \register[30][1]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X66_Y35_N5
dffeas \register[30][1] (
	.clk(!CLK),
	.d(\register[30][1]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~56_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\register[30][1]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \register[30][1] .is_wysiwyg = "true";
defparam \register[30][1] .power_up = "low";
// synopsys translate_on

// Location: FF_X67_Y37_N3
dffeas \register[22][1] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\register~92_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~55_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\register[22][1]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \register[22][1] .is_wysiwyg = "true";
defparam \register[22][1] .power_up = "low";
// synopsys translate_on

// Location: FF_X67_Y37_N9
dffeas \register[18][1] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\register~92_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~33_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\register[18][1]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \register[18][1] .is_wysiwyg = "true";
defparam \register[18][1] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X67_Y37_N8
cycloneive_lcell_comb \Mux30~2 (
// Equation(s):
// \Mux30~2_combout  = (Selector3 & (((Selector2)))) # (!Selector3 & ((Selector2 & (\register[26][1]~q )) # (!Selector2 & ((\register[18][1]~q )))))

	.dataa(\register[26][1]~q ),
	.datab(Selector3),
	.datac(\register[18][1]~q ),
	.datad(Selector2),
	.cin(gnd),
	.combout(\Mux30~2_combout ),
	.cout());
// synopsys translate_off
defparam \Mux30~2 .lut_mask = 16'hEE30;
defparam \Mux30~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X66_Y36_N28
cycloneive_lcell_comb \Mux30~3 (
// Equation(s):
// \Mux30~3_combout  = (Selector3 & ((\Mux30~2_combout  & (\register[30][1]~q )) # (!\Mux30~2_combout  & ((\register[22][1]~q ))))) # (!Selector3 & (((\Mux30~2_combout ))))

	.dataa(Selector3),
	.datab(\register[30][1]~q ),
	.datac(\register[22][1]~q ),
	.datad(\Mux30~2_combout ),
	.cin(gnd),
	.combout(\Mux30~3_combout ),
	.cout());
// synopsys translate_off
defparam \Mux30~3 .lut_mask = 16'hDDA0;
defparam \Mux30~3 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X66_Y35_N14
cycloneive_lcell_comb \register[28][1]~feeder (
// Equation(s):
// \register[28][1]~feeder_combout  = \register~92_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(\register~92_combout ),
	.cin(gnd),
	.combout(\register[28][1]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \register[28][1]~feeder .lut_mask = 16'hFF00;
defparam \register[28][1]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X66_Y35_N15
dffeas \register[28][1] (
	.clk(!CLK),
	.d(\register[28][1]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~57_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\register[28][1]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \register[28][1] .is_wysiwyg = "true";
defparam \register[28][1] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X65_Y39_N6
cycloneive_lcell_comb \register[16][1]~feeder (
// Equation(s):
// \register[16][1]~feeder_combout  = \register~92_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(\register~92_combout ),
	.datad(gnd),
	.cin(gnd),
	.combout(\register[16][1]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \register[16][1]~feeder .lut_mask = 16'hF0F0;
defparam \register[16][1]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X65_Y39_N7
dffeas \register[16][1] (
	.clk(!CLK),
	.d(\register[16][1]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~36_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\register[16][1]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \register[16][1] .is_wysiwyg = "true";
defparam \register[16][1] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X70_Y35_N2
cycloneive_lcell_comb \Mux30~4 (
// Equation(s):
// \Mux30~4_combout  = (Selector3 & (((Selector2)))) # (!Selector3 & ((Selector2 & (\register[24][1]~q )) # (!Selector2 & ((\register[16][1]~q )))))

	.dataa(\register[24][1]~q ),
	.datab(Selector3),
	.datac(Selector2),
	.datad(\register[16][1]~q ),
	.cin(gnd),
	.combout(\Mux30~4_combout ),
	.cout());
// synopsys translate_off
defparam \Mux30~4 .lut_mask = 16'hE3E0;
defparam \Mux30~4 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X66_Y35_N28
cycloneive_lcell_comb \Mux30~5 (
// Equation(s):
// \Mux30~5_combout  = (\Mux30~4_combout  & (((\register[28][1]~q ) # (!Selector3)))) # (!\Mux30~4_combout  & (\register[20][1]~q  & ((Selector3))))

	.dataa(\register[20][1]~q ),
	.datab(\register[28][1]~q ),
	.datac(\Mux30~4_combout ),
	.datad(Selector3),
	.cin(gnd),
	.combout(\Mux30~5_combout ),
	.cout());
// synopsys translate_off
defparam \Mux30~5 .lut_mask = 16'hCAF0;
defparam \Mux30~5 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X65_Y31_N26
cycloneive_lcell_comb \Mux30~6 (
// Equation(s):
// \Mux30~6_combout  = (Selector41 & ((Selector5) # ((\Mux30~3_combout )))) # (!Selector41 & (!Selector5 & ((\Mux30~5_combout ))))

	.dataa(Selector41),
	.datab(Selector5),
	.datac(\Mux30~3_combout ),
	.datad(\Mux30~5_combout ),
	.cin(gnd),
	.combout(\Mux30~6_combout ),
	.cout());
// synopsys translate_off
defparam \Mux30~6 .lut_mask = 16'hB9A8;
defparam \Mux30~6 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X63_Y31_N10
cycloneive_lcell_comb \register[27][1]~feeder (
// Equation(s):
// \register[27][1]~feeder_combout  = \register~92_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(\register~92_combout ),
	.datad(gnd),
	.cin(gnd),
	.combout(\register[27][1]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \register[27][1]~feeder .lut_mask = 16'hF0F0;
defparam \register[27][1]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X63_Y31_N11
dffeas \register[27][1] (
	.clk(!CLK),
	.d(\register[27][1]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~38_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\register[27][1]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \register[27][1] .is_wysiwyg = "true";
defparam \register[27][1] .power_up = "low";
// synopsys translate_on

// Location: FF_X65_Y31_N21
dffeas \register[31][1] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\register~92_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~40_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\register[31][1]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \register[31][1] .is_wysiwyg = "true";
defparam \register[31][1] .power_up = "low";
// synopsys translate_on

// Location: FF_X62_Y31_N23
dffeas \register[19][1] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\register~92_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~39_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\register[19][1]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \register[19][1] .is_wysiwyg = "true";
defparam \register[19][1] .power_up = "low";
// synopsys translate_on

// Location: FF_X62_Y31_N29
dffeas \register[23][1] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\register~92_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~37_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\register[23][1]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \register[23][1] .is_wysiwyg = "true";
defparam \register[23][1] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X62_Y31_N22
cycloneive_lcell_comb \Mux30~7 (
// Equation(s):
// \Mux30~7_combout  = (Selector3 & ((Selector2) # ((\register[23][1]~q )))) # (!Selector3 & (!Selector2 & (\register[19][1]~q )))

	.dataa(Selector3),
	.datab(Selector2),
	.datac(\register[19][1]~q ),
	.datad(\register[23][1]~q ),
	.cin(gnd),
	.combout(\Mux30~7_combout ),
	.cout());
// synopsys translate_off
defparam \Mux30~7 .lut_mask = 16'hBA98;
defparam \Mux30~7 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X65_Y31_N20
cycloneive_lcell_comb \Mux30~8 (
// Equation(s):
// \Mux30~8_combout  = (Selector2 & ((\Mux30~7_combout  & ((\register[31][1]~q ))) # (!\Mux30~7_combout  & (\register[27][1]~q )))) # (!Selector2 & (((\Mux30~7_combout ))))

	.dataa(Selector2),
	.datab(\register[27][1]~q ),
	.datac(\register[31][1]~q ),
	.datad(\Mux30~7_combout ),
	.cin(gnd),
	.combout(\Mux30~8_combout ),
	.cout());
// synopsys translate_off
defparam \Mux30~8 .lut_mask = 16'hF588;
defparam \Mux30~8 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X70_Y34_N9
dffeas \register[3][1] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\register~92_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~48_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\register[3][1]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \register[3][1] .is_wysiwyg = "true";
defparam \register[3][1] .power_up = "low";
// synopsys translate_on

// Location: FF_X70_Y34_N31
dffeas \register[1][1] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\register~92_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~49_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\register[1][1]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \register[1][1] .is_wysiwyg = "true";
defparam \register[1][1] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X70_Y34_N30
cycloneive_lcell_comb \Mux30~14 (
// Equation(s):
// \Mux30~14_combout  = (Selector4 & ((plif_ifidinstr_l_22 & (\register[3][1]~q )) # (!plif_ifidinstr_l_22 & ((\register[1][1]~q ))))) # (!Selector4 & (((\register[1][1]~q ))))

	.dataa(Selector4),
	.datab(\register[3][1]~q ),
	.datac(\register[1][1]~q ),
	.datad(plif_ifidinstr_l_22),
	.cin(gnd),
	.combout(\Mux30~14_combout ),
	.cout());
// synopsys translate_off
defparam \Mux30~14 .lut_mask = 16'hD8F0;
defparam \Mux30~14 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X65_Y31_N8
cycloneive_lcell_comb \Mux30~15 (
// Equation(s):
// \Mux30~15_combout  = (Selector5 & (((\Mux30~14_combout )))) # (!Selector5 & (\register[2][1]~q  & (Selector41)))

	.dataa(\register[2][1]~q ),
	.datab(Selector5),
	.datac(Selector41),
	.datad(\Mux30~14_combout ),
	.cin(gnd),
	.combout(\Mux30~15_combout ),
	.cout());
// synopsys translate_off
defparam \Mux30~15 .lut_mask = 16'hEC20;
defparam \Mux30~15 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X66_Y31_N1
dffeas \register[6][1] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\register~92_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~58_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\register[6][1]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \register[6][1] .is_wysiwyg = "true";
defparam \register[6][1] .power_up = "low";
// synopsys translate_on

// Location: FF_X66_Y31_N7
dffeas \register[7][1] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\register~92_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~43_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\register[7][1]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \register[7][1] .is_wysiwyg = "true";
defparam \register[7][1] .power_up = "low";
// synopsys translate_on

// Location: FF_X67_Y31_N9
dffeas \register[5][1] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\register~92_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~59_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\register[5][1]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \register[5][1] .is_wysiwyg = "true";
defparam \register[5][1] .power_up = "low";
// synopsys translate_on

// Location: FF_X67_Y31_N31
dffeas \register[4][1] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\register~92_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~60_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\register[4][1]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \register[4][1] .is_wysiwyg = "true";
defparam \register[4][1] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X67_Y31_N30
cycloneive_lcell_comb \Mux30~12 (
// Equation(s):
// \Mux30~12_combout  = (Selector41 & (((Selector5)))) # (!Selector41 & ((Selector5 & (\register[5][1]~q )) # (!Selector5 & ((\register[4][1]~q )))))

	.dataa(Selector41),
	.datab(\register[5][1]~q ),
	.datac(\register[4][1]~q ),
	.datad(Selector5),
	.cin(gnd),
	.combout(\Mux30~12_combout ),
	.cout());
// synopsys translate_off
defparam \Mux30~12 .lut_mask = 16'hEE50;
defparam \Mux30~12 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X66_Y31_N6
cycloneive_lcell_comb \Mux30~13 (
// Equation(s):
// \Mux30~13_combout  = (Selector41 & ((\Mux30~12_combout  & ((\register[7][1]~q ))) # (!\Mux30~12_combout  & (\register[6][1]~q )))) # (!Selector41 & (((\Mux30~12_combout ))))

	.dataa(Selector41),
	.datab(\register[6][1]~q ),
	.datac(\register[7][1]~q ),
	.datad(\Mux30~12_combout ),
	.cin(gnd),
	.combout(\Mux30~13_combout ),
	.cout());
// synopsys translate_off
defparam \Mux30~13 .lut_mask = 16'hF588;
defparam \Mux30~13 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X65_Y31_N18
cycloneive_lcell_comb \Mux30~16 (
// Equation(s):
// \Mux30~16_combout  = (Selector2 & (((Selector3)))) # (!Selector2 & ((Selector3 & ((\Mux30~13_combout ))) # (!Selector3 & (\Mux30~15_combout ))))

	.dataa(Selector2),
	.datab(\Mux30~15_combout ),
	.datac(Selector3),
	.datad(\Mux30~13_combout ),
	.cin(gnd),
	.combout(\Mux30~16_combout ),
	.cout());
// synopsys translate_off
defparam \Mux30~16 .lut_mask = 16'hF4A4;
defparam \Mux30~16 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X66_Y38_N31
dffeas \register[11][1] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\register~92_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~47_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\register[11][1]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \register[11][1] .is_wysiwyg = "true";
defparam \register[11][1] .power_up = "low";
// synopsys translate_on

// Location: FF_X67_Y38_N17
dffeas \register[10][1] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\register~92_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~45_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\register[10][1]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \register[10][1] .is_wysiwyg = "true";
defparam \register[10][1] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X67_Y38_N16
cycloneive_lcell_comb \Mux30~10 (
// Equation(s):
// \Mux30~10_combout  = (Selector41 & (((\register[10][1]~q ) # (Selector5)))) # (!Selector41 & (\register[8][1]~q  & ((!Selector5))))

	.dataa(\register[8][1]~q ),
	.datab(Selector41),
	.datac(\register[10][1]~q ),
	.datad(Selector5),
	.cin(gnd),
	.combout(\Mux30~10_combout ),
	.cout());
// synopsys translate_off
defparam \Mux30~10 .lut_mask = 16'hCCE2;
defparam \Mux30~10 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X66_Y38_N1
dffeas \register[9][1] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\register~92_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~44_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\register[9][1]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \register[9][1] .is_wysiwyg = "true";
defparam \register[9][1] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X66_Y38_N0
cycloneive_lcell_comb \Mux30~11 (
// Equation(s):
// \Mux30~11_combout  = (\Mux30~10_combout  & ((\register[11][1]~q ) # ((!Selector5)))) # (!\Mux30~10_combout  & (((\register[9][1]~q  & Selector5))))

	.dataa(\register[11][1]~q ),
	.datab(\Mux30~10_combout ),
	.datac(\register[9][1]~q ),
	.datad(Selector5),
	.cin(gnd),
	.combout(\Mux30~11_combout ),
	.cout());
// synopsys translate_off
defparam \Mux30~11 .lut_mask = 16'hB8CC;
defparam \Mux30~11 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X63_Y30_N29
dffeas \register[13][1] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\register~92_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~62_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\register[13][1]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \register[13][1] .is_wysiwyg = "true";
defparam \register[13][1] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X63_Y30_N28
cycloneive_lcell_comb \Mux30~17 (
// Equation(s):
// \Mux30~17_combout  = (Selector41 & (((Selector5)))) # (!Selector41 & ((Selector5 & ((\register[13][1]~q ))) # (!Selector5 & (\register[12][1]~q ))))

	.dataa(\register[12][1]~q ),
	.datab(Selector41),
	.datac(\register[13][1]~q ),
	.datad(Selector5),
	.cin(gnd),
	.combout(\Mux30~17_combout ),
	.cout());
// synopsys translate_off
defparam \Mux30~17 .lut_mask = 16'hFC22;
defparam \Mux30~17 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y33_N8
cycloneive_lcell_comb \register[14][1]~feeder (
// Equation(s):
// \register[14][1]~feeder_combout  = \register~92_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(\register~92_combout ),
	.datad(gnd),
	.cin(gnd),
	.combout(\register[14][1]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \register[14][1]~feeder .lut_mask = 16'hF0F0;
defparam \register[14][1]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X62_Y33_N9
dffeas \register[14][1] (
	.clk(!CLK),
	.d(\register[14][1]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~61_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\register[14][1]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \register[14][1] .is_wysiwyg = "true";
defparam \register[14][1] .power_up = "low";
// synopsys translate_on

// Location: FF_X63_Y37_N19
dffeas \register[15][1] (
	.clk(!CLK),
	.d(\register~92_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~53_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\register[15][1]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \register[15][1] .is_wysiwyg = "true";
defparam \register[15][1] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X69_Y34_N16
cycloneive_lcell_comb \Mux30~18 (
// Equation(s):
// \Mux30~18_combout  = (\Mux30~17_combout  & (((\register[15][1]~q )) # (!Selector41))) # (!\Mux30~17_combout  & (Selector41 & (\register[14][1]~q )))

	.dataa(\Mux30~17_combout ),
	.datab(Selector41),
	.datac(\register[14][1]~q ),
	.datad(\register[15][1]~q ),
	.cin(gnd),
	.combout(\Mux30~18_combout ),
	.cout());
// synopsys translate_off
defparam \Mux30~18 .lut_mask = 16'hEA62;
defparam \Mux30~18 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y36_N18
cycloneive_lcell_comb \register~93 (
// Equation(s):
// \register~93_combout  = (WideOr01 & ((\wdat[0]~58_combout ) # ((plif_memwbrtnaddr_l_0 & plif_memwbregsrc_l_1))))

	.dataa(plif_memwbrtnaddr_l_0),
	.datab(plif_memwbregsrc_l_1),
	.datac(wdat_0),
	.datad(WideOr0),
	.cin(gnd),
	.combout(\register~93_combout ),
	.cout());
// synopsys translate_off
defparam \register~93 .lut_mask = 16'hF800;
defparam \register~93 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y38_N10
cycloneive_lcell_comb \register[29][0]~feeder (
// Equation(s):
// \register[29][0]~feeder_combout  = \register~93_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(\register~93_combout ),
	.cin(gnd),
	.combout(\register[29][0]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \register[29][0]~feeder .lut_mask = 16'hFF00;
defparam \register[29][0]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X61_Y38_N11
dffeas \register[29][0] (
	.clk(!CLK),
	.d(\register[29][0]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~28_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\register[29][0]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \register[29][0] .is_wysiwyg = "true";
defparam \register[29][0] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X59_Y35_N22
cycloneive_lcell_comb \register[25][0]~feeder (
// Equation(s):
// \register[25][0]~feeder_combout  = \register~93_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(\register~93_combout ),
	.datad(gnd),
	.cin(gnd),
	.combout(\register[25][0]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \register[25][0]~feeder .lut_mask = 16'hF0F0;
defparam \register[25][0]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X59_Y35_N23
dffeas \register[25][0] (
	.clk(!CLK),
	.d(\register[25][0]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~24_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\register[25][0]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \register[25][0] .is_wysiwyg = "true";
defparam \register[25][0] .power_up = "low";
// synopsys translate_on

// Location: FF_X62_Y35_N29
dffeas \register[17][0] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\register~93_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~26_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\register[17][0]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \register[17][0] .is_wysiwyg = "true";
defparam \register[17][0] .power_up = "low";
// synopsys translate_on

// Location: FF_X63_Y35_N27
dffeas \register[21][0] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\register~93_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~22_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\register[21][0]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \register[21][0] .is_wysiwyg = "true";
defparam \register[21][0] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X63_Y35_N26
cycloneive_lcell_comb \Mux63~0 (
// Equation(s):
// \Mux63~0_combout  = (Selector7 & (((Selector8)))) # (!Selector7 & ((Selector8 & ((\register[21][0]~q ))) # (!Selector8 & (\register[17][0]~q ))))

	.dataa(Selector7),
	.datab(\register[17][0]~q ),
	.datac(\register[21][0]~q ),
	.datad(Selector8),
	.cin(gnd),
	.combout(\Mux63~0_combout ),
	.cout());
// synopsys translate_off
defparam \Mux63~0 .lut_mask = 16'hFA44;
defparam \Mux63~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y35_N16
cycloneive_lcell_comb \Mux63~1 (
// Equation(s):
// \Mux63~1_combout  = (Selector7 & ((\Mux63~0_combout  & (\register[29][0]~q )) # (!\Mux63~0_combout  & ((\register[25][0]~q ))))) # (!Selector7 & (((\Mux63~0_combout ))))

	.dataa(Selector7),
	.datab(\register[29][0]~q ),
	.datac(\register[25][0]~q ),
	.datad(\Mux63~0_combout ),
	.cin(gnd),
	.combout(\Mux63~1_combout ),
	.cout());
// synopsys translate_off
defparam \Mux63~1 .lut_mask = 16'hDDA0;
defparam \Mux63~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X63_Y35_N16
cycloneive_lcell_comb \register[27][0]~feeder (
// Equation(s):
// \register[27][0]~feeder_combout  = \register~93_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(\register~93_combout ),
	.datad(gnd),
	.cin(gnd),
	.combout(\register[27][0]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \register[27][0]~feeder .lut_mask = 16'hF0F0;
defparam \register[27][0]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X63_Y35_N17
dffeas \register[27][0] (
	.clk(!CLK),
	.d(\register[27][0]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~38_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\register[27][0]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \register[27][0] .is_wysiwyg = "true";
defparam \register[27][0] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X61_Y38_N24
cycloneive_lcell_comb \register[31][0]~feeder (
// Equation(s):
// \register[31][0]~feeder_combout  = \register~93_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(\register~93_combout ),
	.cin(gnd),
	.combout(\register[31][0]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \register[31][0]~feeder .lut_mask = 16'hFF00;
defparam \register[31][0]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X61_Y38_N25
dffeas \register[31][0] (
	.clk(!CLK),
	.d(\register[31][0]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~40_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\register[31][0]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \register[31][0] .is_wysiwyg = "true";
defparam \register[31][0] .power_up = "low";
// synopsys translate_on

// Location: FF_X60_Y38_N23
dffeas \register[19][0] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\register~93_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~39_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\register[19][0]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \register[19][0] .is_wysiwyg = "true";
defparam \register[19][0] .power_up = "low";
// synopsys translate_on

// Location: FF_X62_Y38_N25
dffeas \register[23][0] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\register~93_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~37_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\register[23][0]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \register[23][0] .is_wysiwyg = "true";
defparam \register[23][0] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X62_Y38_N24
cycloneive_lcell_comb \Mux63~7 (
// Equation(s):
// \Mux63~7_combout  = (Selector8 & (((\register[23][0]~q ) # (Selector7)))) # (!Selector8 & (\register[19][0]~q  & ((!Selector7))))

	.dataa(Selector8),
	.datab(\register[19][0]~q ),
	.datac(\register[23][0]~q ),
	.datad(Selector7),
	.cin(gnd),
	.combout(\Mux63~7_combout ),
	.cout());
// synopsys translate_off
defparam \Mux63~7 .lut_mask = 16'hAAE4;
defparam \Mux63~7 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y38_N14
cycloneive_lcell_comb \Mux63~8 (
// Equation(s):
// \Mux63~8_combout  = (Selector7 & ((\Mux63~7_combout  & ((\register[31][0]~q ))) # (!\Mux63~7_combout  & (\register[27][0]~q )))) # (!Selector7 & (((\Mux63~7_combout ))))

	.dataa(Selector7),
	.datab(\register[27][0]~q ),
	.datac(\register[31][0]~q ),
	.datad(\Mux63~7_combout ),
	.cin(gnd),
	.combout(\Mux63~8_combout ),
	.cout());
// synopsys translate_off
defparam \Mux63~8 .lut_mask = 16'hF588;
defparam \Mux63~8 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X61_Y36_N25
dffeas \register[30][0] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\register~93_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~56_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\register[30][0]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \register[30][0] .is_wysiwyg = "true";
defparam \register[30][0] .power_up = "low";
// synopsys translate_on

// Location: FF_X69_Y39_N5
dffeas \register[18][0] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\register~93_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~33_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\register[18][0]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \register[18][0] .is_wysiwyg = "true";
defparam \register[18][0] .power_up = "low";
// synopsys translate_on

// Location: FF_X69_Y39_N31
dffeas \register[26][0] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\register~93_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~54_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\register[26][0]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \register[26][0] .is_wysiwyg = "true";
defparam \register[26][0] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X69_Y39_N30
cycloneive_lcell_comb \Mux63~2 (
// Equation(s):
// \Mux63~2_combout  = (Selector8 & (((Selector7)))) # (!Selector8 & ((Selector7 & ((\register[26][0]~q ))) # (!Selector7 & (\register[18][0]~q ))))

	.dataa(Selector8),
	.datab(\register[18][0]~q ),
	.datac(\register[26][0]~q ),
	.datad(Selector7),
	.cin(gnd),
	.combout(\Mux63~2_combout ),
	.cout());
// synopsys translate_off
defparam \Mux63~2 .lut_mask = 16'hFA44;
defparam \Mux63~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X69_Y37_N12
cycloneive_lcell_comb \Mux63~3 (
// Equation(s):
// \Mux63~3_combout  = (Selector8 & ((\Mux63~2_combout  & ((\register[30][0]~q ))) # (!\Mux63~2_combout  & (\register[22][0]~q )))) # (!Selector8 & (((\Mux63~2_combout ))))

	.dataa(\register[22][0]~q ),
	.datab(Selector8),
	.datac(\register[30][0]~q ),
	.datad(\Mux63~2_combout ),
	.cin(gnd),
	.combout(\Mux63~3_combout ),
	.cout());
// synopsys translate_off
defparam \Mux63~3 .lut_mask = 16'hF388;
defparam \Mux63~3 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X65_Y38_N3
dffeas \register[28][0] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\register~93_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~57_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\register[28][0]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \register[28][0] .is_wysiwyg = "true";
defparam \register[28][0] .power_up = "low";
// synopsys translate_on

// Location: FF_X65_Y38_N13
dffeas \register[24][0] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\register~93_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~34_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\register[24][0]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \register[24][0] .is_wysiwyg = "true";
defparam \register[24][0] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X66_Y36_N24
cycloneive_lcell_comb \register[16][0]~feeder (
// Equation(s):
// \register[16][0]~feeder_combout  = \register~93_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(\register~93_combout ),
	.cin(gnd),
	.combout(\register[16][0]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \register[16][0]~feeder .lut_mask = 16'hFF00;
defparam \register[16][0]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X66_Y36_N25
dffeas \register[16][0] (
	.clk(!CLK),
	.d(\register[16][0]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~36_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\register[16][0]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \register[16][0] .is_wysiwyg = "true";
defparam \register[16][0] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X65_Y38_N12
cycloneive_lcell_comb \Mux63~4 (
// Equation(s):
// \Mux63~4_combout  = (Selector8 & (Selector7)) # (!Selector8 & ((Selector7 & (\register[24][0]~q )) # (!Selector7 & ((\register[16][0]~q )))))

	.dataa(Selector8),
	.datab(Selector7),
	.datac(\register[24][0]~q ),
	.datad(\register[16][0]~q ),
	.cin(gnd),
	.combout(\Mux63~4_combout ),
	.cout());
// synopsys translate_off
defparam \Mux63~4 .lut_mask = 16'hD9C8;
defparam \Mux63~4 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X65_Y38_N2
cycloneive_lcell_comb \Mux63~5 (
// Equation(s):
// \Mux63~5_combout  = (Selector8 & ((\Mux63~4_combout  & ((\register[28][0]~q ))) # (!\Mux63~4_combout  & (\register[20][0]~q )))) # (!Selector8 & (((\Mux63~4_combout ))))

	.dataa(\register[20][0]~q ),
	.datab(Selector8),
	.datac(\register[28][0]~q ),
	.datad(\Mux63~4_combout ),
	.cin(gnd),
	.combout(\Mux63~5_combout ),
	.cout());
// synopsys translate_off
defparam \Mux63~5 .lut_mask = 16'hF388;
defparam \Mux63~5 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y35_N2
cycloneive_lcell_comb \Mux63~6 (
// Equation(s):
// \Mux63~6_combout  = (Selector91 & ((\Mux63~3_combout ) # ((Selector10)))) # (!Selector91 & (((\Mux63~5_combout  & !Selector10))))

	.dataa(\Mux63~3_combout ),
	.datab(\Mux63~5_combout ),
	.datac(Selector91),
	.datad(Selector10),
	.cin(gnd),
	.combout(\Mux63~6_combout ),
	.cout());
// synopsys translate_off
defparam \Mux63~6 .lut_mask = 16'hF0AC;
defparam \Mux63~6 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X63_Y40_N7
dffeas \register[11][0] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\register~93_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~47_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\register[11][0]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \register[11][0] .is_wysiwyg = "true";
defparam \register[11][0] .power_up = "low";
// synopsys translate_on

// Location: FF_X63_Y40_N25
dffeas \register[9][0] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\register~93_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~44_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\register[9][0]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \register[9][0] .is_wysiwyg = "true";
defparam \register[9][0] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X63_Y41_N0
cycloneive_lcell_comb \register[10][0]~feeder (
// Equation(s):
// \register[10][0]~feeder_combout  = \register~93_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(\register~93_combout ),
	.cin(gnd),
	.combout(\register[10][0]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \register[10][0]~feeder .lut_mask = 16'hFF00;
defparam \register[10][0]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X63_Y41_N1
dffeas \register[10][0] (
	.clk(!CLK),
	.d(\register[10][0]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~45_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\register[10][0]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \register[10][0] .is_wysiwyg = "true";
defparam \register[10][0] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X63_Y41_N4
cycloneive_lcell_comb \Mux63~10 (
// Equation(s):
// \Mux63~10_combout  = (Selector91 & (((\register[10][0]~q ) # (Selector10)))) # (!Selector91 & (\register[8][0]~q  & ((!Selector10))))

	.dataa(\register[8][0]~q ),
	.datab(\register[10][0]~q ),
	.datac(Selector91),
	.datad(Selector10),
	.cin(gnd),
	.combout(\Mux63~10_combout ),
	.cout());
// synopsys translate_off
defparam \Mux63~10 .lut_mask = 16'hF0CA;
defparam \Mux63~10 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X63_Y40_N24
cycloneive_lcell_comb \Mux63~11 (
// Equation(s):
// \Mux63~11_combout  = (Selector10 & ((\Mux63~10_combout  & (\register[11][0]~q )) # (!\Mux63~10_combout  & ((\register[9][0]~q ))))) # (!Selector10 & (((\Mux63~10_combout ))))

	.dataa(\register[11][0]~q ),
	.datab(Selector10),
	.datac(\register[9][0]~q ),
	.datad(\Mux63~10_combout ),
	.cin(gnd),
	.combout(\Mux63~11_combout ),
	.cout());
// synopsys translate_off
defparam \Mux63~11 .lut_mask = 16'hBBC0;
defparam \Mux63~11 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X62_Y32_N13
dffeas \register[6][0] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\register~93_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~58_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\register[6][0]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \register[6][0] .is_wysiwyg = "true";
defparam \register[6][0] .power_up = "low";
// synopsys translate_on

// Location: FF_X68_Y33_N31
dffeas \register[7][0] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\register~93_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~43_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\register[7][0]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \register[7][0] .is_wysiwyg = "true";
defparam \register[7][0] .power_up = "low";
// synopsys translate_on

// Location: FF_X67_Y32_N7
dffeas \register[4][0] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\register~93_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~60_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\register[4][0]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \register[4][0] .is_wysiwyg = "true";
defparam \register[4][0] .power_up = "low";
// synopsys translate_on

// Location: FF_X67_Y32_N17
dffeas \register[5][0] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\register~93_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~59_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\register[5][0]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \register[5][0] .is_wysiwyg = "true";
defparam \register[5][0] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X67_Y32_N6
cycloneive_lcell_comb \Mux63~12 (
// Equation(s):
// \Mux63~12_combout  = (Selector10 & ((Selector91) # ((\register[5][0]~q )))) # (!Selector10 & (!Selector91 & (\register[4][0]~q )))

	.dataa(Selector10),
	.datab(Selector91),
	.datac(\register[4][0]~q ),
	.datad(\register[5][0]~q ),
	.cin(gnd),
	.combout(\Mux63~12_combout ),
	.cout());
// synopsys translate_off
defparam \Mux63~12 .lut_mask = 16'hBA98;
defparam \Mux63~12 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X68_Y33_N30
cycloneive_lcell_comb \Mux63~13 (
// Equation(s):
// \Mux63~13_combout  = (Selector91 & ((\Mux63~12_combout  & ((\register[7][0]~q ))) # (!\Mux63~12_combout  & (\register[6][0]~q )))) # (!Selector91 & (((\Mux63~12_combout ))))

	.dataa(Selector91),
	.datab(\register[6][0]~q ),
	.datac(\register[7][0]~q ),
	.datad(\Mux63~12_combout ),
	.cin(gnd),
	.combout(\Mux63~13_combout ),
	.cout());
// synopsys translate_off
defparam \Mux63~13 .lut_mask = 16'hF588;
defparam \Mux63~13 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X68_Y33_N0
cycloneive_lcell_comb \register[2][0]~feeder (
// Equation(s):
// \register[2][0]~feeder_combout  = \register~93_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(\register~93_combout ),
	.datad(gnd),
	.cin(gnd),
	.combout(\register[2][0]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \register[2][0]~feeder .lut_mask = 16'hF0F0;
defparam \register[2][0]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X68_Y33_N1
dffeas \register[2][0] (
	.clk(!CLK),
	.d(\register[2][0]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~50_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\register[2][0]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \register[2][0] .is_wysiwyg = "true";
defparam \register[2][0] .power_up = "low";
// synopsys translate_on

// Location: FF_X65_Y36_N1
dffeas \register[3][0] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\register~93_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~48_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\register[3][0]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \register[3][0] .is_wysiwyg = "true";
defparam \register[3][0] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X65_Y36_N0
cycloneive_lcell_comb \Mux63~14 (
// Equation(s):
// \Mux63~14_combout  = (Selector10 & ((Selector91 & ((\register[3][0]~q ))) # (!Selector91 & (\register[1][0]~q ))))

	.dataa(\register[1][0]~q ),
	.datab(Selector10),
	.datac(\register[3][0]~q ),
	.datad(Selector91),
	.cin(gnd),
	.combout(\Mux63~14_combout ),
	.cout());
// synopsys translate_off
defparam \Mux63~14 .lut_mask = 16'hC088;
defparam \Mux63~14 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X66_Y33_N20
cycloneive_lcell_comb \Mux63~15 (
// Equation(s):
// \Mux63~15_combout  = (\Mux63~14_combout ) # ((!Selector10 & (Selector91 & \register[2][0]~q )))

	.dataa(Selector10),
	.datab(Selector91),
	.datac(\register[2][0]~q ),
	.datad(\Mux63~14_combout ),
	.cin(gnd),
	.combout(\Mux63~15_combout ),
	.cout());
// synopsys translate_off
defparam \Mux63~15 .lut_mask = 16'hFF40;
defparam \Mux63~15 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y35_N26
cycloneive_lcell_comb \Mux63~16 (
// Equation(s):
// \Mux63~16_combout  = (Selector7 & (Selector8)) # (!Selector7 & ((Selector8 & (\Mux63~13_combout )) # (!Selector8 & ((\Mux63~15_combout )))))

	.dataa(Selector7),
	.datab(Selector8),
	.datac(\Mux63~13_combout ),
	.datad(\Mux63~15_combout ),
	.cin(gnd),
	.combout(\Mux63~16_combout ),
	.cout());
// synopsys translate_off
defparam \Mux63~16 .lut_mask = 16'hD9C8;
defparam \Mux63~16 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X61_Y36_N19
dffeas \register[15][0] (
	.clk(!CLK),
	.d(\register~93_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~53_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\register[15][0]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \register[15][0] .is_wysiwyg = "true";
defparam \register[15][0] .power_up = "low";
// synopsys translate_on

// Location: FF_X62_Y32_N7
dffeas \register[14][0] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\register~93_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~61_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\register[14][0]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \register[14][0] .is_wysiwyg = "true";
defparam \register[14][0] .power_up = "low";
// synopsys translate_on

// Location: FF_X60_Y33_N23
dffeas \register[12][0] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\register~93_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~52_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\register[12][0]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \register[12][0] .is_wysiwyg = "true";
defparam \register[12][0] .power_up = "low";
// synopsys translate_on

// Location: FF_X60_Y33_N21
dffeas \register[13][0] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\register~93_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~62_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\register[13][0]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \register[13][0] .is_wysiwyg = "true";
defparam \register[13][0] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X60_Y33_N22
cycloneive_lcell_comb \Mux63~17 (
// Equation(s):
// \Mux63~17_combout  = (Selector10 & ((Selector91) # ((\register[13][0]~q )))) # (!Selector10 & (!Selector91 & (\register[12][0]~q )))

	.dataa(Selector10),
	.datab(Selector91),
	.datac(\register[12][0]~q ),
	.datad(\register[13][0]~q ),
	.cin(gnd),
	.combout(\Mux63~17_combout ),
	.cout());
// synopsys translate_off
defparam \Mux63~17 .lut_mask = 16'hBA98;
defparam \Mux63~17 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X65_Y34_N26
cycloneive_lcell_comb \Mux63~18 (
// Equation(s):
// \Mux63~18_combout  = (Selector91 & ((\Mux63~17_combout  & (\register[15][0]~q )) # (!\Mux63~17_combout  & ((\register[14][0]~q ))))) # (!Selector91 & (((\Mux63~17_combout ))))

	.dataa(\register[15][0]~q ),
	.datab(Selector91),
	.datac(\register[14][0]~q ),
	.datad(\Mux63~17_combout ),
	.cin(gnd),
	.combout(\Mux63~18_combout ),
	.cout());
// synopsys translate_off
defparam \Mux63~18 .lut_mask = 16'hBBC0;
defparam \Mux63~18 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X67_Y37_N2
cycloneive_lcell_comb \Mux62~2 (
// Equation(s):
// \Mux62~2_combout  = (Selector8 & (((\register[22][1]~q ) # (Selector7)))) # (!Selector8 & (\register[18][1]~q  & ((!Selector7))))

	.dataa(Selector8),
	.datab(\register[18][1]~q ),
	.datac(\register[22][1]~q ),
	.datad(Selector7),
	.cin(gnd),
	.combout(\Mux62~2_combout ),
	.cout());
// synopsys translate_off
defparam \Mux62~2 .lut_mask = 16'hAAE4;
defparam \Mux62~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X68_Y37_N10
cycloneive_lcell_comb \register[26][1]~feeder (
// Equation(s):
// \register[26][1]~feeder_combout  = \register~92_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(\register~92_combout ),
	.cin(gnd),
	.combout(\register[26][1]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \register[26][1]~feeder .lut_mask = 16'hFF00;
defparam \register[26][1]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X68_Y37_N11
dffeas \register[26][1] (
	.clk(!CLK),
	.d(\register[26][1]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~54_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\register[26][1]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \register[26][1] .is_wysiwyg = "true";
defparam \register[26][1] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X66_Y35_N30
cycloneive_lcell_comb \Mux62~3 (
// Equation(s):
// \Mux62~3_combout  = (Selector7 & ((\Mux62~2_combout  & (\register[30][1]~q )) # (!\Mux62~2_combout  & ((\register[26][1]~q ))))) # (!Selector7 & (\Mux62~2_combout ))

	.dataa(Selector7),
	.datab(\Mux62~2_combout ),
	.datac(\register[30][1]~q ),
	.datad(\register[26][1]~q ),
	.cin(gnd),
	.combout(\Mux62~3_combout ),
	.cout());
// synopsys translate_off
defparam \Mux62~3 .lut_mask = 16'hE6C4;
defparam \Mux62~3 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X65_Y39_N5
dffeas \register[20][1] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\register~92_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~35_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\register[20][1]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \register[20][1] .is_wysiwyg = "true";
defparam \register[20][1] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X65_Y39_N4
cycloneive_lcell_comb \Mux62~4 (
// Equation(s):
// \Mux62~4_combout  = (Selector7 & (Selector8)) # (!Selector7 & ((Selector8 & (\register[20][1]~q )) # (!Selector8 & ((\register[16][1]~q )))))

	.dataa(Selector7),
	.datab(Selector8),
	.datac(\register[20][1]~q ),
	.datad(\register[16][1]~q ),
	.cin(gnd),
	.combout(\Mux62~4_combout ),
	.cout());
// synopsys translate_off
defparam \Mux62~4 .lut_mask = 16'hD9C8;
defparam \Mux62~4 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X66_Y35_N0
cycloneive_lcell_comb \Mux62~5 (
// Equation(s):
// \Mux62~5_combout  = (\Mux62~4_combout  & (((\register[28][1]~q ) # (!Selector7)))) # (!\Mux62~4_combout  & (\register[24][1]~q  & ((Selector7))))

	.dataa(\register[24][1]~q ),
	.datab(\Mux62~4_combout ),
	.datac(\register[28][1]~q ),
	.datad(Selector7),
	.cin(gnd),
	.combout(\Mux62~5_combout ),
	.cout());
// synopsys translate_off
defparam \Mux62~5 .lut_mask = 16'hE2CC;
defparam \Mux62~5 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X66_Y35_N6
cycloneive_lcell_comb \Mux62~6 (
// Equation(s):
// \Mux62~6_combout  = (Selector10 & (((Selector91)))) # (!Selector10 & ((Selector91 & (\Mux62~3_combout )) # (!Selector91 & ((\Mux62~5_combout )))))

	.dataa(\Mux62~3_combout ),
	.datab(Selector10),
	.datac(Selector91),
	.datad(\Mux62~5_combout ),
	.cin(gnd),
	.combout(\Mux62~6_combout ),
	.cout());
// synopsys translate_off
defparam \Mux62~6 .lut_mask = 16'hE3E0;
defparam \Mux62~6 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y34_N14
cycloneive_lcell_comb \Mux62~0 (
// Equation(s):
// \Mux62~0_combout  = (Selector7 & ((Selector8) # ((\register[25][1]~q )))) # (!Selector7 & (!Selector8 & (\register[17][1]~q )))

	.dataa(Selector7),
	.datab(Selector8),
	.datac(\register[17][1]~q ),
	.datad(\register[25][1]~q ),
	.cin(gnd),
	.combout(\Mux62~0_combout ),
	.cout());
// synopsys translate_off
defparam \Mux62~0 .lut_mask = 16'hBA98;
defparam \Mux62~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X63_Y33_N12
cycloneive_lcell_comb \Mux62~1 (
// Equation(s):
// \Mux62~1_combout  = (Selector8 & ((\Mux62~0_combout  & ((\register[29][1]~q ))) # (!\Mux62~0_combout  & (\register[21][1]~q )))) # (!Selector8 & (((\Mux62~0_combout ))))

	.dataa(Selector8),
	.datab(\register[21][1]~q ),
	.datac(\register[29][1]~q ),
	.datad(\Mux62~0_combout ),
	.cin(gnd),
	.combout(\Mux62~1_combout ),
	.cout());
// synopsys translate_off
defparam \Mux62~1 .lut_mask = 16'hF588;
defparam \Mux62~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X63_Y31_N28
cycloneive_lcell_comb \Mux62~7 (
// Equation(s):
// \Mux62~7_combout  = (Selector7 & ((\register[27][1]~q ) # ((Selector8)))) # (!Selector7 & (((!Selector8 & \register[19][1]~q ))))

	.dataa(\register[27][1]~q ),
	.datab(Selector7),
	.datac(Selector8),
	.datad(\register[19][1]~q ),
	.cin(gnd),
	.combout(\Mux62~7_combout ),
	.cout());
// synopsys translate_off
defparam \Mux62~7 .lut_mask = 16'hCBC8;
defparam \Mux62~7 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y31_N28
cycloneive_lcell_comb \Mux62~8 (
// Equation(s):
// \Mux62~8_combout  = (Selector8 & ((\Mux62~7_combout  & (\register[31][1]~q )) # (!\Mux62~7_combout  & ((\register[23][1]~q ))))) # (!Selector8 & (((\Mux62~7_combout ))))

	.dataa(Selector8),
	.datab(\register[31][1]~q ),
	.datac(\register[23][1]~q ),
	.datad(\Mux62~7_combout ),
	.cin(gnd),
	.combout(\Mux62~8_combout ),
	.cout());
// synopsys translate_off
defparam \Mux62~8 .lut_mask = 16'hDDA0;
defparam \Mux62~8 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X67_Y31_N8
cycloneive_lcell_comb \Mux62~10 (
// Equation(s):
// \Mux62~10_combout  = (Selector91 & (((Selector10)))) # (!Selector91 & ((Selector10 & ((\register[5][1]~q ))) # (!Selector10 & (\register[4][1]~q ))))

	.dataa(\register[4][1]~q ),
	.datab(Selector91),
	.datac(\register[5][1]~q ),
	.datad(Selector10),
	.cin(gnd),
	.combout(\Mux62~10_combout ),
	.cout());
// synopsys translate_off
defparam \Mux62~10 .lut_mask = 16'hFC22;
defparam \Mux62~10 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X66_Y31_N0
cycloneive_lcell_comb \Mux62~11 (
// Equation(s):
// \Mux62~11_combout  = (Selector91 & ((\Mux62~10_combout  & ((\register[7][1]~q ))) # (!\Mux62~10_combout  & (\register[6][1]~q )))) # (!Selector91 & (\Mux62~10_combout ))

	.dataa(Selector91),
	.datab(\Mux62~10_combout ),
	.datac(\register[6][1]~q ),
	.datad(\register[7][1]~q ),
	.cin(gnd),
	.combout(\Mux62~11_combout ),
	.cout());
// synopsys translate_off
defparam \Mux62~11 .lut_mask = 16'hEC64;
defparam \Mux62~11 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X63_Y30_N27
dffeas \register[12][1] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\register~92_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~52_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\register[12][1]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \register[12][1] .is_wysiwyg = "true";
defparam \register[12][1] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X63_Y30_N26
cycloneive_lcell_comb \Mux62~17 (
// Equation(s):
// \Mux62~17_combout  = (Selector91 & (((Selector10)))) # (!Selector91 & ((Selector10 & (\register[13][1]~q )) # (!Selector10 & ((\register[12][1]~q )))))

	.dataa(Selector91),
	.datab(\register[13][1]~q ),
	.datac(\register[12][1]~q ),
	.datad(Selector10),
	.cin(gnd),
	.combout(\Mux62~17_combout ),
	.cout());
// synopsys translate_off
defparam \Mux62~17 .lut_mask = 16'hEE50;
defparam \Mux62~17 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y33_N2
cycloneive_lcell_comb \Mux62~18 (
// Equation(s):
// \Mux62~18_combout  = (Selector91 & ((\Mux62~17_combout  & (\register[15][1]~q )) # (!\Mux62~17_combout  & ((\register[14][1]~q ))))) # (!Selector91 & (((\Mux62~17_combout ))))

	.dataa(Selector91),
	.datab(\register[15][1]~q ),
	.datac(\register[14][1]~q ),
	.datad(\Mux62~17_combout ),
	.cin(gnd),
	.combout(\Mux62~18_combout ),
	.cout());
// synopsys translate_off
defparam \Mux62~18 .lut_mask = 16'hDDA0;
defparam \Mux62~18 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X67_Y38_N27
dffeas \register[8][1] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\register~92_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~46_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\register[8][1]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \register[8][1] .is_wysiwyg = "true";
defparam \register[8][1] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X67_Y38_N26
cycloneive_lcell_comb \Mux62~12 (
// Equation(s):
// \Mux62~12_combout  = (Selector10 & (((Selector91)))) # (!Selector10 & ((Selector91 & (\register[10][1]~q )) # (!Selector91 & ((\register[8][1]~q )))))

	.dataa(Selector10),
	.datab(\register[10][1]~q ),
	.datac(\register[8][1]~q ),
	.datad(Selector91),
	.cin(gnd),
	.combout(\Mux62~12_combout ),
	.cout());
// synopsys translate_off
defparam \Mux62~12 .lut_mask = 16'hEE50;
defparam \Mux62~12 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X66_Y38_N30
cycloneive_lcell_comb \Mux62~13 (
// Equation(s):
// \Mux62~13_combout  = (Selector10 & ((\Mux62~12_combout  & ((\register[11][1]~q ))) # (!\Mux62~12_combout  & (\register[9][1]~q )))) # (!Selector10 & (((\Mux62~12_combout ))))

	.dataa(Selector10),
	.datab(\register[9][1]~q ),
	.datac(\register[11][1]~q ),
	.datad(\Mux62~12_combout ),
	.cin(gnd),
	.combout(\Mux62~13_combout ),
	.cout());
// synopsys translate_off
defparam \Mux62~13 .lut_mask = 16'hF588;
defparam \Mux62~13 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X68_Y33_N13
dffeas \register[2][1] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\register~92_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~50_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\register[2][1]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \register[2][1] .is_wysiwyg = "true";
defparam \register[2][1] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X70_Y34_N8
cycloneive_lcell_comb \Mux62~14 (
// Equation(s):
// \Mux62~14_combout  = (Selector10 & ((Selector91 & ((\register[3][1]~q ))) # (!Selector91 & (\register[1][1]~q ))))

	.dataa(\register[1][1]~q ),
	.datab(Selector91),
	.datac(\register[3][1]~q ),
	.datad(Selector10),
	.cin(gnd),
	.combout(\Mux62~14_combout ),
	.cout());
// synopsys translate_off
defparam \Mux62~14 .lut_mask = 16'hE200;
defparam \Mux62~14 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X68_Y33_N12
cycloneive_lcell_comb \Mux62~15 (
// Equation(s):
// \Mux62~15_combout  = (\Mux62~14_combout ) # ((!Selector10 & (Selector91 & \register[2][1]~q )))

	.dataa(Selector10),
	.datab(Selector91),
	.datac(\register[2][1]~q ),
	.datad(\Mux62~14_combout ),
	.cin(gnd),
	.combout(\Mux62~15_combout ),
	.cout());
// synopsys translate_off
defparam \Mux62~15 .lut_mask = 16'hFF40;
defparam \Mux62~15 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y35_N18
cycloneive_lcell_comb \Mux62~16 (
// Equation(s):
// \Mux62~16_combout  = (Selector7 & ((Selector8) # ((\Mux62~13_combout )))) # (!Selector7 & (!Selector8 & ((\Mux62~15_combout ))))

	.dataa(Selector7),
	.datab(Selector8),
	.datac(\Mux62~13_combout ),
	.datad(\Mux62~15_combout ),
	.cin(gnd),
	.combout(\Mux62~16_combout ),
	.cout());
// synopsys translate_off
defparam \Mux62~16 .lut_mask = 16'hB9A8;
defparam \Mux62~16 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X63_Y37_N6
cycloneive_lcell_comb \register~94 (
// Equation(s):
// \register~94_combout  = (WideOr01 & ((\wdat[4]~60_combout ) # ((plif_memwbregsrc_l_1 & plif_memwbrtnaddr_l_4))))

	.dataa(plif_memwbregsrc_l_1),
	.datab(plif_memwbrtnaddr_l_4),
	.datac(WideOr0),
	.datad(wdat_4),
	.cin(gnd),
	.combout(\register~94_combout ),
	.cout());
// synopsys translate_off
defparam \register~94 .lut_mask = 16'hF080;
defparam \register~94 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y34_N26
cycloneive_lcell_comb \register[21][4]~feeder (
// Equation(s):
// \register[21][4]~feeder_combout  = \register~94_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(\register~94_combout ),
	.datad(gnd),
	.cin(gnd),
	.combout(\register[21][4]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \register[21][4]~feeder .lut_mask = 16'hF0F0;
defparam \register[21][4]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X59_Y34_N27
dffeas \register[21][4] (
	.clk(!CLK),
	.d(\register[21][4]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~22_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\register[21][4]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \register[21][4] .is_wysiwyg = "true";
defparam \register[21][4] .power_up = "low";
// synopsys translate_on

// Location: FF_X60_Y34_N17
dffeas \register[25][4] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\register~94_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~24_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\register[25][4]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \register[25][4] .is_wysiwyg = "true";
defparam \register[25][4] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X60_Y34_N16
cycloneive_lcell_comb \Mux27~0 (
// Equation(s):
// \Mux27~0_combout  = (Selector3 & (((Selector2)))) # (!Selector3 & ((Selector2 & ((\register[25][4]~q ))) # (!Selector2 & (\register[17][4]~q ))))

	.dataa(\register[17][4]~q ),
	.datab(Selector3),
	.datac(\register[25][4]~q ),
	.datad(Selector2),
	.cin(gnd),
	.combout(\Mux27~0_combout ),
	.cout());
// synopsys translate_off
defparam \Mux27~0 .lut_mask = 16'hFC22;
defparam \Mux27~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y41_N28
cycloneive_lcell_comb \register[29][4]~feeder (
// Equation(s):
// \register[29][4]~feeder_combout  = \register~94_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(\register~94_combout ),
	.cin(gnd),
	.combout(\register[29][4]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \register[29][4]~feeder .lut_mask = 16'hFF00;
defparam \register[29][4]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X60_Y41_N29
dffeas \register[29][4] (
	.clk(!CLK),
	.d(\register[29][4]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~28_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\register[29][4]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \register[29][4] .is_wysiwyg = "true";
defparam \register[29][4] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X59_Y34_N4
cycloneive_lcell_comb \Mux27~1 (
// Equation(s):
// \Mux27~1_combout  = (\Mux27~0_combout  & (((\register[29][4]~q ) # (!Selector3)))) # (!\Mux27~0_combout  & (\register[21][4]~q  & (Selector3)))

	.dataa(\register[21][4]~q ),
	.datab(\Mux27~0_combout ),
	.datac(Selector3),
	.datad(\register[29][4]~q ),
	.cin(gnd),
	.combout(\Mux27~1_combout ),
	.cout());
// synopsys translate_off
defparam \Mux27~1 .lut_mask = 16'hEC2C;
defparam \Mux27~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y38_N30
cycloneive_lcell_comb \register[23][4]~feeder (
// Equation(s):
// \register[23][4]~feeder_combout  = \register~94_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(\register~94_combout ),
	.cin(gnd),
	.combout(\register[23][4]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \register[23][4]~feeder .lut_mask = 16'hFF00;
defparam \register[23][4]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X62_Y38_N31
dffeas \register[23][4] (
	.clk(!CLK),
	.d(\register[23][4]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~37_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\register[23][4]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \register[23][4] .is_wysiwyg = "true";
defparam \register[23][4] .power_up = "low";
// synopsys translate_on

// Location: FF_X62_Y39_N15
dffeas \register[31][4] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\register~94_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~40_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\register[31][4]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \register[31][4] .is_wysiwyg = "true";
defparam \register[31][4] .power_up = "low";
// synopsys translate_on

// Location: FF_X60_Y37_N17
dffeas \register[19][4] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\register~94_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~39_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\register[19][4]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \register[19][4] .is_wysiwyg = "true";
defparam \register[19][4] .power_up = "low";
// synopsys translate_on

// Location: FF_X62_Y39_N25
dffeas \register[27][4] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\register~94_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~38_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\register[27][4]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \register[27][4] .is_wysiwyg = "true";
defparam \register[27][4] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X62_Y39_N24
cycloneive_lcell_comb \Mux27~7 (
// Equation(s):
// \Mux27~7_combout  = (Selector3 & (((Selector2)))) # (!Selector3 & ((Selector2 & ((\register[27][4]~q ))) # (!Selector2 & (\register[19][4]~q ))))

	.dataa(Selector3),
	.datab(\register[19][4]~q ),
	.datac(\register[27][4]~q ),
	.datad(Selector2),
	.cin(gnd),
	.combout(\Mux27~7_combout ),
	.cout());
// synopsys translate_off
defparam \Mux27~7 .lut_mask = 16'hFA44;
defparam \Mux27~7 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y39_N14
cycloneive_lcell_comb \Mux27~8 (
// Equation(s):
// \Mux27~8_combout  = (Selector3 & ((\Mux27~7_combout  & ((\register[31][4]~q ))) # (!\Mux27~7_combout  & (\register[23][4]~q )))) # (!Selector3 & (((\Mux27~7_combout ))))

	.dataa(Selector3),
	.datab(\register[23][4]~q ),
	.datac(\register[31][4]~q ),
	.datad(\Mux27~7_combout ),
	.cin(gnd),
	.combout(\Mux27~8_combout ),
	.cout());
// synopsys translate_off
defparam \Mux27~8 .lut_mask = 16'hF588;
defparam \Mux27~8 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X68_Y37_N9
dffeas \register[26][4] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\register~94_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~54_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\register[26][4]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \register[26][4] .is_wysiwyg = "true";
defparam \register[26][4] .power_up = "low";
// synopsys translate_on

// Location: FF_X68_Y37_N3
dffeas \register[30][4] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\register~94_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~56_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\register[30][4]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \register[30][4] .is_wysiwyg = "true";
defparam \register[30][4] .power_up = "low";
// synopsys translate_on

// Location: FF_X67_Y37_N17
dffeas \register[18][4] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\register~94_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~33_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\register[18][4]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \register[18][4] .is_wysiwyg = "true";
defparam \register[18][4] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X67_Y37_N16
cycloneive_lcell_comb \Mux27~2 (
// Equation(s):
// \Mux27~2_combout  = (Selector3 & ((\register[22][4]~q ) # ((Selector2)))) # (!Selector3 & (((\register[18][4]~q  & !Selector2))))

	.dataa(\register[22][4]~q ),
	.datab(Selector3),
	.datac(\register[18][4]~q ),
	.datad(Selector2),
	.cin(gnd),
	.combout(\Mux27~2_combout ),
	.cout());
// synopsys translate_off
defparam \Mux27~2 .lut_mask = 16'hCCB8;
defparam \Mux27~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X68_Y37_N2
cycloneive_lcell_comb \Mux27~3 (
// Equation(s):
// \Mux27~3_combout  = (Selector2 & ((\Mux27~2_combout  & ((\register[30][4]~q ))) # (!\Mux27~2_combout  & (\register[26][4]~q )))) # (!Selector2 & (((\Mux27~2_combout ))))

	.dataa(Selector2),
	.datab(\register[26][4]~q ),
	.datac(\register[30][4]~q ),
	.datad(\Mux27~2_combout ),
	.cin(gnd),
	.combout(\Mux27~3_combout ),
	.cout());
// synopsys translate_off
defparam \Mux27~3 .lut_mask = 16'hF588;
defparam \Mux27~3 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X65_Y38_N5
dffeas \register[24][4] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\register~94_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~34_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\register[24][4]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \register[24][4] .is_wysiwyg = "true";
defparam \register[24][4] .power_up = "low";
// synopsys translate_on

// Location: FF_X65_Y37_N23
dffeas \register[20][4] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\register~94_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~35_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\register[20][4]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \register[20][4] .is_wysiwyg = "true";
defparam \register[20][4] .power_up = "low";
// synopsys translate_on

// Location: FF_X65_Y37_N29
dffeas \register[16][4] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\register~94_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~36_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\register[16][4]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \register[16][4] .is_wysiwyg = "true";
defparam \register[16][4] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X65_Y37_N22
cycloneive_lcell_comb \Mux27~4 (
// Equation(s):
// \Mux27~4_combout  = (Selector3 & ((Selector2) # ((\register[20][4]~q )))) # (!Selector3 & (!Selector2 & ((\register[16][4]~q ))))

	.dataa(Selector3),
	.datab(Selector2),
	.datac(\register[20][4]~q ),
	.datad(\register[16][4]~q ),
	.cin(gnd),
	.combout(\Mux27~4_combout ),
	.cout());
// synopsys translate_off
defparam \Mux27~4 .lut_mask = 16'hB9A8;
defparam \Mux27~4 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X65_Y38_N4
cycloneive_lcell_comb \Mux27~5 (
// Equation(s):
// \Mux27~5_combout  = (Selector2 & ((\Mux27~4_combout  & (\register[28][4]~q )) # (!\Mux27~4_combout  & ((\register[24][4]~q ))))) # (!Selector2 & (((\Mux27~4_combout ))))

	.dataa(\register[28][4]~q ),
	.datab(Selector2),
	.datac(\register[24][4]~q ),
	.datad(\Mux27~4_combout ),
	.cin(gnd),
	.combout(\Mux27~5_combout ),
	.cout());
// synopsys translate_off
defparam \Mux27~5 .lut_mask = 16'hBBC0;
defparam \Mux27~5 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y34_N18
cycloneive_lcell_comb \Mux27~6 (
// Equation(s):
// \Mux27~6_combout  = (Selector5 & (Selector41)) # (!Selector5 & ((Selector41 & (\Mux27~3_combout )) # (!Selector41 & ((\Mux27~5_combout )))))

	.dataa(Selector5),
	.datab(Selector41),
	.datac(\Mux27~3_combout ),
	.datad(\Mux27~5_combout ),
	.cin(gnd),
	.combout(\Mux27~6_combout ),
	.cout());
// synopsys translate_off
defparam \Mux27~6 .lut_mask = 16'hD9C8;
defparam \Mux27~6 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X66_Y31_N11
dffeas \register[7][4] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\register~94_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~43_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\register[7][4]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \register[7][4] .is_wysiwyg = "true";
defparam \register[7][4] .power_up = "low";
// synopsys translate_on

// Location: FF_X66_Y31_N17
dffeas \register[6][4] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\register~94_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~58_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\register[6][4]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \register[6][4] .is_wysiwyg = "true";
defparam \register[6][4] .power_up = "low";
// synopsys translate_on

// Location: FF_X67_Y31_N5
dffeas \register[5][4] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\register~94_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~59_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\register[5][4]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \register[5][4] .is_wysiwyg = "true";
defparam \register[5][4] .power_up = "low";
// synopsys translate_on

// Location: FF_X67_Y31_N19
dffeas \register[4][4] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\register~94_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~60_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\register[4][4]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \register[4][4] .is_wysiwyg = "true";
defparam \register[4][4] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X67_Y31_N18
cycloneive_lcell_comb \Mux27~10 (
// Equation(s):
// \Mux27~10_combout  = (Selector41 & (((Selector5)))) # (!Selector41 & ((Selector5 & (\register[5][4]~q )) # (!Selector5 & ((\register[4][4]~q )))))

	.dataa(Selector41),
	.datab(\register[5][4]~q ),
	.datac(\register[4][4]~q ),
	.datad(Selector5),
	.cin(gnd),
	.combout(\Mux27~10_combout ),
	.cout());
// synopsys translate_off
defparam \Mux27~10 .lut_mask = 16'hEE50;
defparam \Mux27~10 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X66_Y31_N16
cycloneive_lcell_comb \Mux27~11 (
// Equation(s):
// \Mux27~11_combout  = (Selector41 & ((\Mux27~10_combout  & (\register[7][4]~q )) # (!\Mux27~10_combout  & ((\register[6][4]~q ))))) # (!Selector41 & (((\Mux27~10_combout ))))

	.dataa(\register[7][4]~q ),
	.datab(Selector41),
	.datac(\register[6][4]~q ),
	.datad(\Mux27~10_combout ),
	.cin(gnd),
	.combout(\Mux27~11_combout ),
	.cout());
// synopsys translate_off
defparam \Mux27~11 .lut_mask = 16'hBBC0;
defparam \Mux27~11 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X60_Y34_N23
dffeas \register[14][4] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\register~94_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~61_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\register[14][4]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \register[14][4] .is_wysiwyg = "true";
defparam \register[14][4] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X63_Y37_N0
cycloneive_lcell_comb \register[15][4]~feeder (
// Equation(s):
// \register[15][4]~feeder_combout  = \register~94_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(\register~94_combout ),
	.cin(gnd),
	.combout(\register[15][4]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \register[15][4]~feeder .lut_mask = 16'hFF00;
defparam \register[15][4]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X63_Y37_N1
dffeas \register[15][4] (
	.clk(!CLK),
	.d(\register[15][4]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~53_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\register[15][4]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \register[15][4] .is_wysiwyg = "true";
defparam \register[15][4] .power_up = "low";
// synopsys translate_on

// Location: FF_X60_Y33_N3
dffeas \register[12][4] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\register~94_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~52_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\register[12][4]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \register[12][4] .is_wysiwyg = "true";
defparam \register[12][4] .power_up = "low";
// synopsys translate_on

// Location: FF_X60_Y33_N13
dffeas \register[13][4] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\register~94_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~62_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\register[13][4]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \register[13][4] .is_wysiwyg = "true";
defparam \register[13][4] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X60_Y33_N12
cycloneive_lcell_comb \Mux27~17 (
// Equation(s):
// \Mux27~17_combout  = (Selector5 & (((\register[13][4]~q ) # (Selector41)))) # (!Selector5 & (\register[12][4]~q  & ((!Selector41))))

	.dataa(Selector5),
	.datab(\register[12][4]~q ),
	.datac(\register[13][4]~q ),
	.datad(Selector41),
	.cin(gnd),
	.combout(\Mux27~17_combout ),
	.cout());
// synopsys translate_off
defparam \Mux27~17 .lut_mask = 16'hAAE4;
defparam \Mux27~17 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y34_N28
cycloneive_lcell_comb \Mux27~18 (
// Equation(s):
// \Mux27~18_combout  = (Selector41 & ((\Mux27~17_combout  & ((\register[15][4]~q ))) # (!\Mux27~17_combout  & (\register[14][4]~q )))) # (!Selector41 & (((\Mux27~17_combout ))))

	.dataa(\register[14][4]~q ),
	.datab(\register[15][4]~q ),
	.datac(Selector41),
	.datad(\Mux27~17_combout ),
	.cin(gnd),
	.combout(\Mux27~18_combout ),
	.cout());
// synopsys translate_off
defparam \Mux27~18 .lut_mask = 16'hCFA0;
defparam \Mux27~18 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X70_Y34_N3
dffeas \register[1][4] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\register~94_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~49_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\register[1][4]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \register[1][4] .is_wysiwyg = "true";
defparam \register[1][4] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X70_Y34_N2
cycloneive_lcell_comb \Mux27~14 (
// Equation(s):
// \Mux27~14_combout  = (plif_ifidinstr_l_22 & ((Selector4 & (\register[3][4]~q )) # (!Selector4 & ((\register[1][4]~q ))))) # (!plif_ifidinstr_l_22 & (((\register[1][4]~q ))))

	.dataa(\register[3][4]~q ),
	.datab(plif_ifidinstr_l_22),
	.datac(\register[1][4]~q ),
	.datad(Selector4),
	.cin(gnd),
	.combout(\Mux27~14_combout ),
	.cout());
// synopsys translate_off
defparam \Mux27~14 .lut_mask = 16'hB8F0;
defparam \Mux27~14 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X67_Y34_N24
cycloneive_lcell_comb \Mux27~15 (
// Equation(s):
// \Mux27~15_combout  = (Selector5 & (((\Mux27~14_combout )))) # (!Selector5 & (\register[2][4]~q  & (Selector41)))

	.dataa(\register[2][4]~q ),
	.datab(Selector41),
	.datac(Selector5),
	.datad(\Mux27~14_combout ),
	.cin(gnd),
	.combout(\Mux27~15_combout ),
	.cout());
// synopsys translate_off
defparam \Mux27~15 .lut_mask = 16'hF808;
defparam \Mux27~15 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X63_Y34_N27
dffeas \register[9][4] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\register~94_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~44_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\register[9][4]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \register[9][4] .is_wysiwyg = "true";
defparam \register[9][4] .power_up = "low";
// synopsys translate_on

// Location: FF_X67_Y34_N17
dffeas \register[11][4] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\register~94_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~47_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\register[11][4]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \register[11][4] .is_wysiwyg = "true";
defparam \register[11][4] .power_up = "low";
// synopsys translate_on

// Location: FF_X67_Y38_N15
dffeas \register[8][4] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\register~94_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~46_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\register[8][4]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \register[8][4] .is_wysiwyg = "true";
defparam \register[8][4] .power_up = "low";
// synopsys translate_on

// Location: FF_X67_Y38_N9
dffeas \register[10][4] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\register~94_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~45_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\register[10][4]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \register[10][4] .is_wysiwyg = "true";
defparam \register[10][4] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X67_Y38_N14
cycloneive_lcell_comb \Mux27~12 (
// Equation(s):
// \Mux27~12_combout  = (Selector5 & (Selector41)) # (!Selector5 & ((Selector41 & ((\register[10][4]~q ))) # (!Selector41 & (\register[8][4]~q ))))

	.dataa(Selector5),
	.datab(Selector41),
	.datac(\register[8][4]~q ),
	.datad(\register[10][4]~q ),
	.cin(gnd),
	.combout(\Mux27~12_combout ),
	.cout());
// synopsys translate_off
defparam \Mux27~12 .lut_mask = 16'hDC98;
defparam \Mux27~12 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X67_Y34_N16
cycloneive_lcell_comb \Mux27~13 (
// Equation(s):
// \Mux27~13_combout  = (Selector5 & ((\Mux27~12_combout  & ((\register[11][4]~q ))) # (!\Mux27~12_combout  & (\register[9][4]~q )))) # (!Selector5 & (((\Mux27~12_combout ))))

	.dataa(Selector5),
	.datab(\register[9][4]~q ),
	.datac(\register[11][4]~q ),
	.datad(\Mux27~12_combout ),
	.cin(gnd),
	.combout(\Mux27~13_combout ),
	.cout());
// synopsys translate_off
defparam \Mux27~13 .lut_mask = 16'hF588;
defparam \Mux27~13 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y34_N6
cycloneive_lcell_comb \Mux27~16 (
// Equation(s):
// \Mux27~16_combout  = (Selector2 & (((Selector3) # (\Mux27~13_combout )))) # (!Selector2 & (\Mux27~15_combout  & (!Selector3)))

	.dataa(\Mux27~15_combout ),
	.datab(Selector2),
	.datac(Selector3),
	.datad(\Mux27~13_combout ),
	.cin(gnd),
	.combout(\Mux27~16_combout ),
	.cout());
// synopsys translate_off
defparam \Mux27~16 .lut_mask = 16'hCEC2;
defparam \Mux27~16 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y35_N22
cycloneive_lcell_comb \register~95 (
// Equation(s):
// \register~95_combout  = (WideOr01 & ((\wdat[3]~62_combout ) # ((plif_memwbrtnaddr_l_3 & plif_memwbregsrc_l_1))))

	.dataa(plif_memwbrtnaddr_l_3),
	.datab(wdat_3),
	.datac(WideOr0),
	.datad(plif_memwbregsrc_l_1),
	.cin(gnd),
	.combout(\register~95_combout ),
	.cout());
// synopsys translate_off
defparam \register~95 .lut_mask = 16'hE0C0;
defparam \register~95 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X65_Y34_N17
dffeas \register[20][3] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\register~95_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~35_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\register[20][3]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \register[20][3] .is_wysiwyg = "true";
defparam \register[20][3] .power_up = "low";
// synopsys translate_on

// Location: FF_X65_Y34_N11
dffeas \register[16][3] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\register~95_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~36_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\register[16][3]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \register[16][3] .is_wysiwyg = "true";
defparam \register[16][3] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X66_Y33_N24
cycloneive_lcell_comb \register[24][3]~feeder (
// Equation(s):
// \register[24][3]~feeder_combout  = \register~95_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(\register~95_combout ),
	.datad(gnd),
	.cin(gnd),
	.combout(\register[24][3]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \register[24][3]~feeder .lut_mask = 16'hF0F0;
defparam \register[24][3]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X66_Y33_N25
dffeas \register[24][3] (
	.clk(!CLK),
	.d(\register[24][3]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~34_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\register[24][3]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \register[24][3] .is_wysiwyg = "true";
defparam \register[24][3] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X65_Y34_N10
cycloneive_lcell_comb \Mux28~4 (
// Equation(s):
// \Mux28~4_combout  = (Selector2 & ((Selector3) # ((\register[24][3]~q )))) # (!Selector2 & (!Selector3 & (\register[16][3]~q )))

	.dataa(Selector2),
	.datab(Selector3),
	.datac(\register[16][3]~q ),
	.datad(\register[24][3]~q ),
	.cin(gnd),
	.combout(\Mux28~4_combout ),
	.cout());
// synopsys translate_off
defparam \Mux28~4 .lut_mask = 16'hBA98;
defparam \Mux28~4 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X65_Y34_N8
cycloneive_lcell_comb \Mux28~5 (
// Equation(s):
// \Mux28~5_combout  = (Selector3 & ((\Mux28~4_combout  & (\register[28][3]~q )) # (!\Mux28~4_combout  & ((\register[20][3]~q ))))) # (!Selector3 & (((\Mux28~4_combout ))))

	.dataa(\register[28][3]~q ),
	.datab(\register[20][3]~q ),
	.datac(Selector3),
	.datad(\Mux28~4_combout ),
	.cin(gnd),
	.combout(\Mux28~5_combout ),
	.cout());
// synopsys translate_off
defparam \Mux28~5 .lut_mask = 16'hAFC0;
defparam \Mux28~5 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X67_Y37_N7
dffeas \register[22][3] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\register~95_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~55_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\register[22][3]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \register[22][3] .is_wysiwyg = "true";
defparam \register[22][3] .power_up = "low";
// synopsys translate_on

// Location: FF_X68_Y35_N7
dffeas \register[30][3] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\register~95_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~56_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\register[30][3]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \register[30][3] .is_wysiwyg = "true";
defparam \register[30][3] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X68_Y35_N20
cycloneive_lcell_comb \register[26][3]~feeder (
// Equation(s):
// \register[26][3]~feeder_combout  = \register~95_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(\register~95_combout ),
	.datad(gnd),
	.cin(gnd),
	.combout(\register[26][3]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \register[26][3]~feeder .lut_mask = 16'hF0F0;
defparam \register[26][3]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X68_Y35_N21
dffeas \register[26][3] (
	.clk(!CLK),
	.d(\register[26][3]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~54_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\register[26][3]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \register[26][3] .is_wysiwyg = "true";
defparam \register[26][3] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X67_Y37_N24
cycloneive_lcell_comb \register[18][3]~feeder (
// Equation(s):
// \register[18][3]~feeder_combout  = \register~95_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(\register~95_combout ),
	.datad(gnd),
	.cin(gnd),
	.combout(\register[18][3]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \register[18][3]~feeder .lut_mask = 16'hF0F0;
defparam \register[18][3]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X67_Y37_N25
dffeas \register[18][3] (
	.clk(!CLK),
	.d(\register[18][3]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~33_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\register[18][3]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \register[18][3] .is_wysiwyg = "true";
defparam \register[18][3] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X67_Y37_N26
cycloneive_lcell_comb \Mux28~2 (
// Equation(s):
// \Mux28~2_combout  = (Selector3 & (((Selector2)))) # (!Selector3 & ((Selector2 & (\register[26][3]~q )) # (!Selector2 & ((\register[18][3]~q )))))

	.dataa(Selector3),
	.datab(\register[26][3]~q ),
	.datac(Selector2),
	.datad(\register[18][3]~q ),
	.cin(gnd),
	.combout(\Mux28~2_combout ),
	.cout());
// synopsys translate_off
defparam \Mux28~2 .lut_mask = 16'hE5E0;
defparam \Mux28~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X70_Y37_N16
cycloneive_lcell_comb \Mux28~3 (
// Equation(s):
// \Mux28~3_combout  = (Selector3 & ((\Mux28~2_combout  & ((\register[30][3]~q ))) # (!\Mux28~2_combout  & (\register[22][3]~q )))) # (!Selector3 & (((\Mux28~2_combout ))))

	.dataa(Selector3),
	.datab(\register[22][3]~q ),
	.datac(\register[30][3]~q ),
	.datad(\Mux28~2_combout ),
	.cin(gnd),
	.combout(\Mux28~3_combout ),
	.cout());
// synopsys translate_off
defparam \Mux28~3 .lut_mask = 16'hF588;
defparam \Mux28~3 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X70_Y37_N2
cycloneive_lcell_comb \Mux28~6 (
// Equation(s):
// \Mux28~6_combout  = (Selector41 & (((Selector5) # (\Mux28~3_combout )))) # (!Selector41 & (\Mux28~5_combout  & (!Selector5)))

	.dataa(\Mux28~5_combout ),
	.datab(Selector41),
	.datac(Selector5),
	.datad(\Mux28~3_combout ),
	.cin(gnd),
	.combout(\Mux28~6_combout ),
	.cout());
// synopsys translate_off
defparam \Mux28~6 .lut_mask = 16'hCEC2;
defparam \Mux28~6 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y38_N28
cycloneive_lcell_comb \register[31][3]~feeder (
// Equation(s):
// \register[31][3]~feeder_combout  = \register~95_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(\register~95_combout ),
	.cin(gnd),
	.combout(\register[31][3]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \register[31][3]~feeder .lut_mask = 16'hFF00;
defparam \register[31][3]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X61_Y38_N29
dffeas \register[31][3] (
	.clk(!CLK),
	.d(\register[31][3]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~40_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\register[31][3]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \register[31][3] .is_wysiwyg = "true";
defparam \register[31][3] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X63_Y35_N22
cycloneive_lcell_comb \register[27][3]~feeder (
// Equation(s):
// \register[27][3]~feeder_combout  = \register~95_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(\register~95_combout ),
	.cin(gnd),
	.combout(\register[27][3]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \register[27][3]~feeder .lut_mask = 16'hFF00;
defparam \register[27][3]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X63_Y35_N23
dffeas \register[27][3] (
	.clk(!CLK),
	.d(\register[27][3]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~38_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\register[27][3]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \register[27][3] .is_wysiwyg = "true";
defparam \register[27][3] .power_up = "low";
// synopsys translate_on

// Location: FF_X62_Y31_N5
dffeas \register[23][3] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\register~95_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~37_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\register[23][3]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \register[23][3] .is_wysiwyg = "true";
defparam \register[23][3] .power_up = "low";
// synopsys translate_on

// Location: FF_X62_Y31_N7
dffeas \register[19][3] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\register~95_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~39_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\register[19][3]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \register[19][3] .is_wysiwyg = "true";
defparam \register[19][3] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X62_Y31_N4
cycloneive_lcell_comb \Mux28~7 (
// Equation(s):
// \Mux28~7_combout  = (Selector3 & ((Selector2) # ((\register[23][3]~q )))) # (!Selector3 & (!Selector2 & ((\register[19][3]~q ))))

	.dataa(Selector3),
	.datab(Selector2),
	.datac(\register[23][3]~q ),
	.datad(\register[19][3]~q ),
	.cin(gnd),
	.combout(\Mux28~7_combout ),
	.cout());
// synopsys translate_off
defparam \Mux28~7 .lut_mask = 16'hB9A8;
defparam \Mux28~7 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y38_N30
cycloneive_lcell_comb \Mux28~8 (
// Equation(s):
// \Mux28~8_combout  = (Selector2 & ((\Mux28~7_combout  & (\register[31][3]~q )) # (!\Mux28~7_combout  & ((\register[27][3]~q ))))) # (!Selector2 & (((\Mux28~7_combout ))))

	.dataa(\register[31][3]~q ),
	.datab(Selector2),
	.datac(\register[27][3]~q ),
	.datad(\Mux28~7_combout ),
	.cin(gnd),
	.combout(\Mux28~8_combout ),
	.cout());
// synopsys translate_off
defparam \Mux28~8 .lut_mask = 16'hBBC0;
defparam \Mux28~8 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y36_N8
cycloneive_lcell_comb \register[29][3]~feeder (
// Equation(s):
// \register[29][3]~feeder_combout  = \register~95_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(\register~95_combout ),
	.cin(gnd),
	.combout(\register[29][3]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \register[29][3]~feeder .lut_mask = 16'hFF00;
defparam \register[29][3]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X58_Y36_N9
dffeas \register[29][3] (
	.clk(!CLK),
	.d(\register[29][3]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~28_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\register[29][3]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \register[29][3] .is_wysiwyg = "true";
defparam \register[29][3] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X63_Y31_N14
cycloneive_lcell_comb \register[25][3]~feeder (
// Equation(s):
// \register[25][3]~feeder_combout  = \register~95_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(\register~95_combout ),
	.cin(gnd),
	.combout(\register[25][3]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \register[25][3]~feeder .lut_mask = 16'hFF00;
defparam \register[25][3]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X63_Y31_N15
dffeas \register[25][3] (
	.clk(!CLK),
	.d(\register[25][3]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~24_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\register[25][3]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \register[25][3] .is_wysiwyg = "true";
defparam \register[25][3] .power_up = "low";
// synopsys translate_on

// Location: FF_X62_Y33_N1
dffeas \register[21][3] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\register~95_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~22_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\register[21][3]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \register[21][3] .is_wysiwyg = "true";
defparam \register[21][3] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X60_Y37_N6
cycloneive_lcell_comb \register[17][3]~feeder (
// Equation(s):
// \register[17][3]~feeder_combout  = \register~95_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(\register~95_combout ),
	.cin(gnd),
	.combout(\register[17][3]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \register[17][3]~feeder .lut_mask = 16'hFF00;
defparam \register[17][3]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X60_Y37_N7
dffeas \register[17][3] (
	.clk(!CLK),
	.d(\register[17][3]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~26_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\register[17][3]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \register[17][3] .is_wysiwyg = "true";
defparam \register[17][3] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X62_Y33_N0
cycloneive_lcell_comb \Mux28~0 (
// Equation(s):
// \Mux28~0_combout  = (Selector2 & (Selector3)) # (!Selector2 & ((Selector3 & (\register[21][3]~q )) # (!Selector3 & ((\register[17][3]~q )))))

	.dataa(Selector2),
	.datab(Selector3),
	.datac(\register[21][3]~q ),
	.datad(\register[17][3]~q ),
	.cin(gnd),
	.combout(\Mux28~0_combout ),
	.cout());
// synopsys translate_off
defparam \Mux28~0 .lut_mask = 16'hD9C8;
defparam \Mux28~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X63_Y31_N20
cycloneive_lcell_comb \Mux28~1 (
// Equation(s):
// \Mux28~1_combout  = (Selector2 & ((\Mux28~0_combout  & (\register[29][3]~q )) # (!\Mux28~0_combout  & ((\register[25][3]~q ))))) # (!Selector2 & (((\Mux28~0_combout ))))

	.dataa(\register[29][3]~q ),
	.datab(\register[25][3]~q ),
	.datac(Selector2),
	.datad(\Mux28~0_combout ),
	.cin(gnd),
	.combout(\Mux28~1_combout ),
	.cout());
// synopsys translate_off
defparam \Mux28~1 .lut_mask = 16'hAFC0;
defparam \Mux28~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X61_Y35_N23
dffeas \register[15][3] (
	.clk(!CLK),
	.d(\register~95_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~53_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\register[15][3]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \register[15][3] .is_wysiwyg = "true";
defparam \register[15][3] .power_up = "low";
// synopsys translate_on

// Location: FF_X62_Y33_N19
dffeas \register[14][3] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\register~95_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~61_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\register[14][3]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \register[14][3] .is_wysiwyg = "true";
defparam \register[14][3] .power_up = "low";
// synopsys translate_on

// Location: FF_X60_Y33_N17
dffeas \register[13][3] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\register~95_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~62_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\register[13][3]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \register[13][3] .is_wysiwyg = "true";
defparam \register[13][3] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X60_Y33_N16
cycloneive_lcell_comb \Mux28~17 (
// Equation(s):
// \Mux28~17_combout  = (Selector41 & (((Selector5)))) # (!Selector41 & ((Selector5 & ((\register[13][3]~q ))) # (!Selector5 & (\register[12][3]~q ))))

	.dataa(\register[12][3]~q ),
	.datab(Selector41),
	.datac(\register[13][3]~q ),
	.datad(Selector5),
	.cin(gnd),
	.combout(\Mux28~17_combout ),
	.cout());
// synopsys translate_off
defparam \Mux28~17 .lut_mask = 16'hFC22;
defparam \Mux28~17 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y33_N18
cycloneive_lcell_comb \Mux28~18 (
// Equation(s):
// \Mux28~18_combout  = (Selector41 & ((\Mux28~17_combout  & (\register[15][3]~q )) # (!\Mux28~17_combout  & ((\register[14][3]~q ))))) # (!Selector41 & (((\Mux28~17_combout ))))

	.dataa(Selector41),
	.datab(\register[15][3]~q ),
	.datac(\register[14][3]~q ),
	.datad(\Mux28~17_combout ),
	.cin(gnd),
	.combout(\Mux28~18_combout ),
	.cout());
// synopsys translate_off
defparam \Mux28~18 .lut_mask = 16'hDDA0;
defparam \Mux28~18 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X67_Y34_N29
dffeas \register[2][3] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\register~95_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~50_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\register[2][3]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \register[2][3] .is_wysiwyg = "true";
defparam \register[2][3] .power_up = "low";
// synopsys translate_on

// Location: FF_X70_Y34_N23
dffeas \register[1][3] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\register~95_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~49_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\register[1][3]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \register[1][3] .is_wysiwyg = "true";
defparam \register[1][3] .power_up = "low";
// synopsys translate_on

// Location: FF_X70_Y34_N21
dffeas \register[3][3] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\register~95_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~48_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\register[3][3]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \register[3][3] .is_wysiwyg = "true";
defparam \register[3][3] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X70_Y34_N22
cycloneive_lcell_comb \Mux28~14 (
// Equation(s):
// \Mux28~14_combout  = (Selector4 & ((plif_ifidinstr_l_22 & ((\register[3][3]~q ))) # (!plif_ifidinstr_l_22 & (\register[1][3]~q )))) # (!Selector4 & (((\register[1][3]~q ))))

	.dataa(Selector4),
	.datab(plif_ifidinstr_l_22),
	.datac(\register[1][3]~q ),
	.datad(\register[3][3]~q ),
	.cin(gnd),
	.combout(\Mux28~14_combout ),
	.cout());
// synopsys translate_off
defparam \Mux28~14 .lut_mask = 16'hF870;
defparam \Mux28~14 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X70_Y38_N8
cycloneive_lcell_comb \Mux28~15 (
// Equation(s):
// \Mux28~15_combout  = (Selector5 & (((\Mux28~14_combout )))) # (!Selector5 & (Selector41 & (\register[2][3]~q )))

	.dataa(Selector41),
	.datab(\register[2][3]~q ),
	.datac(Selector5),
	.datad(\Mux28~14_combout ),
	.cin(gnd),
	.combout(\Mux28~15_combout ),
	.cout());
// synopsys translate_off
defparam \Mux28~15 .lut_mask = 16'hF808;
defparam \Mux28~15 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X66_Y31_N9
dffeas \register[6][3] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\register~95_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~58_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\register[6][3]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \register[6][3] .is_wysiwyg = "true";
defparam \register[6][3] .power_up = "low";
// synopsys translate_on

// Location: FF_X66_Y31_N15
dffeas \register[7][3] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\register~95_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~43_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\register[7][3]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \register[7][3] .is_wysiwyg = "true";
defparam \register[7][3] .power_up = "low";
// synopsys translate_on

// Location: FF_X67_Y31_N17
dffeas \register[5][3] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\register~95_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~59_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\register[5][3]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \register[5][3] .is_wysiwyg = "true";
defparam \register[5][3] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X67_Y31_N16
cycloneive_lcell_comb \Mux28~12 (
// Equation(s):
// \Mux28~12_combout  = (Selector41 & (((Selector5)))) # (!Selector41 & ((Selector5 & ((\register[5][3]~q ))) # (!Selector5 & (\register[4][3]~q ))))

	.dataa(\register[4][3]~q ),
	.datab(Selector41),
	.datac(\register[5][3]~q ),
	.datad(Selector5),
	.cin(gnd),
	.combout(\Mux28~12_combout ),
	.cout());
// synopsys translate_off
defparam \Mux28~12 .lut_mask = 16'hFC22;
defparam \Mux28~12 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X66_Y31_N14
cycloneive_lcell_comb \Mux28~13 (
// Equation(s):
// \Mux28~13_combout  = (Selector41 & ((\Mux28~12_combout  & ((\register[7][3]~q ))) # (!\Mux28~12_combout  & (\register[6][3]~q )))) # (!Selector41 & (((\Mux28~12_combout ))))

	.dataa(Selector41),
	.datab(\register[6][3]~q ),
	.datac(\register[7][3]~q ),
	.datad(\Mux28~12_combout ),
	.cin(gnd),
	.combout(\Mux28~13_combout ),
	.cout());
// synopsys translate_off
defparam \Mux28~13 .lut_mask = 16'hF588;
defparam \Mux28~13 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X70_Y38_N22
cycloneive_lcell_comb \Mux28~16 (
// Equation(s):
// \Mux28~16_combout  = (Selector3 & (((Selector2) # (\Mux28~13_combout )))) # (!Selector3 & (\Mux28~15_combout  & (!Selector2)))

	.dataa(Selector3),
	.datab(\Mux28~15_combout ),
	.datac(Selector2),
	.datad(\Mux28~13_combout ),
	.cin(gnd),
	.combout(\Mux28~16_combout ),
	.cout());
// synopsys translate_off
defparam \Mux28~16 .lut_mask = 16'hAEA4;
defparam \Mux28~16 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X70_Y37_N22
cycloneive_lcell_comb \register[9][3]~feeder (
// Equation(s):
// \register[9][3]~feeder_combout  = \register~95_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(\register~95_combout ),
	.datad(gnd),
	.cin(gnd),
	.combout(\register[9][3]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \register[9][3]~feeder .lut_mask = 16'hF0F0;
defparam \register[9][3]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X70_Y37_N23
dffeas \register[9][3] (
	.clk(!CLK),
	.d(\register[9][3]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~44_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\register[9][3]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \register[9][3] .is_wysiwyg = "true";
defparam \register[9][3] .power_up = "low";
// synopsys translate_on

// Location: FF_X67_Y34_N7
dffeas \register[11][3] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\register~95_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~47_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\register[11][3]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \register[11][3] .is_wysiwyg = "true";
defparam \register[11][3] .power_up = "low";
// synopsys translate_on

// Location: FF_X67_Y38_N31
dffeas \register[8][3] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\register~95_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~46_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\register[8][3]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \register[8][3] .is_wysiwyg = "true";
defparam \register[8][3] .power_up = "low";
// synopsys translate_on

// Location: FF_X67_Y38_N25
dffeas \register[10][3] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\register~95_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~45_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\register[10][3]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \register[10][3] .is_wysiwyg = "true";
defparam \register[10][3] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X67_Y38_N30
cycloneive_lcell_comb \Mux28~10 (
// Equation(s):
// \Mux28~10_combout  = (Selector5 & (Selector41)) # (!Selector5 & ((Selector41 & ((\register[10][3]~q ))) # (!Selector41 & (\register[8][3]~q ))))

	.dataa(Selector5),
	.datab(Selector41),
	.datac(\register[8][3]~q ),
	.datad(\register[10][3]~q ),
	.cin(gnd),
	.combout(\Mux28~10_combout ),
	.cout());
// synopsys translate_off
defparam \Mux28~10 .lut_mask = 16'hDC98;
defparam \Mux28~10 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X70_Y37_N0
cycloneive_lcell_comb \Mux28~11 (
// Equation(s):
// \Mux28~11_combout  = (Selector5 & ((\Mux28~10_combout  & ((\register[11][3]~q ))) # (!\Mux28~10_combout  & (\register[9][3]~q )))) # (!Selector5 & (((\Mux28~10_combout ))))

	.dataa(\register[9][3]~q ),
	.datab(\register[11][3]~q ),
	.datac(Selector5),
	.datad(\Mux28~10_combout ),
	.cin(gnd),
	.combout(\Mux28~11_combout ),
	.cout());
// synopsys translate_off
defparam \Mux28~11 .lut_mask = 16'hCFA0;
defparam \Mux28~11 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y31_N16
cycloneive_lcell_comb \Mux61~7 (
// Equation(s):
// \Mux61~7_combout  = (Selector7 & (((Selector8)))) # (!Selector7 & ((Selector8 & ((\register[23][2]~q ))) # (!Selector8 & (\register[19][2]~q ))))

	.dataa(\register[19][2]~q ),
	.datab(Selector7),
	.datac(\register[23][2]~q ),
	.datad(Selector8),
	.cin(gnd),
	.combout(\Mux61~7_combout ),
	.cout());
// synopsys translate_off
defparam \Mux61~7 .lut_mask = 16'hFC22;
defparam \Mux61~7 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y31_N20
cycloneive_lcell_comb \Mux61~8 (
// Equation(s):
// \Mux61~8_combout  = (\Mux61~7_combout  & (((\register[31][2]~q ) # (!Selector7)))) # (!\Mux61~7_combout  & (\register[27][2]~q  & ((Selector7))))

	.dataa(\register[27][2]~q ),
	.datab(\register[31][2]~q ),
	.datac(\Mux61~7_combout ),
	.datad(Selector7),
	.cin(gnd),
	.combout(\Mux61~8_combout ),
	.cout());
// synopsys translate_off
defparam \Mux61~8 .lut_mask = 16'hCAF0;
defparam \Mux61~8 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X60_Y37_N9
dffeas \register[17][2] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\register~91_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~26_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\register[17][2]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \register[17][2] .is_wysiwyg = "true";
defparam \register[17][2] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X60_Y37_N8
cycloneive_lcell_comb \Mux61~0 (
// Equation(s):
// \Mux61~0_combout  = (Selector8 & ((Selector7) # ((\register[21][2]~q )))) # (!Selector8 & (!Selector7 & (\register[17][2]~q )))

	.dataa(Selector8),
	.datab(Selector7),
	.datac(\register[17][2]~q ),
	.datad(\register[21][2]~q ),
	.cin(gnd),
	.combout(\Mux61~0_combout ),
	.cout());
// synopsys translate_off
defparam \Mux61~0 .lut_mask = 16'hBA98;
defparam \Mux61~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X63_Y33_N30
cycloneive_lcell_comb \Mux61~1 (
// Equation(s):
// \Mux61~1_combout  = (Selector7 & ((\Mux61~0_combout  & ((\register[29][2]~q ))) # (!\Mux61~0_combout  & (\register[25][2]~q )))) # (!Selector7 & (((\Mux61~0_combout ))))

	.dataa(\register[25][2]~q ),
	.datab(Selector7),
	.datac(\register[29][2]~q ),
	.datad(\Mux61~0_combout ),
	.cin(gnd),
	.combout(\Mux61~1_combout ),
	.cout());
// synopsys translate_off
defparam \Mux61~1 .lut_mask = 16'hF388;
defparam \Mux61~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X65_Y34_N20
cycloneive_lcell_comb \Mux61~4 (
// Equation(s):
// \Mux61~4_combout  = (Selector7 & ((Selector8) # ((\register[24][2]~q )))) # (!Selector7 & (!Selector8 & (\register[16][2]~q )))

	.dataa(Selector7),
	.datab(Selector8),
	.datac(\register[16][2]~q ),
	.datad(\register[24][2]~q ),
	.cin(gnd),
	.combout(\Mux61~4_combout ),
	.cout());
// synopsys translate_off
defparam \Mux61~4 .lut_mask = 16'hBA98;
defparam \Mux61~4 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X65_Y34_N2
cycloneive_lcell_comb \Mux61~5 (
// Equation(s):
// \Mux61~5_combout  = (\Mux61~4_combout  & (((\register[28][2]~q ) # (!Selector8)))) # (!\Mux61~4_combout  & (\register[20][2]~q  & (Selector8)))

	.dataa(\register[20][2]~q ),
	.datab(\Mux61~4_combout ),
	.datac(Selector8),
	.datad(\register[28][2]~q ),
	.cin(gnd),
	.combout(\Mux61~5_combout ),
	.cout());
// synopsys translate_off
defparam \Mux61~5 .lut_mask = 16'hEC2C;
defparam \Mux61~5 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X68_Y37_N31
dffeas \register[26][2] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\register~91_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~54_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\register[26][2]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \register[26][2] .is_wysiwyg = "true";
defparam \register[26][2] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X68_Y37_N30
cycloneive_lcell_comb \Mux61~2 (
// Equation(s):
// \Mux61~2_combout  = (Selector7 & (((\register[26][2]~q ) # (Selector8)))) # (!Selector7 & (\register[18][2]~q  & ((!Selector8))))

	.dataa(Selector7),
	.datab(\register[18][2]~q ),
	.datac(\register[26][2]~q ),
	.datad(Selector8),
	.cin(gnd),
	.combout(\Mux61~2_combout ),
	.cout());
// synopsys translate_off
defparam \Mux61~2 .lut_mask = 16'hAAE4;
defparam \Mux61~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X69_Y37_N24
cycloneive_lcell_comb \Mux61~3 (
// Equation(s):
// \Mux61~3_combout  = (Selector8 & ((\Mux61~2_combout  & (\register[30][2]~q )) # (!\Mux61~2_combout  & ((\register[22][2]~q ))))) # (!Selector8 & (((\Mux61~2_combout ))))

	.dataa(\register[30][2]~q ),
	.datab(Selector8),
	.datac(\register[22][2]~q ),
	.datad(\Mux61~2_combout ),
	.cin(gnd),
	.combout(\Mux61~3_combout ),
	.cout());
// synopsys translate_off
defparam \Mux61~3 .lut_mask = 16'hBBC0;
defparam \Mux61~3 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X65_Y34_N0
cycloneive_lcell_comb \Mux61~6 (
// Equation(s):
// \Mux61~6_combout  = (Selector91 & (((Selector10) # (\Mux61~3_combout )))) # (!Selector91 & (\Mux61~5_combout  & (!Selector10)))

	.dataa(Selector91),
	.datab(\Mux61~5_combout ),
	.datac(Selector10),
	.datad(\Mux61~3_combout ),
	.cin(gnd),
	.combout(\Mux61~6_combout ),
	.cout());
// synopsys translate_off
defparam \Mux61~6 .lut_mask = 16'hAEA4;
defparam \Mux61~6 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y33_N18
cycloneive_lcell_comb \Mux61~17 (
// Equation(s):
// \Mux61~17_combout  = (Selector10 & ((\register[13][2]~q ) # ((Selector91)))) # (!Selector10 & (((\register[12][2]~q  & !Selector91))))

	.dataa(Selector10),
	.datab(\register[13][2]~q ),
	.datac(\register[12][2]~q ),
	.datad(Selector91),
	.cin(gnd),
	.combout(\Mux61~17_combout ),
	.cout());
// synopsys translate_off
defparam \Mux61~17 .lut_mask = 16'hAAD8;
defparam \Mux61~17 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y35_N14
cycloneive_lcell_comb \Mux61~18 (
// Equation(s):
// \Mux61~18_combout  = (Selector91 & ((\Mux61~17_combout  & ((\register[15][2]~q ))) # (!\Mux61~17_combout  & (\register[14][2]~q )))) # (!Selector91 & (((\Mux61~17_combout ))))

	.dataa(\register[14][2]~q ),
	.datab(Selector91),
	.datac(\Mux61~17_combout ),
	.datad(\register[15][2]~q ),
	.cin(gnd),
	.combout(\Mux61~18_combout ),
	.cout());
// synopsys translate_off
defparam \Mux61~18 .lut_mask = 16'hF838;
defparam \Mux61~18 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X67_Y38_N28
cycloneive_lcell_comb \Mux61~10 (
// Equation(s):
// \Mux61~10_combout  = (Selector91 & (((\register[10][2]~q ) # (Selector10)))) # (!Selector91 & (\register[8][2]~q  & ((!Selector10))))

	.dataa(\register[8][2]~q ),
	.datab(Selector91),
	.datac(\register[10][2]~q ),
	.datad(Selector10),
	.cin(gnd),
	.combout(\Mux61~10_combout ),
	.cout());
// synopsys translate_off
defparam \Mux61~10 .lut_mask = 16'hCCE2;
defparam \Mux61~10 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X66_Y38_N8
cycloneive_lcell_comb \Mux61~11 (
// Equation(s):
// \Mux61~11_combout  = (Selector10 & ((\Mux61~10_combout  & (\register[11][2]~q )) # (!\Mux61~10_combout  & ((\register[9][2]~q ))))) # (!Selector10 & (((\Mux61~10_combout ))))

	.dataa(\register[11][2]~q ),
	.datab(Selector10),
	.datac(\register[9][2]~q ),
	.datad(\Mux61~10_combout ),
	.cin(gnd),
	.combout(\Mux61~11_combout ),
	.cout());
// synopsys translate_off
defparam \Mux61~11 .lut_mask = 16'hBBC0;
defparam \Mux61~11 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X67_Y31_N2
cycloneive_lcell_comb \Mux61~12 (
// Equation(s):
// \Mux61~12_combout  = (Selector10 & ((Selector91) # ((\register[5][2]~q )))) # (!Selector10 & (!Selector91 & (\register[4][2]~q )))

	.dataa(Selector10),
	.datab(Selector91),
	.datac(\register[4][2]~q ),
	.datad(\register[5][2]~q ),
	.cin(gnd),
	.combout(\Mux61~12_combout ),
	.cout());
// synopsys translate_off
defparam \Mux61~12 .lut_mask = 16'hBA98;
defparam \Mux61~12 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X66_Y31_N18
cycloneive_lcell_comb \Mux61~13 (
// Equation(s):
// \Mux61~13_combout  = (Selector91 & ((\Mux61~12_combout  & ((\register[7][2]~q ))) # (!\Mux61~12_combout  & (\register[6][2]~q )))) # (!Selector91 & (((\Mux61~12_combout ))))

	.dataa(Selector91),
	.datab(\register[6][2]~q ),
	.datac(\register[7][2]~q ),
	.datad(\Mux61~12_combout ),
	.cin(gnd),
	.combout(\Mux61~13_combout ),
	.cout());
// synopsys translate_off
defparam \Mux61~13 .lut_mask = 16'hF588;
defparam \Mux61~13 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X68_Y33_N10
cycloneive_lcell_comb \Mux61~15 (
// Equation(s):
// \Mux61~15_combout  = (\Mux61~14_combout ) # ((Selector91 & (\register[2][2]~q  & !Selector10)))

	.dataa(\Mux61~14_combout ),
	.datab(Selector91),
	.datac(\register[2][2]~q ),
	.datad(Selector10),
	.cin(gnd),
	.combout(\Mux61~15_combout ),
	.cout());
// synopsys translate_off
defparam \Mux61~15 .lut_mask = 16'hAAEA;
defparam \Mux61~15 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y35_N0
cycloneive_lcell_comb \Mux61~16 (
// Equation(s):
// \Mux61~16_combout  = (Selector7 & (Selector8)) # (!Selector7 & ((Selector8 & (\Mux61~13_combout )) # (!Selector8 & ((\Mux61~15_combout )))))

	.dataa(Selector7),
	.datab(Selector8),
	.datac(\Mux61~13_combout ),
	.datad(\Mux61~15_combout ),
	.cin(gnd),
	.combout(\Mux61~16_combout ),
	.cout());
// synopsys translate_off
defparam \Mux61~16 .lut_mask = 16'hD9C8;
defparam \Mux61~16 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y39_N30
cycloneive_lcell_comb \Mux23~7 (
// Equation(s):
// \Mux23~7_combout  = (Selector3 & (((Selector2)))) # (!Selector3 & ((Selector2 & ((\register[27][8]~q ))) # (!Selector2 & (\register[19][8]~q ))))

	.dataa(Selector3),
	.datab(\register[19][8]~q ),
	.datac(\register[27][8]~q ),
	.datad(Selector2),
	.cin(gnd),
	.combout(\Mux23~7_combout ),
	.cout());
// synopsys translate_off
defparam \Mux23~7 .lut_mask = 16'hFA44;
defparam \Mux23~7 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y38_N12
cycloneive_lcell_comb \Mux23~8 (
// Equation(s):
// \Mux23~8_combout  = (\Mux23~7_combout  & (((\register[31][8]~q )) # (!Selector3))) # (!\Mux23~7_combout  & (Selector3 & (\register[23][8]~q )))

	.dataa(\Mux23~7_combout ),
	.datab(Selector3),
	.datac(\register[23][8]~q ),
	.datad(\register[31][8]~q ),
	.cin(gnd),
	.combout(\Mux23~8_combout ),
	.cout());
// synopsys translate_off
defparam \Mux23~8 .lut_mask = 16'hEA62;
defparam \Mux23~8 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X70_Y39_N28
cycloneive_lcell_comb \Mux23~4 (
// Equation(s):
// \Mux23~4_combout  = (Selector3 & ((\register[20][8]~q ) # ((Selector2)))) # (!Selector3 & (((!Selector2 & \register[16][8]~q ))))

	.dataa(\register[20][8]~q ),
	.datab(Selector3),
	.datac(Selector2),
	.datad(\register[16][8]~q ),
	.cin(gnd),
	.combout(\Mux23~4_combout ),
	.cout());
// synopsys translate_off
defparam \Mux23~4 .lut_mask = 16'hCBC8;
defparam \Mux23~4 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X68_Y36_N6
cycloneive_lcell_comb \Mux23~5 (
// Equation(s):
// \Mux23~5_combout  = (Selector2 & ((\Mux23~4_combout  & ((\register[28][8]~q ))) # (!\Mux23~4_combout  & (\register[24][8]~q )))) # (!Selector2 & (((\Mux23~4_combout ))))

	.dataa(Selector2),
	.datab(\register[24][8]~q ),
	.datac(\register[28][8]~q ),
	.datad(\Mux23~4_combout ),
	.cin(gnd),
	.combout(\Mux23~5_combout ),
	.cout());
// synopsys translate_off
defparam \Mux23~5 .lut_mask = 16'hF588;
defparam \Mux23~5 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X69_Y37_N28
cycloneive_lcell_comb \register[18][8]~feeder (
// Equation(s):
// \register[18][8]~feeder_combout  = \register~87_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(\register~87_combout ),
	.cin(gnd),
	.combout(\register[18][8]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \register[18][8]~feeder .lut_mask = 16'hFF00;
defparam \register[18][8]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X69_Y37_N29
dffeas \register[18][8] (
	.clk(!CLK),
	.d(\register[18][8]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~33_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\register[18][8]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \register[18][8] .is_wysiwyg = "true";
defparam \register[18][8] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X69_Y37_N18
cycloneive_lcell_comb \Mux23~2 (
// Equation(s):
// \Mux23~2_combout  = (Selector2 & (((Selector3)))) # (!Selector2 & ((Selector3 & (\register[22][8]~q )) # (!Selector3 & ((\register[18][8]~q )))))

	.dataa(\register[22][8]~q ),
	.datab(\register[18][8]~q ),
	.datac(Selector2),
	.datad(Selector3),
	.cin(gnd),
	.combout(\Mux23~2_combout ),
	.cout());
// synopsys translate_off
defparam \Mux23~2 .lut_mask = 16'hFA0C;
defparam \Mux23~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X69_Y37_N8
cycloneive_lcell_comb \Mux23~3 (
// Equation(s):
// \Mux23~3_combout  = (\Mux23~2_combout  & (((\register[30][8]~q ) # (!Selector2)))) # (!\Mux23~2_combout  & (\register[26][8]~q  & (Selector2)))

	.dataa(\register[26][8]~q ),
	.datab(\Mux23~2_combout ),
	.datac(Selector2),
	.datad(\register[30][8]~q ),
	.cin(gnd),
	.combout(\Mux23~3_combout ),
	.cout());
// synopsys translate_off
defparam \Mux23~3 .lut_mask = 16'hEC2C;
defparam \Mux23~3 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X68_Y36_N4
cycloneive_lcell_comb \Mux23~6 (
// Equation(s):
// \Mux23~6_combout  = (Selector5 & (((Selector41)))) # (!Selector5 & ((Selector41 & ((\Mux23~3_combout ))) # (!Selector41 & (\Mux23~5_combout ))))

	.dataa(\Mux23~5_combout ),
	.datab(Selector5),
	.datac(Selector41),
	.datad(\Mux23~3_combout ),
	.cin(gnd),
	.combout(\Mux23~6_combout ),
	.cout());
// synopsys translate_off
defparam \Mux23~6 .lut_mask = 16'hF2C2;
defparam \Mux23~6 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y35_N0
cycloneive_lcell_comb \Mux23~0 (
// Equation(s):
// \Mux23~0_combout  = (Selector3 & (((Selector2)))) # (!Selector3 & ((Selector2 & (\register[25][8]~q )) # (!Selector2 & ((\register[17][8]~q )))))

	.dataa(\register[25][8]~q ),
	.datab(Selector3),
	.datac(\register[17][8]~q ),
	.datad(Selector2),
	.cin(gnd),
	.combout(\Mux23~0_combout ),
	.cout());
// synopsys translate_off
defparam \Mux23~0 .lut_mask = 16'hEE30;
defparam \Mux23~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X63_Y33_N6
cycloneive_lcell_comb \Mux23~1 (
// Equation(s):
// \Mux23~1_combout  = (Selector3 & ((\Mux23~0_combout  & ((\register[29][8]~q ))) # (!\Mux23~0_combout  & (\register[21][8]~q )))) # (!Selector3 & (((\Mux23~0_combout ))))

	.dataa(Selector3),
	.datab(\register[21][8]~q ),
	.datac(\register[29][8]~q ),
	.datad(\Mux23~0_combout ),
	.cin(gnd),
	.combout(\Mux23~1_combout ),
	.cout());
// synopsys translate_off
defparam \Mux23~1 .lut_mask = 16'hF588;
defparam \Mux23~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X60_Y33_N11
dffeas \register[12][8] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\register~87_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~52_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\register[12][8]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \register[12][8] .is_wysiwyg = "true";
defparam \register[12][8] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X60_Y33_N10
cycloneive_lcell_comb \Mux23~17 (
// Equation(s):
// \Mux23~17_combout  = (Selector5 & ((\register[13][8]~q ) # ((Selector41)))) # (!Selector5 & (((\register[12][8]~q  & !Selector41))))

	.dataa(Selector5),
	.datab(\register[13][8]~q ),
	.datac(\register[12][8]~q ),
	.datad(Selector41),
	.cin(gnd),
	.combout(\Mux23~17_combout ),
	.cout());
// synopsys translate_off
defparam \Mux23~17 .lut_mask = 16'hAAD8;
defparam \Mux23~17 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X68_Y36_N12
cycloneive_lcell_comb \Mux23~18 (
// Equation(s):
// \Mux23~18_combout  = (Selector41 & ((\Mux23~17_combout  & ((\register[15][8]~q ))) # (!\Mux23~17_combout  & (\register[14][8]~q )))) # (!Selector41 & (((\Mux23~17_combout ))))

	.dataa(Selector41),
	.datab(\register[14][8]~q ),
	.datac(\register[15][8]~q ),
	.datad(\Mux23~17_combout ),
	.cin(gnd),
	.combout(\Mux23~18_combout ),
	.cout());
// synopsys translate_off
defparam \Mux23~18 .lut_mask = 16'hF588;
defparam \Mux23~18 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X68_Y33_N4
cycloneive_lcell_comb \register[7][8]~feeder (
// Equation(s):
// \register[7][8]~feeder_combout  = \register~87_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(\register~87_combout ),
	.datad(gnd),
	.cin(gnd),
	.combout(\register[7][8]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \register[7][8]~feeder .lut_mask = 16'hF0F0;
defparam \register[7][8]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X68_Y33_N5
dffeas \register[7][8] (
	.clk(!CLK),
	.d(\register[7][8]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~43_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\register[7][8]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \register[7][8] .is_wysiwyg = "true";
defparam \register[7][8] .power_up = "low";
// synopsys translate_on

// Location: FF_X67_Y31_N23
dffeas \register[4][8] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\register~87_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~60_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\register[4][8]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \register[4][8] .is_wysiwyg = "true";
defparam \register[4][8] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X67_Y31_N22
cycloneive_lcell_comb \Mux23~10 (
// Equation(s):
// \Mux23~10_combout  = (Selector41 & (((Selector5)))) # (!Selector41 & ((Selector5 & (\register[5][8]~q )) # (!Selector5 & ((\register[4][8]~q )))))

	.dataa(Selector41),
	.datab(\register[5][8]~q ),
	.datac(\register[4][8]~q ),
	.datad(Selector5),
	.cin(gnd),
	.combout(\Mux23~10_combout ),
	.cout());
// synopsys translate_off
defparam \Mux23~10 .lut_mask = 16'hEE50;
defparam \Mux23~10 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X68_Y33_N14
cycloneive_lcell_comb \Mux23~11 (
// Equation(s):
// \Mux23~11_combout  = (Selector41 & ((\Mux23~10_combout  & ((\register[7][8]~q ))) # (!\Mux23~10_combout  & (\register[6][8]~q )))) # (!Selector41 & (((\Mux23~10_combout ))))

	.dataa(\register[6][8]~q ),
	.datab(\register[7][8]~q ),
	.datac(Selector41),
	.datad(\Mux23~10_combout ),
	.cin(gnd),
	.combout(\Mux23~11_combout ),
	.cout());
// synopsys translate_off
defparam \Mux23~11 .lut_mask = 16'hCFA0;
defparam \Mux23~11 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X70_Y34_N10
cycloneive_lcell_comb \Mux23~14 (
// Equation(s):
// \Mux23~14_combout  = (Selector4 & ((plif_ifidinstr_l_22 & ((\register[3][8]~q ))) # (!plif_ifidinstr_l_22 & (\register[1][8]~q )))) # (!Selector4 & (((\register[1][8]~q ))))

	.dataa(Selector4),
	.datab(plif_ifidinstr_l_22),
	.datac(\register[1][8]~q ),
	.datad(\register[3][8]~q ),
	.cin(gnd),
	.combout(\Mux23~14_combout ),
	.cout());
// synopsys translate_off
defparam \Mux23~14 .lut_mask = 16'hF870;
defparam \Mux23~14 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X68_Y36_N0
cycloneive_lcell_comb \Mux23~15 (
// Equation(s):
// \Mux23~15_combout  = (Selector5 & (((\Mux23~14_combout )))) # (!Selector5 & (\register[2][8]~q  & (Selector41)))

	.dataa(\register[2][8]~q ),
	.datab(Selector5),
	.datac(Selector41),
	.datad(\Mux23~14_combout ),
	.cin(gnd),
	.combout(\Mux23~15_combout ),
	.cout());
// synopsys translate_off
defparam \Mux23~15 .lut_mask = 16'hEC20;
defparam \Mux23~15 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X67_Y38_N7
dffeas \register[8][8] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\register~87_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~46_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\register[8][8]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \register[8][8] .is_wysiwyg = "true";
defparam \register[8][8] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X67_Y38_N6
cycloneive_lcell_comb \Mux23~12 (
// Equation(s):
// \Mux23~12_combout  = (Selector5 & (((Selector41)))) # (!Selector5 & ((Selector41 & (\register[10][8]~q )) # (!Selector41 & ((\register[8][8]~q )))))

	.dataa(Selector5),
	.datab(\register[10][8]~q ),
	.datac(\register[8][8]~q ),
	.datad(Selector41),
	.cin(gnd),
	.combout(\Mux23~12_combout ),
	.cout());
// synopsys translate_off
defparam \Mux23~12 .lut_mask = 16'hEE50;
defparam \Mux23~12 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X66_Y38_N2
cycloneive_lcell_comb \Mux23~13 (
// Equation(s):
// \Mux23~13_combout  = (Selector5 & ((\Mux23~12_combout  & ((\register[11][8]~q ))) # (!\Mux23~12_combout  & (\register[9][8]~q )))) # (!Selector5 & (((\Mux23~12_combout ))))

	.dataa(Selector5),
	.datab(\register[9][8]~q ),
	.datac(\register[11][8]~q ),
	.datad(\Mux23~12_combout ),
	.cin(gnd),
	.combout(\Mux23~13_combout ),
	.cout());
// synopsys translate_off
defparam \Mux23~13 .lut_mask = 16'hF588;
defparam \Mux23~13 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X68_Y36_N18
cycloneive_lcell_comb \Mux23~16 (
// Equation(s):
// \Mux23~16_combout  = (Selector3 & (((Selector2)))) # (!Selector3 & ((Selector2 & ((\Mux23~13_combout ))) # (!Selector2 & (\Mux23~15_combout ))))

	.dataa(\Mux23~15_combout ),
	.datab(Selector3),
	.datac(Selector2),
	.datad(\Mux23~13_combout ),
	.cin(gnd),
	.combout(\Mux23~16_combout ),
	.cout());
// synopsys translate_off
defparam \Mux23~16 .lut_mask = 16'hF2C2;
defparam \Mux23~16 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y31_N12
cycloneive_lcell_comb \Mux24~7 (
// Equation(s):
// \Mux24~7_combout  = (Selector3 & (((\register[23][7]~q ) # (Selector2)))) # (!Selector3 & (\register[19][7]~q  & ((!Selector2))))

	.dataa(Selector3),
	.datab(\register[19][7]~q ),
	.datac(\register[23][7]~q ),
	.datad(Selector2),
	.cin(gnd),
	.combout(\Mux24~7_combout ),
	.cout());
// synopsys translate_off
defparam \Mux24~7 .lut_mask = 16'hAAE4;
defparam \Mux24~7 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y31_N0
cycloneive_lcell_comb \Mux24~8 (
// Equation(s):
// \Mux24~8_combout  = (Selector2 & ((\Mux24~7_combout  & (\register[31][7]~q )) # (!\Mux24~7_combout  & ((\register[27][7]~q ))))) # (!Selector2 & (((\Mux24~7_combout ))))

	.dataa(\register[31][7]~q ),
	.datab(Selector2),
	.datac(\Mux24~7_combout ),
	.datad(\register[27][7]~q ),
	.cin(gnd),
	.combout(\Mux24~8_combout ),
	.cout());
// synopsys translate_off
defparam \Mux24~8 .lut_mask = 16'hBCB0;
defparam \Mux24~8 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y35_N10
cycloneive_lcell_comb \Mux24~0 (
// Equation(s):
// \Mux24~0_combout  = (Selector3 & ((\register[21][7]~q ) # ((Selector2)))) # (!Selector3 & (((\register[17][7]~q  & !Selector2))))

	.dataa(\register[21][7]~q ),
	.datab(Selector3),
	.datac(\register[17][7]~q ),
	.datad(Selector2),
	.cin(gnd),
	.combout(\Mux24~0_combout ),
	.cout());
// synopsys translate_off
defparam \Mux24~0 .lut_mask = 16'hCCB8;
defparam \Mux24~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y31_N26
cycloneive_lcell_comb \Mux24~1 (
// Equation(s):
// \Mux24~1_combout  = (Selector2 & ((\Mux24~0_combout  & (\register[29][7]~q )) # (!\Mux24~0_combout  & ((\register[25][7]~q ))))) # (!Selector2 & (((\Mux24~0_combout ))))

	.dataa(\register[29][7]~q ),
	.datab(Selector2),
	.datac(\register[25][7]~q ),
	.datad(\Mux24~0_combout ),
	.cin(gnd),
	.combout(\Mux24~1_combout ),
	.cout());
// synopsys translate_off
defparam \Mux24~1 .lut_mask = 16'hBBC0;
defparam \Mux24~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X68_Y38_N18
cycloneive_lcell_comb \Mux24~2 (
// Equation(s):
// \Mux24~2_combout  = (Selector3 & (((Selector2)))) # (!Selector3 & ((Selector2 & ((\register[26][7]~q ))) # (!Selector2 & (\register[18][7]~q ))))

	.dataa(Selector3),
	.datab(\register[18][7]~q ),
	.datac(\register[26][7]~q ),
	.datad(Selector2),
	.cin(gnd),
	.combout(\Mux24~2_combout ),
	.cout());
// synopsys translate_off
defparam \Mux24~2 .lut_mask = 16'hFA44;
defparam \Mux24~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X67_Y37_N0
cycloneive_lcell_comb \Mux24~3 (
// Equation(s):
// \Mux24~3_combout  = (Selector3 & ((\Mux24~2_combout  & (\register[30][7]~q )) # (!\Mux24~2_combout  & ((\register[22][7]~q ))))) # (!Selector3 & (((\Mux24~2_combout ))))

	.dataa(Selector3),
	.datab(\register[30][7]~q ),
	.datac(\register[22][7]~q ),
	.datad(\Mux24~2_combout ),
	.cin(gnd),
	.combout(\Mux24~3_combout ),
	.cout());
// synopsys translate_off
defparam \Mux24~3 .lut_mask = 16'hDDA0;
defparam \Mux24~3 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X69_Y38_N7
dffeas \register[20][7] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\register~88_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~35_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\register[20][7]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \register[20][7] .is_wysiwyg = "true";
defparam \register[20][7] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X69_Y38_N6
cycloneive_lcell_comb \Mux24~5 (
// Equation(s):
// \Mux24~5_combout  = (\Mux24~4_combout  & ((\register[28][7]~q ) # ((!Selector3)))) # (!\Mux24~4_combout  & (((\register[20][7]~q  & Selector3))))

	.dataa(\Mux24~4_combout ),
	.datab(\register[28][7]~q ),
	.datac(\register[20][7]~q ),
	.datad(Selector3),
	.cin(gnd),
	.combout(\Mux24~5_combout ),
	.cout());
// synopsys translate_off
defparam \Mux24~5 .lut_mask = 16'hD8AA;
defparam \Mux24~5 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y40_N18
cycloneive_lcell_comb \Mux24~6 (
// Equation(s):
// \Mux24~6_combout  = (Selector5 & (Selector41)) # (!Selector5 & ((Selector41 & (\Mux24~3_combout )) # (!Selector41 & ((\Mux24~5_combout )))))

	.dataa(Selector5),
	.datab(Selector41),
	.datac(\Mux24~3_combout ),
	.datad(\Mux24~5_combout ),
	.cin(gnd),
	.combout(\Mux24~6_combout ),
	.cout());
// synopsys translate_off
defparam \Mux24~6 .lut_mask = 16'hD9C8;
defparam \Mux24~6 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X63_Y30_N6
cycloneive_lcell_comb \Mux24~17 (
// Equation(s):
// \Mux24~17_combout  = (Selector5 & ((\register[13][7]~q ) # ((Selector41)))) # (!Selector5 & (((\register[12][7]~q  & !Selector41))))

	.dataa(Selector5),
	.datab(\register[13][7]~q ),
	.datac(\register[12][7]~q ),
	.datad(Selector41),
	.cin(gnd),
	.combout(\Mux24~17_combout ),
	.cout());
// synopsys translate_off
defparam \Mux24~17 .lut_mask = 16'hAAD8;
defparam \Mux24~17 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X66_Y33_N28
cycloneive_lcell_comb \Mux24~18 (
// Equation(s):
// \Mux24~18_combout  = (Selector41 & ((\Mux24~17_combout  & (\register[15][7]~q )) # (!\Mux24~17_combout  & ((\register[14][7]~q ))))) # (!Selector41 & (((\Mux24~17_combout ))))

	.dataa(Selector41),
	.datab(\register[15][7]~q ),
	.datac(\Mux24~17_combout ),
	.datad(\register[14][7]~q ),
	.cin(gnd),
	.combout(\Mux24~18_combout ),
	.cout());
// synopsys translate_off
defparam \Mux24~18 .lut_mask = 16'hDAD0;
defparam \Mux24~18 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X67_Y38_N21
dffeas \register[10][7] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\register~88_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~45_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\register[10][7]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \register[10][7] .is_wysiwyg = "true";
defparam \register[10][7] .power_up = "low";
// synopsys translate_on

// Location: FF_X67_Y38_N11
dffeas \register[8][7] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\register~88_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~46_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\register[8][7]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \register[8][7] .is_wysiwyg = "true";
defparam \register[8][7] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X67_Y38_N10
cycloneive_lcell_comb \Mux24~10 (
// Equation(s):
// \Mux24~10_combout  = (Selector5 & (((Selector41)))) # (!Selector5 & ((Selector41 & (\register[10][7]~q )) # (!Selector41 & ((\register[8][7]~q )))))

	.dataa(Selector5),
	.datab(\register[10][7]~q ),
	.datac(\register[8][7]~q ),
	.datad(Selector41),
	.cin(gnd),
	.combout(\Mux24~10_combout ),
	.cout());
// synopsys translate_off
defparam \Mux24~10 .lut_mask = 16'hEE50;
defparam \Mux24~10 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X66_Y38_N16
cycloneive_lcell_comb \Mux24~11 (
// Equation(s):
// \Mux24~11_combout  = (\Mux24~10_combout  & ((\register[11][7]~q ) # ((!Selector5)))) # (!\Mux24~10_combout  & (((\register[9][7]~q  & Selector5))))

	.dataa(\register[11][7]~q ),
	.datab(\Mux24~10_combout ),
	.datac(\register[9][7]~q ),
	.datad(Selector5),
	.cin(gnd),
	.combout(\Mux24~11_combout ),
	.cout());
// synopsys translate_off
defparam \Mux24~11 .lut_mask = 16'hB8CC;
defparam \Mux24~11 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X67_Y31_N14
cycloneive_lcell_comb \Mux24~12 (
// Equation(s):
// \Mux24~12_combout  = (Selector41 & (((Selector5)))) # (!Selector41 & ((Selector5 & (\register[5][7]~q )) # (!Selector5 & ((\register[4][7]~q )))))

	.dataa(Selector41),
	.datab(\register[5][7]~q ),
	.datac(\register[4][7]~q ),
	.datad(Selector5),
	.cin(gnd),
	.combout(\Mux24~12_combout ),
	.cout());
// synopsys translate_off
defparam \Mux24~12 .lut_mask = 16'hEE50;
defparam \Mux24~12 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X68_Y32_N10
cycloneive_lcell_comb \Mux24~13 (
// Equation(s):
// \Mux24~13_combout  = (Selector41 & ((\Mux24~12_combout  & ((\register[7][7]~q ))) # (!\Mux24~12_combout  & (\register[6][7]~q )))) # (!Selector41 & (((\Mux24~12_combout ))))

	.dataa(Selector41),
	.datab(\register[6][7]~q ),
	.datac(\register[7][7]~q ),
	.datad(\Mux24~12_combout ),
	.cin(gnd),
	.combout(\Mux24~13_combout ),
	.cout());
// synopsys translate_off
defparam \Mux24~13 .lut_mask = 16'hF588;
defparam \Mux24~13 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X70_Y33_N16
cycloneive_lcell_comb \Mux24~14 (
// Equation(s):
// \Mux24~14_combout  = (Selector5 & ((Selector41 & ((\register[3][7]~q ))) # (!Selector41 & (\register[1][7]~q ))))

	.dataa(\register[1][7]~q ),
	.datab(Selector41),
	.datac(Selector5),
	.datad(\register[3][7]~q ),
	.cin(gnd),
	.combout(\Mux24~14_combout ),
	.cout());
// synopsys translate_off
defparam \Mux24~14 .lut_mask = 16'hE020;
defparam \Mux24~14 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y40_N6
cycloneive_lcell_comb \Mux24~15 (
// Equation(s):
// \Mux24~15_combout  = (\Mux24~14_combout ) # ((!Selector5 & (Selector41 & \register[2][7]~q )))

	.dataa(Selector5),
	.datab(Selector41),
	.datac(\Mux24~14_combout ),
	.datad(\register[2][7]~q ),
	.cin(gnd),
	.combout(\Mux24~15_combout ),
	.cout());
// synopsys translate_off
defparam \Mux24~15 .lut_mask = 16'hF4F0;
defparam \Mux24~15 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y40_N0
cycloneive_lcell_comb \Mux24~16 (
// Equation(s):
// \Mux24~16_combout  = (Selector3 & ((Selector2) # ((\Mux24~13_combout )))) # (!Selector3 & (!Selector2 & ((\Mux24~15_combout ))))

	.dataa(Selector3),
	.datab(Selector2),
	.datac(\Mux24~13_combout ),
	.datad(\Mux24~15_combout ),
	.cin(gnd),
	.combout(\Mux24~16_combout ),
	.cout());
// synopsys translate_off
defparam \Mux24~16 .lut_mask = 16'hB9A8;
defparam \Mux24~16 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y39_N26
cycloneive_lcell_comb \Mux25~7 (
// Equation(s):
// \Mux25~7_combout  = (Selector3 & (((Selector2)))) # (!Selector3 & ((Selector2 & ((\register[27][6]~q ))) # (!Selector2 & (\register[19][6]~q ))))

	.dataa(Selector3),
	.datab(\register[19][6]~q ),
	.datac(\register[27][6]~q ),
	.datad(Selector2),
	.cin(gnd),
	.combout(\Mux25~7_combout ),
	.cout());
// synopsys translate_off
defparam \Mux25~7 .lut_mask = 16'hFA44;
defparam \Mux25~7 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y38_N4
cycloneive_lcell_comb \Mux25~8 (
// Equation(s):
// \Mux25~8_combout  = (\Mux25~7_combout  & (((\register[31][6]~q )) # (!Selector3))) # (!\Mux25~7_combout  & (Selector3 & (\register[23][6]~q )))

	.dataa(\Mux25~7_combout ),
	.datab(Selector3),
	.datac(\register[23][6]~q ),
	.datad(\register[31][6]~q ),
	.cin(gnd),
	.combout(\Mux25~8_combout ),
	.cout());
// synopsys translate_off
defparam \Mux25~8 .lut_mask = 16'hEA62;
defparam \Mux25~8 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X68_Y37_N23
dffeas \register[26][6] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\register~89_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~54_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\register[26][6]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \register[26][6] .is_wysiwyg = "true";
defparam \register[26][6] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X68_Y38_N14
cycloneive_lcell_comb \Mux25~3 (
// Equation(s):
// \Mux25~3_combout  = (\Mux25~2_combout  & ((\register[30][6]~q ) # ((!Selector2)))) # (!\Mux25~2_combout  & (((\register[26][6]~q  & Selector2))))

	.dataa(\Mux25~2_combout ),
	.datab(\register[30][6]~q ),
	.datac(\register[26][6]~q ),
	.datad(Selector2),
	.cin(gnd),
	.combout(\Mux25~3_combout ),
	.cout());
// synopsys translate_off
defparam \Mux25~3 .lut_mask = 16'hD8AA;
defparam \Mux25~3 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X65_Y37_N20
cycloneive_lcell_comb \register[16][6]~feeder (
// Equation(s):
// \register[16][6]~feeder_combout  = \register~89_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(\register~89_combout ),
	.datad(gnd),
	.cin(gnd),
	.combout(\register[16][6]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \register[16][6]~feeder .lut_mask = 16'hF0F0;
defparam \register[16][6]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X65_Y37_N21
dffeas \register[16][6] (
	.clk(!CLK),
	.d(\register[16][6]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~36_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\register[16][6]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \register[16][6] .is_wysiwyg = "true";
defparam \register[16][6] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X65_Y37_N26
cycloneive_lcell_comb \Mux25~4 (
// Equation(s):
// \Mux25~4_combout  = (Selector3 & ((Selector2) # ((\register[20][6]~q )))) # (!Selector3 & (!Selector2 & ((\register[16][6]~q ))))

	.dataa(Selector3),
	.datab(Selector2),
	.datac(\register[20][6]~q ),
	.datad(\register[16][6]~q ),
	.cin(gnd),
	.combout(\Mux25~4_combout ),
	.cout());
// synopsys translate_off
defparam \Mux25~4 .lut_mask = 16'hB9A8;
defparam \Mux25~4 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X65_Y38_N30
cycloneive_lcell_comb \Mux25~5 (
// Equation(s):
// \Mux25~5_combout  = (\Mux25~4_combout  & (((\register[28][6]~q ) # (!Selector2)))) # (!\Mux25~4_combout  & (\register[24][6]~q  & ((Selector2))))

	.dataa(\register[24][6]~q ),
	.datab(\Mux25~4_combout ),
	.datac(\register[28][6]~q ),
	.datad(Selector2),
	.cin(gnd),
	.combout(\Mux25~5_combout ),
	.cout());
// synopsys translate_off
defparam \Mux25~5 .lut_mask = 16'hE2CC;
defparam \Mux25~5 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X67_Y36_N24
cycloneive_lcell_comb \Mux25~6 (
// Equation(s):
// \Mux25~6_combout  = (Selector41 & ((\Mux25~3_combout ) # ((Selector5)))) # (!Selector41 & (((!Selector5 & \Mux25~5_combout ))))

	.dataa(Selector41),
	.datab(\Mux25~3_combout ),
	.datac(Selector5),
	.datad(\Mux25~5_combout ),
	.cin(gnd),
	.combout(\Mux25~6_combout ),
	.cout());
// synopsys translate_off
defparam \Mux25~6 .lut_mask = 16'hADA8;
defparam \Mux25~6 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X62_Y34_N5
dffeas \register[17][6] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\register~89_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~26_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\register[17][6]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \register[17][6] .is_wysiwyg = "true";
defparam \register[17][6] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X62_Y34_N4
cycloneive_lcell_comb \Mux25~0 (
// Equation(s):
// \Mux25~0_combout  = (Selector3 & (((Selector2)))) # (!Selector3 & ((Selector2 & (\register[25][6]~q )) # (!Selector2 & ((\register[17][6]~q )))))

	.dataa(\register[25][6]~q ),
	.datab(Selector3),
	.datac(\register[17][6]~q ),
	.datad(Selector2),
	.cin(gnd),
	.combout(\Mux25~0_combout ),
	.cout());
// synopsys translate_off
defparam \Mux25~0 .lut_mask = 16'hEE30;
defparam \Mux25~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X63_Y33_N16
cycloneive_lcell_comb \Mux25~1 (
// Equation(s):
// \Mux25~1_combout  = (Selector3 & ((\Mux25~0_combout  & ((\register[29][6]~q ))) # (!\Mux25~0_combout  & (\register[21][6]~q )))) # (!Selector3 & (((\Mux25~0_combout ))))

	.dataa(Selector3),
	.datab(\register[21][6]~q ),
	.datac(\register[29][6]~q ),
	.datad(\Mux25~0_combout ),
	.cin(gnd),
	.combout(\Mux25~1_combout ),
	.cout());
// synopsys translate_off
defparam \Mux25~1 .lut_mask = 16'hF588;
defparam \Mux25~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X63_Y30_N18
cycloneive_lcell_comb \Mux25~17 (
// Equation(s):
// \Mux25~17_combout  = (Selector41 & (((Selector5)))) # (!Selector41 & ((Selector5 & (\register[13][6]~q )) # (!Selector5 & ((\register[12][6]~q )))))

	.dataa(\register[13][6]~q ),
	.datab(Selector41),
	.datac(\register[12][6]~q ),
	.datad(Selector5),
	.cin(gnd),
	.combout(\Mux25~17_combout ),
	.cout());
// synopsys translate_off
defparam \Mux25~17 .lut_mask = 16'hEE30;
defparam \Mux25~17 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X66_Y33_N2
cycloneive_lcell_comb \Mux25~18 (
// Equation(s):
// \Mux25~18_combout  = (Selector41 & ((\Mux25~17_combout  & ((\register[15][6]~q ))) # (!\Mux25~17_combout  & (\register[14][6]~q )))) # (!Selector41 & (((\Mux25~17_combout ))))

	.dataa(\register[14][6]~q ),
	.datab(\register[15][6]~q ),
	.datac(Selector41),
	.datad(\Mux25~17_combout ),
	.cin(gnd),
	.combout(\Mux25~18_combout ),
	.cout());
// synopsys translate_off
defparam \Mux25~18 .lut_mask = 16'hCFA0;
defparam \Mux25~18 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X67_Y31_N13
dffeas \register[5][6] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\register~89_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~59_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\register[5][6]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \register[5][6] .is_wysiwyg = "true";
defparam \register[5][6] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X67_Y31_N12
cycloneive_lcell_comb \Mux25~10 (
// Equation(s):
// \Mux25~10_combout  = (Selector5 & (((\register[5][6]~q ) # (Selector41)))) # (!Selector5 & (\register[4][6]~q  & ((!Selector41))))

	.dataa(\register[4][6]~q ),
	.datab(Selector5),
	.datac(\register[5][6]~q ),
	.datad(Selector41),
	.cin(gnd),
	.combout(\Mux25~10_combout ),
	.cout());
// synopsys translate_off
defparam \Mux25~10 .lut_mask = 16'hCCE2;
defparam \Mux25~10 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X66_Y31_N3
dffeas \register[6][6] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\register~89_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~58_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\register[6][6]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \register[6][6] .is_wysiwyg = "true";
defparam \register[6][6] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X66_Y31_N2
cycloneive_lcell_comb \Mux25~11 (
// Equation(s):
// \Mux25~11_combout  = (\Mux25~10_combout  & ((\register[7][6]~q ) # ((!Selector41)))) # (!\Mux25~10_combout  & (((\register[6][6]~q  & Selector41))))

	.dataa(\Mux25~10_combout ),
	.datab(\register[7][6]~q ),
	.datac(\register[6][6]~q ),
	.datad(Selector41),
	.cin(gnd),
	.combout(\Mux25~11_combout ),
	.cout());
// synopsys translate_off
defparam \Mux25~11 .lut_mask = 16'hD8AA;
defparam \Mux25~11 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X70_Y33_N6
cycloneive_lcell_comb \Mux25~14 (
// Equation(s):
// \Mux25~14_combout  = (Selector5 & ((Selector41 & (\register[3][6]~q )) # (!Selector41 & ((\register[1][6]~q )))))

	.dataa(Selector5),
	.datab(\register[3][6]~q ),
	.datac(Selector41),
	.datad(\register[1][6]~q ),
	.cin(gnd),
	.combout(\Mux25~14_combout ),
	.cout());
// synopsys translate_off
defparam \Mux25~14 .lut_mask = 16'h8A80;
defparam \Mux25~14 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X67_Y36_N8
cycloneive_lcell_comb \Mux25~15 (
// Equation(s):
// \Mux25~15_combout  = (\Mux25~14_combout ) # ((!Selector5 & (\register[2][6]~q  & Selector41)))

	.dataa(Selector5),
	.datab(\register[2][6]~q ),
	.datac(\Mux25~14_combout ),
	.datad(Selector41),
	.cin(gnd),
	.combout(\Mux25~15_combout ),
	.cout());
// synopsys translate_off
defparam \Mux25~15 .lut_mask = 16'hF4F0;
defparam \Mux25~15 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X67_Y38_N18
cycloneive_lcell_comb \Mux25~12 (
// Equation(s):
// \Mux25~12_combout  = (Selector5 & (Selector41)) # (!Selector5 & ((Selector41 & ((\register[10][6]~q ))) # (!Selector41 & (\register[8][6]~q ))))

	.dataa(Selector5),
	.datab(Selector41),
	.datac(\register[8][6]~q ),
	.datad(\register[10][6]~q ),
	.cin(gnd),
	.combout(\Mux25~12_combout ),
	.cout());
// synopsys translate_off
defparam \Mux25~12 .lut_mask = 16'hDC98;
defparam \Mux25~12 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X66_Y34_N24
cycloneive_lcell_comb \Mux25~13 (
// Equation(s):
// \Mux25~13_combout  = (Selector5 & ((\Mux25~12_combout  & ((\register[11][6]~q ))) # (!\Mux25~12_combout  & (\register[9][6]~q )))) # (!Selector5 & (((\Mux25~12_combout ))))

	.dataa(Selector5),
	.datab(\register[9][6]~q ),
	.datac(\register[11][6]~q ),
	.datad(\Mux25~12_combout ),
	.cin(gnd),
	.combout(\Mux25~13_combout ),
	.cout());
// synopsys translate_off
defparam \Mux25~13 .lut_mask = 16'hF588;
defparam \Mux25~13 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X67_Y36_N10
cycloneive_lcell_comb \Mux25~16 (
// Equation(s):
// \Mux25~16_combout  = (Selector2 & (((Selector3) # (\Mux25~13_combout )))) # (!Selector2 & (\Mux25~15_combout  & (!Selector3)))

	.dataa(\Mux25~15_combout ),
	.datab(Selector2),
	.datac(Selector3),
	.datad(\Mux25~13_combout ),
	.cin(gnd),
	.combout(\Mux25~16_combout ),
	.cout());
// synopsys translate_off
defparam \Mux25~16 .lut_mask = 16'hCEC2;
defparam \Mux25~16 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y31_N8
cycloneive_lcell_comb \Mux26~7 (
// Equation(s):
// \Mux26~7_combout  = (Selector3 & ((Selector2) # ((\register[23][5]~q )))) # (!Selector3 & (!Selector2 & ((\register[19][5]~q ))))

	.dataa(Selector3),
	.datab(Selector2),
	.datac(\register[23][5]~q ),
	.datad(\register[19][5]~q ),
	.cin(gnd),
	.combout(\Mux26~7_combout ),
	.cout());
// synopsys translate_off
defparam \Mux26~7 .lut_mask = 16'hB9A8;
defparam \Mux26~7 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X63_Y31_N2
cycloneive_lcell_comb \Mux26~8 (
// Equation(s):
// \Mux26~8_combout  = (Selector2 & ((\Mux26~7_combout  & ((\register[31][5]~q ))) # (!\Mux26~7_combout  & (\register[27][5]~q )))) # (!Selector2 & (((\Mux26~7_combout ))))

	.dataa(Selector2),
	.datab(\register[27][5]~q ),
	.datac(\register[31][5]~q ),
	.datad(\Mux26~7_combout ),
	.cin(gnd),
	.combout(\Mux26~8_combout ),
	.cout());
// synopsys translate_off
defparam \Mux26~8 .lut_mask = 16'hF588;
defparam \Mux26~8 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X68_Y38_N30
cycloneive_lcell_comb \Mux26~2 (
// Equation(s):
// \Mux26~2_combout  = (Selector3 & (((Selector2)))) # (!Selector3 & ((Selector2 & ((\register[26][5]~q ))) # (!Selector2 & (\register[18][5]~q ))))

	.dataa(Selector3),
	.datab(\register[18][5]~q ),
	.datac(\register[26][5]~q ),
	.datad(Selector2),
	.cin(gnd),
	.combout(\Mux26~2_combout ),
	.cout());
// synopsys translate_off
defparam \Mux26~2 .lut_mask = 16'hFA44;
defparam \Mux26~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X69_Y37_N10
cycloneive_lcell_comb \Mux26~3 (
// Equation(s):
// \Mux26~3_combout  = (Selector3 & ((\Mux26~2_combout  & (\register[30][5]~q )) # (!\Mux26~2_combout  & ((\register[22][5]~q ))))) # (!Selector3 & (((\Mux26~2_combout ))))

	.dataa(Selector3),
	.datab(\register[30][5]~q ),
	.datac(\register[22][5]~q ),
	.datad(\Mux26~2_combout ),
	.cin(gnd),
	.combout(\Mux26~3_combout ),
	.cout());
// synopsys translate_off
defparam \Mux26~3 .lut_mask = 16'hDDA0;
defparam \Mux26~3 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X70_Y38_N2
cycloneive_lcell_comb \Mux26~4 (
// Equation(s):
// \Mux26~4_combout  = (Selector2 & (((\register[24][5]~q ) # (Selector3)))) # (!Selector2 & (\register[16][5]~q  & ((!Selector3))))

	.dataa(\register[16][5]~q ),
	.datab(\register[24][5]~q ),
	.datac(Selector2),
	.datad(Selector3),
	.cin(gnd),
	.combout(\Mux26~4_combout ),
	.cout());
// synopsys translate_off
defparam \Mux26~4 .lut_mask = 16'hF0CA;
defparam \Mux26~4 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X70_Y38_N24
cycloneive_lcell_comb \Mux26~5 (
// Equation(s):
// \Mux26~5_combout  = (Selector3 & ((\Mux26~4_combout  & (\register[28][5]~q )) # (!\Mux26~4_combout  & ((\register[20][5]~q ))))) # (!Selector3 & (((\Mux26~4_combout ))))

	.dataa(\register[28][5]~q ),
	.datab(\register[20][5]~q ),
	.datac(Selector3),
	.datad(\Mux26~4_combout ),
	.cin(gnd),
	.combout(\Mux26~5_combout ),
	.cout());
// synopsys translate_off
defparam \Mux26~5 .lut_mask = 16'hAFC0;
defparam \Mux26~5 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X70_Y38_N26
cycloneive_lcell_comb \Mux26~6 (
// Equation(s):
// \Mux26~6_combout  = (Selector5 & (Selector41)) # (!Selector5 & ((Selector41 & (\Mux26~3_combout )) # (!Selector41 & ((\Mux26~5_combout )))))

	.dataa(Selector5),
	.datab(Selector41),
	.datac(\Mux26~3_combout ),
	.datad(\Mux26~5_combout ),
	.cin(gnd),
	.combout(\Mux26~6_combout ),
	.cout());
// synopsys translate_off
defparam \Mux26~6 .lut_mask = 16'hD9C8;
defparam \Mux26~6 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y35_N18
cycloneive_lcell_comb \Mux26~0 (
// Equation(s):
// \Mux26~0_combout  = (Selector2 & (Selector3)) # (!Selector2 & ((Selector3 & ((\register[21][5]~q ))) # (!Selector3 & (\register[17][5]~q ))))

	.dataa(Selector2),
	.datab(Selector3),
	.datac(\register[17][5]~q ),
	.datad(\register[21][5]~q ),
	.cin(gnd),
	.combout(\Mux26~0_combout ),
	.cout());
// synopsys translate_off
defparam \Mux26~0 .lut_mask = 16'hDC98;
defparam \Mux26~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y38_N16
cycloneive_lcell_comb \Mux26~1 (
// Equation(s):
// \Mux26~1_combout  = (\Mux26~0_combout  & (((\register[29][5]~q )) # (!Selector2))) # (!\Mux26~0_combout  & (Selector2 & (\register[25][5]~q )))

	.dataa(\Mux26~0_combout ),
	.datab(Selector2),
	.datac(\register[25][5]~q ),
	.datad(\register[29][5]~q ),
	.cin(gnd),
	.combout(\Mux26~1_combout ),
	.cout());
// synopsys translate_off
defparam \Mux26~1 .lut_mask = 16'hEA62;
defparam \Mux26~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X69_Y32_N0
cycloneive_lcell_comb \Mux26~12 (
// Equation(s):
// \Mux26~12_combout  = (Selector5 & (((\register[5][5]~q ) # (Selector41)))) # (!Selector5 & (\register[4][5]~q  & ((!Selector41))))

	.dataa(\register[4][5]~q ),
	.datab(Selector5),
	.datac(\register[5][5]~q ),
	.datad(Selector41),
	.cin(gnd),
	.combout(\Mux26~12_combout ),
	.cout());
// synopsys translate_off
defparam \Mux26~12 .lut_mask = 16'hCCE2;
defparam \Mux26~12 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X66_Y31_N30
cycloneive_lcell_comb \Mux26~13 (
// Equation(s):
// \Mux26~13_combout  = (Selector41 & ((\Mux26~12_combout  & ((\register[7][5]~q ))) # (!\Mux26~12_combout  & (\register[6][5]~q )))) # (!Selector41 & (((\Mux26~12_combout ))))

	.dataa(Selector41),
	.datab(\register[6][5]~q ),
	.datac(\register[7][5]~q ),
	.datad(\Mux26~12_combout ),
	.cin(gnd),
	.combout(\Mux26~13_combout ),
	.cout());
// synopsys translate_off
defparam \Mux26~13 .lut_mask = 16'hF588;
defparam \Mux26~13 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X70_Y34_N28
cycloneive_lcell_comb \Mux26~14 (
// Equation(s):
// \Mux26~14_combout  = (plif_ifidinstr_l_22 & ((Selector4 & ((\register[3][5]~q ))) # (!Selector4 & (\register[1][5]~q )))) # (!plif_ifidinstr_l_22 & (\register[1][5]~q ))

	.dataa(\register[1][5]~q ),
	.datab(plif_ifidinstr_l_22),
	.datac(\register[3][5]~q ),
	.datad(Selector4),
	.cin(gnd),
	.combout(\Mux26~14_combout ),
	.cout());
// synopsys translate_off
defparam \Mux26~14 .lut_mask = 16'hE2AA;
defparam \Mux26~14 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X66_Y34_N0
cycloneive_lcell_comb \Mux26~15 (
// Equation(s):
// \Mux26~15_combout  = (Selector5 & (((\Mux26~14_combout )))) # (!Selector5 & (Selector41 & (\register[2][5]~q )))

	.dataa(Selector41),
	.datab(Selector5),
	.datac(\register[2][5]~q ),
	.datad(\Mux26~14_combout ),
	.cin(gnd),
	.combout(\Mux26~15_combout ),
	.cout());
// synopsys translate_off
defparam \Mux26~15 .lut_mask = 16'hEC20;
defparam \Mux26~15 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X67_Y36_N6
cycloneive_lcell_comb \Mux26~16 (
// Equation(s):
// \Mux26~16_combout  = (Selector3 & ((\Mux26~13_combout ) # ((Selector2)))) # (!Selector3 & (((\Mux26~15_combout  & !Selector2))))

	.dataa(\Mux26~13_combout ),
	.datab(Selector3),
	.datac(\Mux26~15_combout ),
	.datad(Selector2),
	.cin(gnd),
	.combout(\Mux26~16_combout ),
	.cout());
// synopsys translate_off
defparam \Mux26~16 .lut_mask = 16'hCCB8;
defparam \Mux26~16 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X63_Y30_N14
cycloneive_lcell_comb \Mux26~17 (
// Equation(s):
// \Mux26~17_combout  = (Selector5 & ((Selector41) # ((\register[13][5]~q )))) # (!Selector5 & (!Selector41 & (\register[12][5]~q )))

	.dataa(Selector5),
	.datab(Selector41),
	.datac(\register[12][5]~q ),
	.datad(\register[13][5]~q ),
	.cin(gnd),
	.combout(\Mux26~17_combout ),
	.cout());
// synopsys translate_off
defparam \Mux26~17 .lut_mask = 16'hBA98;
defparam \Mux26~17 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X67_Y33_N26
cycloneive_lcell_comb \Mux26~18 (
// Equation(s):
// \Mux26~18_combout  = (Selector41 & ((\Mux26~17_combout  & ((\register[15][5]~q ))) # (!\Mux26~17_combout  & (\register[14][5]~q )))) # (!Selector41 & (((\Mux26~17_combout ))))

	.dataa(Selector41),
	.datab(\register[14][5]~q ),
	.datac(\Mux26~17_combout ),
	.datad(\register[15][5]~q ),
	.cin(gnd),
	.combout(\Mux26~18_combout ),
	.cout());
// synopsys translate_off
defparam \Mux26~18 .lut_mask = 16'hF858;
defparam \Mux26~18 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X62_Y40_N9
dffeas \register[10][5] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\register~90_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~45_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\register[10][5]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \register[10][5] .is_wysiwyg = "true";
defparam \register[10][5] .power_up = "low";
// synopsys translate_on

// Location: FF_X62_Y40_N31
dffeas \register[8][5] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\register~90_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~46_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\register[8][5]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \register[8][5] .is_wysiwyg = "true";
defparam \register[8][5] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X62_Y40_N30
cycloneive_lcell_comb \Mux26~10 (
// Equation(s):
// \Mux26~10_combout  = (Selector41 & ((\register[10][5]~q ) # ((Selector5)))) # (!Selector41 & (((\register[8][5]~q  & !Selector5))))

	.dataa(Selector41),
	.datab(\register[10][5]~q ),
	.datac(\register[8][5]~q ),
	.datad(Selector5),
	.cin(gnd),
	.combout(\Mux26~10_combout ),
	.cout());
// synopsys translate_off
defparam \Mux26~10 .lut_mask = 16'hAAD8;
defparam \Mux26~10 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X66_Y38_N20
cycloneive_lcell_comb \Mux26~11 (
// Equation(s):
// \Mux26~11_combout  = (Selector5 & ((\Mux26~10_combout  & (\register[11][5]~q )) # (!\Mux26~10_combout  & ((\register[9][5]~q ))))) # (!Selector5 & (((\Mux26~10_combout ))))

	.dataa(Selector5),
	.datab(\register[11][5]~q ),
	.datac(\register[9][5]~q ),
	.datad(\Mux26~10_combout ),
	.cin(gnd),
	.combout(\Mux26~11_combout ),
	.cout());
// synopsys translate_off
defparam \Mux26~11 .lut_mask = 16'hDDA0;
defparam \Mux26~11 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y31_N6
cycloneive_lcell_comb \Mux60~7 (
// Equation(s):
// \Mux60~7_combout  = (Selector8 & (Selector7)) # (!Selector8 & ((Selector7 & ((\register[27][3]~q ))) # (!Selector7 & (\register[19][3]~q ))))

	.dataa(Selector8),
	.datab(Selector7),
	.datac(\register[19][3]~q ),
	.datad(\register[27][3]~q ),
	.cin(gnd),
	.combout(\Mux60~7_combout ),
	.cout());
// synopsys translate_off
defparam \Mux60~7 .lut_mask = 16'hDC98;
defparam \Mux60~7 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y36_N30
cycloneive_lcell_comb \Mux60~8 (
// Equation(s):
// \Mux60~8_combout  = (\Mux60~7_combout  & (((\register[31][3]~q )) # (!Selector8))) # (!\Mux60~7_combout  & (Selector8 & ((\register[23][3]~q ))))

	.dataa(\Mux60~7_combout ),
	.datab(Selector8),
	.datac(\register[31][3]~q ),
	.datad(\register[23][3]~q ),
	.cin(gnd),
	.combout(\Mux60~8_combout ),
	.cout());
// synopsys translate_off
defparam \Mux60~8 .lut_mask = 16'hE6A2;
defparam \Mux60~8 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y37_N4
cycloneive_lcell_comb \Mux60~0 (
// Equation(s):
// \Mux60~0_combout  = (Selector8 & (Selector7)) # (!Selector8 & ((Selector7 & (\register[25][3]~q )) # (!Selector7 & ((\register[17][3]~q )))))

	.dataa(Selector8),
	.datab(Selector7),
	.datac(\register[25][3]~q ),
	.datad(\register[17][3]~q ),
	.cin(gnd),
	.combout(\Mux60~0_combout ),
	.cout());
// synopsys translate_off
defparam \Mux60~0 .lut_mask = 16'hD9C8;
defparam \Mux60~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y36_N22
cycloneive_lcell_comb \Mux60~1 (
// Equation(s):
// \Mux60~1_combout  = (Selector8 & ((\Mux60~0_combout  & ((\register[29][3]~q ))) # (!\Mux60~0_combout  & (\register[21][3]~q )))) # (!Selector8 & (((\Mux60~0_combout ))))

	.dataa(\register[21][3]~q ),
	.datab(Selector8),
	.datac(\register[29][3]~q ),
	.datad(\Mux60~0_combout ),
	.cin(gnd),
	.combout(\Mux60~1_combout ),
	.cout());
// synopsys translate_off
defparam \Mux60~1 .lut_mask = 16'hF388;
defparam \Mux60~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X65_Y34_N16
cycloneive_lcell_comb \Mux60~4 (
// Equation(s):
// \Mux60~4_combout  = (Selector7 & (Selector8)) # (!Selector7 & ((Selector8 & (\register[20][3]~q )) # (!Selector8 & ((\register[16][3]~q )))))

	.dataa(Selector7),
	.datab(Selector8),
	.datac(\register[20][3]~q ),
	.datad(\register[16][3]~q ),
	.cin(gnd),
	.combout(\Mux60~4_combout ),
	.cout());
// synopsys translate_off
defparam \Mux60~4 .lut_mask = 16'hD9C8;
defparam \Mux60~4 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X66_Y33_N10
cycloneive_lcell_comb \register[28][3]~feeder (
// Equation(s):
// \register[28][3]~feeder_combout  = \register~95_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(\register~95_combout ),
	.datad(gnd),
	.cin(gnd),
	.combout(\register[28][3]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \register[28][3]~feeder .lut_mask = 16'hF0F0;
defparam \register[28][3]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X66_Y33_N11
dffeas \register[28][3] (
	.clk(!CLK),
	.d(\register[28][3]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~57_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\register[28][3]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \register[28][3] .is_wysiwyg = "true";
defparam \register[28][3] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X66_Y33_N12
cycloneive_lcell_comb \Mux60~5 (
// Equation(s):
// \Mux60~5_combout  = (Selector7 & ((\Mux60~4_combout  & ((\register[28][3]~q ))) # (!\Mux60~4_combout  & (\register[24][3]~q )))) # (!Selector7 & (((\Mux60~4_combout ))))

	.dataa(Selector7),
	.datab(\register[24][3]~q ),
	.datac(\Mux60~4_combout ),
	.datad(\register[28][3]~q ),
	.cin(gnd),
	.combout(\Mux60~5_combout ),
	.cout());
// synopsys translate_off
defparam \Mux60~5 .lut_mask = 16'hF858;
defparam \Mux60~5 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X67_Y37_N6
cycloneive_lcell_comb \Mux60~2 (
// Equation(s):
// \Mux60~2_combout  = (Selector8 & (((\register[22][3]~q ) # (Selector7)))) # (!Selector8 & (\register[18][3]~q  & ((!Selector7))))

	.dataa(Selector8),
	.datab(\register[18][3]~q ),
	.datac(\register[22][3]~q ),
	.datad(Selector7),
	.cin(gnd),
	.combout(\Mux60~2_combout ),
	.cout());
// synopsys translate_off
defparam \Mux60~2 .lut_mask = 16'hAAE4;
defparam \Mux60~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X68_Y35_N6
cycloneive_lcell_comb \Mux60~3 (
// Equation(s):
// \Mux60~3_combout  = (Selector7 & ((\Mux60~2_combout  & ((\register[30][3]~q ))) # (!\Mux60~2_combout  & (\register[26][3]~q )))) # (!Selector7 & (((\Mux60~2_combout ))))

	.dataa(Selector7),
	.datab(\register[26][3]~q ),
	.datac(\register[30][3]~q ),
	.datad(\Mux60~2_combout ),
	.cin(gnd),
	.combout(\Mux60~3_combout ),
	.cout());
// synopsys translate_off
defparam \Mux60~3 .lut_mask = 16'hF588;
defparam \Mux60~3 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y36_N16
cycloneive_lcell_comb \Mux60~6 (
// Equation(s):
// \Mux60~6_combout  = (Selector91 & (((\Mux60~3_combout ) # (Selector10)))) # (!Selector91 & (\Mux60~5_combout  & ((!Selector10))))

	.dataa(\Mux60~5_combout ),
	.datab(Selector91),
	.datac(\Mux60~3_combout ),
	.datad(Selector10),
	.cin(gnd),
	.combout(\Mux60~6_combout ),
	.cout());
// synopsys translate_off
defparam \Mux60~6 .lut_mask = 16'hCCE2;
defparam \Mux60~6 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X67_Y31_N7
dffeas \register[4][3] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\register~95_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~60_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\register[4][3]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \register[4][3] .is_wysiwyg = "true";
defparam \register[4][3] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X67_Y31_N6
cycloneive_lcell_comb \Mux60~10 (
// Equation(s):
// \Mux60~10_combout  = (Selector10 & ((\register[5][3]~q ) # ((Selector91)))) # (!Selector10 & (((\register[4][3]~q  & !Selector91))))

	.dataa(Selector10),
	.datab(\register[5][3]~q ),
	.datac(\register[4][3]~q ),
	.datad(Selector91),
	.cin(gnd),
	.combout(\Mux60~10_combout ),
	.cout());
// synopsys translate_off
defparam \Mux60~10 .lut_mask = 16'hAAD8;
defparam \Mux60~10 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X66_Y31_N8
cycloneive_lcell_comb \Mux60~11 (
// Equation(s):
// \Mux60~11_combout  = (Selector91 & ((\Mux60~10_combout  & (\register[7][3]~q )) # (!\Mux60~10_combout  & ((\register[6][3]~q ))))) # (!Selector91 & (((\Mux60~10_combout ))))

	.dataa(Selector91),
	.datab(\register[7][3]~q ),
	.datac(\register[6][3]~q ),
	.datad(\Mux60~10_combout ),
	.cin(gnd),
	.combout(\Mux60~11_combout ),
	.cout());
// synopsys translate_off
defparam \Mux60~11 .lut_mask = 16'hDDA0;
defparam \Mux60~11 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X60_Y33_N27
dffeas \register[12][3] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\register~95_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~52_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\register[12][3]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \register[12][3] .is_wysiwyg = "true";
defparam \register[12][3] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X60_Y33_N26
cycloneive_lcell_comb \Mux60~17 (
// Equation(s):
// \Mux60~17_combout  = (Selector10 & ((\register[13][3]~q ) # ((Selector91)))) # (!Selector10 & (((\register[12][3]~q  & !Selector91))))

	.dataa(Selector10),
	.datab(\register[13][3]~q ),
	.datac(\register[12][3]~q ),
	.datad(Selector91),
	.cin(gnd),
	.combout(\Mux60~17_combout ),
	.cout());
// synopsys translate_off
defparam \Mux60~17 .lut_mask = 16'hAAD8;
defparam \Mux60~17 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y36_N14
cycloneive_lcell_comb \Mux60~18 (
// Equation(s):
// \Mux60~18_combout  = (\Mux60~17_combout  & (((\register[15][3]~q )) # (!Selector91))) # (!\Mux60~17_combout  & (Selector91 & ((\register[14][3]~q ))))

	.dataa(\Mux60~17_combout ),
	.datab(Selector91),
	.datac(\register[15][3]~q ),
	.datad(\register[14][3]~q ),
	.cin(gnd),
	.combout(\Mux60~18_combout ),
	.cout());
// synopsys translate_off
defparam \Mux60~18 .lut_mask = 16'hE6A2;
defparam \Mux60~18 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X67_Y34_N28
cycloneive_lcell_comb \Mux60~15 (
// Equation(s):
// \Mux60~15_combout  = (\Mux60~14_combout ) # ((!Selector10 & (\register[2][3]~q  & Selector91)))

	.dataa(\Mux60~14_combout ),
	.datab(Selector10),
	.datac(\register[2][3]~q ),
	.datad(Selector91),
	.cin(gnd),
	.combout(\Mux60~15_combout ),
	.cout());
// synopsys translate_off
defparam \Mux60~15 .lut_mask = 16'hBAAA;
defparam \Mux60~15 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X67_Y38_N24
cycloneive_lcell_comb \Mux60~12 (
// Equation(s):
// \Mux60~12_combout  = (Selector91 & (((\register[10][3]~q ) # (Selector10)))) # (!Selector91 & (\register[8][3]~q  & ((!Selector10))))

	.dataa(\register[8][3]~q ),
	.datab(Selector91),
	.datac(\register[10][3]~q ),
	.datad(Selector10),
	.cin(gnd),
	.combout(\Mux60~12_combout ),
	.cout());
// synopsys translate_off
defparam \Mux60~12 .lut_mask = 16'hCCE2;
defparam \Mux60~12 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X67_Y34_N6
cycloneive_lcell_comb \Mux60~13 (
// Equation(s):
// \Mux60~13_combout  = (Selector10 & ((\Mux60~12_combout  & ((\register[11][3]~q ))) # (!\Mux60~12_combout  & (\register[9][3]~q )))) # (!Selector10 & (((\Mux60~12_combout ))))

	.dataa(\register[9][3]~q ),
	.datab(Selector10),
	.datac(\register[11][3]~q ),
	.datad(\Mux60~12_combout ),
	.cin(gnd),
	.combout(\Mux60~13_combout ),
	.cout());
// synopsys translate_off
defparam \Mux60~13 .lut_mask = 16'hF388;
defparam \Mux60~13 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X67_Y34_N10
cycloneive_lcell_comb \Mux60~16 (
// Equation(s):
// \Mux60~16_combout  = (Selector8 & (((Selector7)))) # (!Selector8 & ((Selector7 & ((\Mux60~13_combout ))) # (!Selector7 & (\Mux60~15_combout ))))

	.dataa(Selector8),
	.datab(\Mux60~15_combout ),
	.datac(Selector7),
	.datad(\Mux60~13_combout ),
	.cin(gnd),
	.combout(\Mux60~16_combout ),
	.cout());
// synopsys translate_off
defparam \Mux60~16 .lut_mask = 16'hF4A4;
defparam \Mux60~16 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X68_Y37_N29
dffeas \register[26][16] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\register~79_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~54_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\register[26][16]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \register[26][16] .is_wysiwyg = "true";
defparam \register[26][16] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X67_Y37_N20
cycloneive_lcell_comb \Mux15~2 (
// Equation(s):
// \Mux15~2_combout  = (Selector2 & (((Selector3)))) # (!Selector2 & ((Selector3 & ((\register[22][16]~q ))) # (!Selector3 & (\register[18][16]~q ))))

	.dataa(\register[18][16]~q ),
	.datab(Selector2),
	.datac(\register[22][16]~q ),
	.datad(Selector3),
	.cin(gnd),
	.combout(\Mux15~2_combout ),
	.cout());
// synopsys translate_off
defparam \Mux15~2 .lut_mask = 16'hFC22;
defparam \Mux15~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X68_Y37_N28
cycloneive_lcell_comb \Mux15~3 (
// Equation(s):
// \Mux15~3_combout  = (Selector2 & ((\Mux15~2_combout  & (\register[30][16]~q )) # (!\Mux15~2_combout  & ((\register[26][16]~q ))))) # (!Selector2 & (((\Mux15~2_combout ))))

	.dataa(Selector2),
	.datab(\register[30][16]~q ),
	.datac(\register[26][16]~q ),
	.datad(\Mux15~2_combout ),
	.cin(gnd),
	.combout(\Mux15~3_combout ),
	.cout());
// synopsys translate_off
defparam \Mux15~3 .lut_mask = 16'hDDA0;
defparam \Mux15~3 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X68_Y34_N0
cycloneive_lcell_comb \Mux15~5 (
// Equation(s):
// \Mux15~5_combout  = (\Mux15~4_combout  & (((\register[28][16]~q )) # (!Selector2))) # (!\Mux15~4_combout  & (Selector2 & ((\register[24][16]~q ))))

	.dataa(\Mux15~4_combout ),
	.datab(Selector2),
	.datac(\register[28][16]~q ),
	.datad(\register[24][16]~q ),
	.cin(gnd),
	.combout(\Mux15~5_combout ),
	.cout());
// synopsys translate_off
defparam \Mux15~5 .lut_mask = 16'hE6A2;
defparam \Mux15~5 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X63_Y36_N30
cycloneive_lcell_comb \Mux15~6 (
// Equation(s):
// \Mux15~6_combout  = (Selector41 & ((Selector5) # ((\Mux15~3_combout )))) # (!Selector41 & (!Selector5 & ((\Mux15~5_combout ))))

	.dataa(Selector41),
	.datab(Selector5),
	.datac(\Mux15~3_combout ),
	.datad(\Mux15~5_combout ),
	.cin(gnd),
	.combout(\Mux15~6_combout ),
	.cout());
// synopsys translate_off
defparam \Mux15~6 .lut_mask = 16'hB9A8;
defparam \Mux15~6 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X62_Y31_N27
dffeas \register[19][16] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\register~79_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~39_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\register[19][16]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \register[19][16] .is_wysiwyg = "true";
defparam \register[19][16] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X62_Y31_N26
cycloneive_lcell_comb \Mux15~7 (
// Equation(s):
// \Mux15~7_combout  = (Selector3 & (Selector2)) # (!Selector3 & ((Selector2 & ((\register[27][16]~q ))) # (!Selector2 & (\register[19][16]~q ))))

	.dataa(Selector3),
	.datab(Selector2),
	.datac(\register[19][16]~q ),
	.datad(\register[27][16]~q ),
	.cin(gnd),
	.combout(\Mux15~7_combout ),
	.cout());
// synopsys translate_off
defparam \Mux15~7 .lut_mask = 16'hDC98;
defparam \Mux15~7 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X63_Y36_N4
cycloneive_lcell_comb \Mux15~8 (
// Equation(s):
// \Mux15~8_combout  = (\Mux15~7_combout  & (((\register[31][16]~q )) # (!Selector3))) # (!\Mux15~7_combout  & (Selector3 & ((\register[23][16]~q ))))

	.dataa(\Mux15~7_combout ),
	.datab(Selector3),
	.datac(\register[31][16]~q ),
	.datad(\register[23][16]~q ),
	.cin(gnd),
	.combout(\Mux15~8_combout ),
	.cout());
// synopsys translate_off
defparam \Mux15~8 .lut_mask = 16'hE6A2;
defparam \Mux15~8 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X63_Y35_N1
dffeas \register[21][16] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\register~79_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~22_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\register[21][16]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \register[21][16] .is_wysiwyg = "true";
defparam \register[21][16] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X61_Y37_N26
cycloneive_lcell_comb \Mux15~0 (
// Equation(s):
// \Mux15~0_combout  = (Selector2 & ((Selector3) # ((\register[25][16]~q )))) # (!Selector2 & (!Selector3 & ((\register[17][16]~q ))))

	.dataa(Selector2),
	.datab(Selector3),
	.datac(\register[25][16]~q ),
	.datad(\register[17][16]~q ),
	.cin(gnd),
	.combout(\Mux15~0_combout ),
	.cout());
// synopsys translate_off
defparam \Mux15~0 .lut_mask = 16'hB9A8;
defparam \Mux15~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X63_Y35_N0
cycloneive_lcell_comb \Mux15~1 (
// Equation(s):
// \Mux15~1_combout  = (Selector3 & ((\Mux15~0_combout  & (\register[29][16]~q )) # (!\Mux15~0_combout  & ((\register[21][16]~q ))))) # (!Selector3 & (((\Mux15~0_combout ))))

	.dataa(\register[29][16]~q ),
	.datab(Selector3),
	.datac(\register[21][16]~q ),
	.datad(\Mux15~0_combout ),
	.cin(gnd),
	.combout(\Mux15~1_combout ),
	.cout());
// synopsys translate_off
defparam \Mux15~1 .lut_mask = 16'hBBC0;
defparam \Mux15~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X69_Y32_N28
cycloneive_lcell_comb \Mux15~10 (
// Equation(s):
// \Mux15~10_combout  = (Selector5 & (((\register[5][16]~q ) # (Selector41)))) # (!Selector5 & (\register[4][16]~q  & ((!Selector41))))

	.dataa(\register[4][16]~q ),
	.datab(Selector5),
	.datac(\register[5][16]~q ),
	.datad(Selector41),
	.cin(gnd),
	.combout(\Mux15~10_combout ),
	.cout());
// synopsys translate_off
defparam \Mux15~10 .lut_mask = 16'hCCE2;
defparam \Mux15~10 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X68_Y32_N16
cycloneive_lcell_comb \Mux15~11 (
// Equation(s):
// \Mux15~11_combout  = (Selector41 & ((\Mux15~10_combout  & (\register[7][16]~q )) # (!\Mux15~10_combout  & ((\register[6][16]~q ))))) # (!Selector41 & (((\Mux15~10_combout ))))

	.dataa(\register[7][16]~q ),
	.datab(Selector41),
	.datac(\register[6][16]~q ),
	.datad(\Mux15~10_combout ),
	.cin(gnd),
	.combout(\Mux15~11_combout ),
	.cout());
// synopsys translate_off
defparam \Mux15~11 .lut_mask = 16'hBBC0;
defparam \Mux15~11 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y36_N28
cycloneive_lcell_comb \Mux15~17 (
// Equation(s):
// \Mux15~17_combout  = (Selector41 & (Selector5)) # (!Selector41 & ((Selector5 & (\register[13][16]~q )) # (!Selector5 & ((\register[12][16]~q )))))

	.dataa(Selector41),
	.datab(Selector5),
	.datac(\register[13][16]~q ),
	.datad(\register[12][16]~q ),
	.cin(gnd),
	.combout(\Mux15~17_combout ),
	.cout());
// synopsys translate_off
defparam \Mux15~17 .lut_mask = 16'hD9C8;
defparam \Mux15~17 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X65_Y35_N30
cycloneive_lcell_comb \Mux15~18 (
// Equation(s):
// \Mux15~18_combout  = (Selector41 & ((\Mux15~17_combout  & (\register[15][16]~q )) # (!\Mux15~17_combout  & ((\register[14][16]~q ))))) # (!Selector41 & (((\Mux15~17_combout ))))

	.dataa(Selector41),
	.datab(\register[15][16]~q ),
	.datac(\register[14][16]~q ),
	.datad(\Mux15~17_combout ),
	.cin(gnd),
	.combout(\Mux15~18_combout ),
	.cout());
// synopsys translate_off
defparam \Mux15~18 .lut_mask = 16'hDDA0;
defparam \Mux15~18 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X70_Y34_N0
cycloneive_lcell_comb \Mux15~14 (
// Equation(s):
// \Mux15~14_combout  = (Selector4 & ((plif_ifidinstr_l_22 & (\register[3][16]~q )) # (!plif_ifidinstr_l_22 & ((\register[1][16]~q ))))) # (!Selector4 & (((\register[1][16]~q ))))

	.dataa(Selector4),
	.datab(plif_ifidinstr_l_22),
	.datac(\register[3][16]~q ),
	.datad(\register[1][16]~q ),
	.cin(gnd),
	.combout(\Mux15~14_combout ),
	.cout());
// synopsys translate_off
defparam \Mux15~14 .lut_mask = 16'hF780;
defparam \Mux15~14 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X65_Y35_N22
cycloneive_lcell_comb \Mux15~15 (
// Equation(s):
// \Mux15~15_combout  = (Selector5 & (((\Mux15~14_combout )))) # (!Selector5 & (\register[2][16]~q  & (Selector41)))

	.dataa(Selector5),
	.datab(\register[2][16]~q ),
	.datac(Selector41),
	.datad(\Mux15~14_combout ),
	.cin(gnd),
	.combout(\Mux15~15_combout ),
	.cout());
// synopsys translate_off
defparam \Mux15~15 .lut_mask = 16'hEA40;
defparam \Mux15~15 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y40_N4
cycloneive_lcell_comb \Mux15~12 (
// Equation(s):
// \Mux15~12_combout  = (Selector41 & ((Selector5) # ((\register[10][16]~q )))) # (!Selector41 & (!Selector5 & ((\register[8][16]~q ))))

	.dataa(Selector41),
	.datab(Selector5),
	.datac(\register[10][16]~q ),
	.datad(\register[8][16]~q ),
	.cin(gnd),
	.combout(\Mux15~12_combout ),
	.cout());
// synopsys translate_off
defparam \Mux15~12 .lut_mask = 16'hB9A8;
defparam \Mux15~12 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X63_Y40_N8
cycloneive_lcell_comb \Mux15~13 (
// Equation(s):
// \Mux15~13_combout  = (\Mux15~12_combout  & ((\register[11][16]~q ) # ((!Selector5)))) # (!\Mux15~12_combout  & (((\register[9][16]~q  & Selector5))))

	.dataa(\register[11][16]~q ),
	.datab(\Mux15~12_combout ),
	.datac(\register[9][16]~q ),
	.datad(Selector5),
	.cin(gnd),
	.combout(\Mux15~13_combout ),
	.cout());
// synopsys translate_off
defparam \Mux15~13 .lut_mask = 16'hB8CC;
defparam \Mux15~13 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X65_Y35_N28
cycloneive_lcell_comb \Mux15~16 (
// Equation(s):
// \Mux15~16_combout  = (Selector3 & (Selector2)) # (!Selector3 & ((Selector2 & ((\Mux15~13_combout ))) # (!Selector2 & (\Mux15~15_combout ))))

	.dataa(Selector3),
	.datab(Selector2),
	.datac(\Mux15~15_combout ),
	.datad(\Mux15~13_combout ),
	.cin(gnd),
	.combout(\Mux15~16_combout ),
	.cout());
// synopsys translate_off
defparam \Mux15~16 .lut_mask = 16'hDC98;
defparam \Mux15~16 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y33_N6
cycloneive_lcell_comb \Mux16~0 (
// Equation(s):
// \Mux16~0_combout  = (Selector2 & (Selector3)) # (!Selector2 & ((Selector3 & (\register[21][15]~q )) # (!Selector3 & ((\register[17][15]~q )))))

	.dataa(Selector2),
	.datab(Selector3),
	.datac(\register[21][15]~q ),
	.datad(\register[17][15]~q ),
	.cin(gnd),
	.combout(\Mux16~0_combout ),
	.cout());
// synopsys translate_off
defparam \Mux16~0 .lut_mask = 16'hD9C8;
defparam \Mux16~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y40_N12
cycloneive_lcell_comb \Mux16~1 (
// Equation(s):
// \Mux16~1_combout  = (Selector2 & ((\Mux16~0_combout  & ((\register[29][15]~q ))) # (!\Mux16~0_combout  & (\register[25][15]~q )))) # (!Selector2 & (((\Mux16~0_combout ))))

	.dataa(Selector2),
	.datab(\register[25][15]~q ),
	.datac(\register[29][15]~q ),
	.datad(\Mux16~0_combout ),
	.cin(gnd),
	.combout(\Mux16~1_combout ),
	.cout());
// synopsys translate_off
defparam \Mux16~1 .lut_mask = 16'hF588;
defparam \Mux16~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y31_N14
cycloneive_lcell_comb \Mux16~7 (
// Equation(s):
// \Mux16~7_combout  = (Selector3 & ((Selector2) # ((\register[23][15]~q )))) # (!Selector3 & (!Selector2 & (\register[19][15]~q )))

	.dataa(Selector3),
	.datab(Selector2),
	.datac(\register[19][15]~q ),
	.datad(\register[23][15]~q ),
	.cin(gnd),
	.combout(\Mux16~7_combout ),
	.cout());
// synopsys translate_off
defparam \Mux16~7 .lut_mask = 16'hBA98;
defparam \Mux16~7 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y40_N24
cycloneive_lcell_comb \Mux16~8 (
// Equation(s):
// \Mux16~8_combout  = (\Mux16~7_combout  & (((\register[31][15]~q ) # (!Selector2)))) # (!\Mux16~7_combout  & (\register[27][15]~q  & ((Selector2))))

	.dataa(\register[27][15]~q ),
	.datab(\Mux16~7_combout ),
	.datac(\register[31][15]~q ),
	.datad(Selector2),
	.cin(gnd),
	.combout(\Mux16~8_combout ),
	.cout());
// synopsys translate_off
defparam \Mux16~8 .lut_mask = 16'hE2CC;
defparam \Mux16~8 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X69_Y34_N10
cycloneive_lcell_comb \Mux16~4 (
// Equation(s):
// \Mux16~4_combout  = (Selector3 & (Selector2)) # (!Selector3 & ((Selector2 & ((\register[24][15]~q ))) # (!Selector2 & (\register[16][15]~q ))))

	.dataa(Selector3),
	.datab(Selector2),
	.datac(\register[16][15]~q ),
	.datad(\register[24][15]~q ),
	.cin(gnd),
	.combout(\Mux16~4_combout ),
	.cout());
// synopsys translate_off
defparam \Mux16~4 .lut_mask = 16'hDC98;
defparam \Mux16~4 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X69_Y36_N20
cycloneive_lcell_comb \Mux16~5 (
// Equation(s):
// \Mux16~5_combout  = (\Mux16~4_combout  & ((\register[28][15]~q ) # ((!Selector3)))) # (!\Mux16~4_combout  & (((\register[20][15]~q  & Selector3))))

	.dataa(\register[28][15]~q ),
	.datab(\Mux16~4_combout ),
	.datac(\register[20][15]~q ),
	.datad(Selector3),
	.cin(gnd),
	.combout(\Mux16~5_combout ),
	.cout());
// synopsys translate_off
defparam \Mux16~5 .lut_mask = 16'hB8CC;
defparam \Mux16~5 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X68_Y38_N24
cycloneive_lcell_comb \Mux16~2 (
// Equation(s):
// \Mux16~2_combout  = (Selector3 & (((Selector2)))) # (!Selector3 & ((Selector2 & ((\register[26][15]~q ))) # (!Selector2 & (\register[18][15]~q ))))

	.dataa(Selector3),
	.datab(\register[18][15]~q ),
	.datac(\register[26][15]~q ),
	.datad(Selector2),
	.cin(gnd),
	.combout(\Mux16~2_combout ),
	.cout());
// synopsys translate_off
defparam \Mux16~2 .lut_mask = 16'hFA44;
defparam \Mux16~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X69_Y36_N10
cycloneive_lcell_comb \Mux16~3 (
// Equation(s):
// \Mux16~3_combout  = (Selector3 & ((\Mux16~2_combout  & (\register[30][15]~q )) # (!\Mux16~2_combout  & ((\register[22][15]~q ))))) # (!Selector3 & (((\Mux16~2_combout ))))

	.dataa(Selector3),
	.datab(\register[30][15]~q ),
	.datac(\Mux16~2_combout ),
	.datad(\register[22][15]~q ),
	.cin(gnd),
	.combout(\Mux16~3_combout ),
	.cout());
// synopsys translate_off
defparam \Mux16~3 .lut_mask = 16'hDAD0;
defparam \Mux16~3 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y40_N18
cycloneive_lcell_comb \Mux16~6 (
// Equation(s):
// \Mux16~6_combout  = (Selector41 & ((Selector5) # ((\Mux16~3_combout )))) # (!Selector41 & (!Selector5 & (\Mux16~5_combout )))

	.dataa(Selector41),
	.datab(Selector5),
	.datac(\Mux16~5_combout ),
	.datad(\Mux16~3_combout ),
	.cin(gnd),
	.combout(\Mux16~6_combout ),
	.cout());
// synopsys translate_off
defparam \Mux16~6 .lut_mask = 16'hBA98;
defparam \Mux16~6 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X63_Y30_N2
cycloneive_lcell_comb \Mux16~17 (
// Equation(s):
// \Mux16~17_combout  = (Selector5 & ((Selector41) # ((\register[13][15]~q )))) # (!Selector5 & (!Selector41 & (\register[12][15]~q )))

	.dataa(Selector5),
	.datab(Selector41),
	.datac(\register[12][15]~q ),
	.datad(\register[13][15]~q ),
	.cin(gnd),
	.combout(\Mux16~17_combout ),
	.cout());
// synopsys translate_off
defparam \Mux16~17 .lut_mask = 16'hBA98;
defparam \Mux16~17 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y33_N12
cycloneive_lcell_comb \Mux16~18 (
// Equation(s):
// \Mux16~18_combout  = (Selector41 & ((\Mux16~17_combout  & (\register[15][15]~q )) # (!\Mux16~17_combout  & ((\register[14][15]~q ))))) # (!Selector41 & (((\Mux16~17_combout ))))

	.dataa(Selector41),
	.datab(\register[15][15]~q ),
	.datac(\register[14][15]~q ),
	.datad(\Mux16~17_combout ),
	.cin(gnd),
	.combout(\Mux16~18_combout ),
	.cout());
// synopsys translate_off
defparam \Mux16~18 .lut_mask = 16'hDDA0;
defparam \Mux16~18 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X62_Y40_N17
dffeas \register[10][15] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\register~80_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~45_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\register[10][15]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \register[10][15] .is_wysiwyg = "true";
defparam \register[10][15] .power_up = "low";
// synopsys translate_on

// Location: FF_X62_Y40_N11
dffeas \register[8][15] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\register~80_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~46_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\register[8][15]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \register[8][15] .is_wysiwyg = "true";
defparam \register[8][15] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X62_Y40_N10
cycloneive_lcell_comb \Mux16~10 (
// Equation(s):
// \Mux16~10_combout  = (Selector41 & ((\register[10][15]~q ) # ((Selector5)))) # (!Selector41 & (((\register[8][15]~q  & !Selector5))))

	.dataa(Selector41),
	.datab(\register[10][15]~q ),
	.datac(\register[8][15]~q ),
	.datad(Selector5),
	.cin(gnd),
	.combout(\Mux16~10_combout ),
	.cout());
// synopsys translate_off
defparam \Mux16~10 .lut_mask = 16'hAAD8;
defparam \Mux16~10 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X63_Y40_N28
cycloneive_lcell_comb \Mux16~11 (
// Equation(s):
// \Mux16~11_combout  = (\Mux16~10_combout  & ((\register[11][15]~q ) # ((!Selector5)))) # (!\Mux16~10_combout  & (((\register[9][15]~q  & Selector5))))

	.dataa(\Mux16~10_combout ),
	.datab(\register[11][15]~q ),
	.datac(\register[9][15]~q ),
	.datad(Selector5),
	.cin(gnd),
	.combout(\Mux16~11_combout ),
	.cout());
// synopsys translate_off
defparam \Mux16~11 .lut_mask = 16'hD8AA;
defparam \Mux16~11 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X67_Y34_N3
dffeas \register[2][15] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\register~80_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~50_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\register[2][15]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \register[2][15] .is_wysiwyg = "true";
defparam \register[2][15] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X67_Y34_N2
cycloneive_lcell_comb \Mux16~15 (
// Equation(s):
// \Mux16~15_combout  = (\Mux16~14_combout ) # ((!Selector5 & (\register[2][15]~q  & Selector41)))

	.dataa(\Mux16~14_combout ),
	.datab(Selector5),
	.datac(\register[2][15]~q ),
	.datad(Selector41),
	.cin(gnd),
	.combout(\Mux16~15_combout ),
	.cout());
// synopsys translate_off
defparam \Mux16~15 .lut_mask = 16'hBAAA;
defparam \Mux16~15 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X69_Y32_N4
cycloneive_lcell_comb \Mux16~12 (
// Equation(s):
// \Mux16~12_combout  = (Selector41 & (Selector5)) # (!Selector41 & ((Selector5 & (\register[5][15]~q )) # (!Selector5 & ((\register[4][15]~q )))))

	.dataa(Selector41),
	.datab(Selector5),
	.datac(\register[5][15]~q ),
	.datad(\register[4][15]~q ),
	.cin(gnd),
	.combout(\Mux16~12_combout ),
	.cout());
// synopsys translate_off
defparam \Mux16~12 .lut_mask = 16'hD9C8;
defparam \Mux16~12 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X68_Y32_N18
cycloneive_lcell_comb \Mux16~13 (
// Equation(s):
// \Mux16~13_combout  = (Selector41 & ((\Mux16~12_combout  & ((\register[7][15]~q ))) # (!\Mux16~12_combout  & (\register[6][15]~q )))) # (!Selector41 & (((\Mux16~12_combout ))))

	.dataa(Selector41),
	.datab(\register[6][15]~q ),
	.datac(\register[7][15]~q ),
	.datad(\Mux16~12_combout ),
	.cin(gnd),
	.combout(\Mux16~13_combout ),
	.cout());
// synopsys translate_off
defparam \Mux16~13 .lut_mask = 16'hF588;
defparam \Mux16~13 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y40_N20
cycloneive_lcell_comb \Mux16~16 (
// Equation(s):
// \Mux16~16_combout  = (Selector2 & (((Selector3)))) # (!Selector2 & ((Selector3 & ((\Mux16~13_combout ))) # (!Selector3 & (\Mux16~15_combout ))))

	.dataa(Selector2),
	.datab(\Mux16~15_combout ),
	.datac(Selector3),
	.datad(\Mux16~13_combout ),
	.cin(gnd),
	.combout(\Mux16~16_combout ),
	.cout());
// synopsys translate_off
defparam \Mux16~16 .lut_mask = 16'hF4A4;
defparam \Mux16~16 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X65_Y37_N4
cycloneive_lcell_comb \Mux17~4 (
// Equation(s):
// \Mux17~4_combout  = (Selector3 & ((Selector2) # ((\register[20][14]~q )))) # (!Selector3 & (!Selector2 & ((\register[16][14]~q ))))

	.dataa(Selector3),
	.datab(Selector2),
	.datac(\register[20][14]~q ),
	.datad(\register[16][14]~q ),
	.cin(gnd),
	.combout(\Mux17~4_combout ),
	.cout());
// synopsys translate_off
defparam \Mux17~4 .lut_mask = 16'hB9A8;
defparam \Mux17~4 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X68_Y34_N12
cycloneive_lcell_comb \Mux17~5 (
// Equation(s):
// \Mux17~5_combout  = (Selector2 & ((\Mux17~4_combout  & (\register[28][14]~q )) # (!\Mux17~4_combout  & ((\register[24][14]~q ))))) # (!Selector2 & (((\Mux17~4_combout ))))

	.dataa(\register[28][14]~q ),
	.datab(\register[24][14]~q ),
	.datac(Selector2),
	.datad(\Mux17~4_combout ),
	.cin(gnd),
	.combout(\Mux17~5_combout ),
	.cout());
// synopsys translate_off
defparam \Mux17~5 .lut_mask = 16'hAFC0;
defparam \Mux17~5 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X69_Y35_N5
dffeas \register[22][14] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\register~81_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~55_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\register[22][14]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \register[22][14] .is_wysiwyg = "true";
defparam \register[22][14] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X69_Y35_N4
cycloneive_lcell_comb \Mux17~2 (
// Equation(s):
// \Mux17~2_combout  = (Selector2 & (((Selector3)))) # (!Selector2 & ((Selector3 & ((\register[22][14]~q ))) # (!Selector3 & (\register[18][14]~q ))))

	.dataa(Selector2),
	.datab(\register[18][14]~q ),
	.datac(\register[22][14]~q ),
	.datad(Selector3),
	.cin(gnd),
	.combout(\Mux17~2_combout ),
	.cout());
// synopsys translate_off
defparam \Mux17~2 .lut_mask = 16'hFA44;
defparam \Mux17~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X68_Y35_N4
cycloneive_lcell_comb \Mux17~3 (
// Equation(s):
// \Mux17~3_combout  = (Selector2 & ((\Mux17~2_combout  & (\register[30][14]~q )) # (!\Mux17~2_combout  & ((\register[26][14]~q ))))) # (!Selector2 & (((\Mux17~2_combout ))))

	.dataa(\register[30][14]~q ),
	.datab(Selector2),
	.datac(\register[26][14]~q ),
	.datad(\Mux17~2_combout ),
	.cin(gnd),
	.combout(\Mux17~3_combout ),
	.cout());
// synopsys translate_off
defparam \Mux17~3 .lut_mask = 16'hBBC0;
defparam \Mux17~3 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X66_Y30_N12
cycloneive_lcell_comb \Mux17~6 (
// Equation(s):
// \Mux17~6_combout  = (Selector5 & (((Selector41)))) # (!Selector5 & ((Selector41 & ((\Mux17~3_combout ))) # (!Selector41 & (\Mux17~5_combout ))))

	.dataa(Selector5),
	.datab(\Mux17~5_combout ),
	.datac(Selector41),
	.datad(\Mux17~3_combout ),
	.cin(gnd),
	.combout(\Mux17~6_combout ),
	.cout());
// synopsys translate_off
defparam \Mux17~6 .lut_mask = 16'hF4A4;
defparam \Mux17~6 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y38_N20
cycloneive_lcell_comb \register[19][14]~feeder (
// Equation(s):
// \register[19][14]~feeder_combout  = \register~81_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(\register~81_combout ),
	.datad(gnd),
	.cin(gnd),
	.combout(\register[19][14]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \register[19][14]~feeder .lut_mask = 16'hF0F0;
defparam \register[19][14]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X60_Y38_N21
dffeas \register[19][14] (
	.clk(!CLK),
	.d(\register[19][14]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~39_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\register[19][14]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \register[19][14] .is_wysiwyg = "true";
defparam \register[19][14] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X60_Y38_N10
cycloneive_lcell_comb \Mux17~7 (
// Equation(s):
// \Mux17~7_combout  = (Selector3 & (Selector2)) # (!Selector3 & ((Selector2 & (\register[27][14]~q )) # (!Selector2 & ((\register[19][14]~q )))))

	.dataa(Selector3),
	.datab(Selector2),
	.datac(\register[27][14]~q ),
	.datad(\register[19][14]~q ),
	.cin(gnd),
	.combout(\Mux17~7_combout ),
	.cout());
// synopsys translate_off
defparam \Mux17~7 .lut_mask = 16'hD9C8;
defparam \Mux17~7 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X66_Y30_N22
cycloneive_lcell_comb \Mux17~8 (
// Equation(s):
// \Mux17~8_combout  = (Selector3 & ((\Mux17~7_combout  & ((\register[31][14]~q ))) # (!\Mux17~7_combout  & (\register[23][14]~q )))) # (!Selector3 & (((\Mux17~7_combout ))))

	.dataa(\register[23][14]~q ),
	.datab(\register[31][14]~q ),
	.datac(Selector3),
	.datad(\Mux17~7_combout ),
	.cin(gnd),
	.combout(\Mux17~8_combout ),
	.cout());
// synopsys translate_off
defparam \Mux17~8 .lut_mask = 16'hCFA0;
defparam \Mux17~8 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y34_N2
cycloneive_lcell_comb \Mux17~0 (
// Equation(s):
// \Mux17~0_combout  = (Selector3 & (((Selector2)))) # (!Selector3 & ((Selector2 & ((\register[25][14]~q ))) # (!Selector2 & (\register[17][14]~q ))))

	.dataa(\register[17][14]~q ),
	.datab(Selector3),
	.datac(\register[25][14]~q ),
	.datad(Selector2),
	.cin(gnd),
	.combout(\Mux17~0_combout ),
	.cout());
// synopsys translate_off
defparam \Mux17~0 .lut_mask = 16'hFC22;
defparam \Mux17~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X63_Y34_N28
cycloneive_lcell_comb \Mux17~1 (
// Equation(s):
// \Mux17~1_combout  = (\Mux17~0_combout  & (((\register[29][14]~q ) # (!Selector3)))) # (!\Mux17~0_combout  & (\register[21][14]~q  & ((Selector3))))

	.dataa(\register[21][14]~q ),
	.datab(\register[29][14]~q ),
	.datac(\Mux17~0_combout ),
	.datad(Selector3),
	.cin(gnd),
	.combout(\Mux17~1_combout ),
	.cout());
// synopsys translate_off
defparam \Mux17~1 .lut_mask = 16'hCAF0;
defparam \Mux17~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X63_Y30_N20
cycloneive_lcell_comb \Mux17~17 (
// Equation(s):
// \Mux17~17_combout  = (Selector41 & (((Selector5)))) # (!Selector41 & ((Selector5 & ((\register[13][14]~q ))) # (!Selector5 & (\register[12][14]~q ))))

	.dataa(\register[12][14]~q ),
	.datab(Selector41),
	.datac(\register[13][14]~q ),
	.datad(Selector5),
	.cin(gnd),
	.combout(\Mux17~17_combout ),
	.cout());
// synopsys translate_off
defparam \Mux17~17 .lut_mask = 16'hFC22;
defparam \Mux17~17 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y34_N8
cycloneive_lcell_comb \Mux17~18 (
// Equation(s):
// \Mux17~18_combout  = (Selector41 & ((\Mux17~17_combout  & (\register[15][14]~q )) # (!\Mux17~17_combout  & ((\register[14][14]~q ))))) # (!Selector41 & (((\Mux17~17_combout ))))

	.dataa(\register[15][14]~q ),
	.datab(Selector41),
	.datac(\register[14][14]~q ),
	.datad(\Mux17~17_combout ),
	.cin(gnd),
	.combout(\Mux17~18_combout ),
	.cout());
// synopsys translate_off
defparam \Mux17~18 .lut_mask = 16'hBBC0;
defparam \Mux17~18 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X66_Y34_N14
cycloneive_lcell_comb \Mux17~15 (
// Equation(s):
// \Mux17~15_combout  = (Selector5 & (\Mux17~14_combout )) # (!Selector5 & (((\register[2][14]~q  & Selector41))))

	.dataa(\Mux17~14_combout ),
	.datab(Selector5),
	.datac(\register[2][14]~q ),
	.datad(Selector41),
	.cin(gnd),
	.combout(\Mux17~15_combout ),
	.cout());
// synopsys translate_off
defparam \Mux17~15 .lut_mask = 16'hB888;
defparam \Mux17~15 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y40_N20
cycloneive_lcell_comb \Mux17~12 (
// Equation(s):
// \Mux17~12_combout  = (Selector41 & ((Selector5) # ((\register[10][14]~q )))) # (!Selector41 & (!Selector5 & ((\register[8][14]~q ))))

	.dataa(Selector41),
	.datab(Selector5),
	.datac(\register[10][14]~q ),
	.datad(\register[8][14]~q ),
	.cin(gnd),
	.combout(\Mux17~12_combout ),
	.cout());
// synopsys translate_off
defparam \Mux17~12 .lut_mask = 16'hB9A8;
defparam \Mux17~12 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X66_Y34_N28
cycloneive_lcell_comb \Mux17~13 (
// Equation(s):
// \Mux17~13_combout  = (Selector5 & ((\Mux17~12_combout  & ((\register[11][14]~q ))) # (!\Mux17~12_combout  & (\register[9][14]~q )))) # (!Selector5 & (((\Mux17~12_combout ))))

	.dataa(\register[9][14]~q ),
	.datab(Selector5),
	.datac(\register[11][14]~q ),
	.datad(\Mux17~12_combout ),
	.cin(gnd),
	.combout(\Mux17~13_combout ),
	.cout());
// synopsys translate_off
defparam \Mux17~13 .lut_mask = 16'hF388;
defparam \Mux17~13 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X65_Y37_N14
cycloneive_lcell_comb \Mux17~16 (
// Equation(s):
// \Mux17~16_combout  = (Selector3 & (Selector2)) # (!Selector3 & ((Selector2 & ((\Mux17~13_combout ))) # (!Selector2 & (\Mux17~15_combout ))))

	.dataa(Selector3),
	.datab(Selector2),
	.datac(\Mux17~15_combout ),
	.datad(\Mux17~13_combout ),
	.cin(gnd),
	.combout(\Mux17~16_combout ),
	.cout());
// synopsys translate_off
defparam \Mux17~16 .lut_mask = 16'hDC98;
defparam \Mux17~16 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X69_Y32_N24
cycloneive_lcell_comb \Mux17~10 (
// Equation(s):
// \Mux17~10_combout  = (Selector41 & (((Selector5)))) # (!Selector41 & ((Selector5 & ((\register[5][14]~q ))) # (!Selector5 & (\register[4][14]~q ))))

	.dataa(Selector41),
	.datab(\register[4][14]~q ),
	.datac(\register[5][14]~q ),
	.datad(Selector5),
	.cin(gnd),
	.combout(\Mux17~10_combout ),
	.cout());
// synopsys translate_off
defparam \Mux17~10 .lut_mask = 16'hFA44;
defparam \Mux17~10 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X68_Y32_N20
cycloneive_lcell_comb \Mux17~11 (
// Equation(s):
// \Mux17~11_combout  = (Selector41 & ((\Mux17~10_combout  & ((\register[7][14]~q ))) # (!\Mux17~10_combout  & (\register[6][14]~q )))) # (!Selector41 & (\Mux17~10_combout ))

	.dataa(Selector41),
	.datab(\Mux17~10_combout ),
	.datac(\register[6][14]~q ),
	.datad(\register[7][14]~q ),
	.cin(gnd),
	.combout(\Mux17~11_combout ),
	.cout());
// synopsys translate_off
defparam \Mux17~11 .lut_mask = 16'hEC64;
defparam \Mux17~11 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y38_N28
cycloneive_lcell_comb \Mux18~7 (
// Equation(s):
// \Mux18~7_combout  = (Selector3 & ((Selector2) # ((\register[23][13]~q )))) # (!Selector3 & (!Selector2 & (\register[19][13]~q )))

	.dataa(Selector3),
	.datab(Selector2),
	.datac(\register[19][13]~q ),
	.datad(\register[23][13]~q ),
	.cin(gnd),
	.combout(\Mux18~7_combout ),
	.cout());
// synopsys translate_off
defparam \Mux18~7 .lut_mask = 16'hBA98;
defparam \Mux18~7 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X63_Y38_N22
cycloneive_lcell_comb \Mux18~8 (
// Equation(s):
// \Mux18~8_combout  = (\Mux18~7_combout  & (((\register[31][13]~q ) # (!Selector2)))) # (!\Mux18~7_combout  & (\register[27][13]~q  & (Selector2)))

	.dataa(\register[27][13]~q ),
	.datab(\Mux18~7_combout ),
	.datac(Selector2),
	.datad(\register[31][13]~q ),
	.cin(gnd),
	.combout(\Mux18~8_combout ),
	.cout());
// synopsys translate_off
defparam \Mux18~8 .lut_mask = 16'hEC2C;
defparam \Mux18~8 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X68_Y38_N0
cycloneive_lcell_comb \Mux18~2 (
// Equation(s):
// \Mux18~2_combout  = (Selector3 & (((Selector2)))) # (!Selector3 & ((Selector2 & ((\register[26][13]~q ))) # (!Selector2 & (\register[18][13]~q ))))

	.dataa(Selector3),
	.datab(\register[18][13]~q ),
	.datac(\register[26][13]~q ),
	.datad(Selector2),
	.cin(gnd),
	.combout(\Mux18~2_combout ),
	.cout());
// synopsys translate_off
defparam \Mux18~2 .lut_mask = 16'hFA44;
defparam \Mux18~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X68_Y39_N28
cycloneive_lcell_comb \Mux18~3 (
// Equation(s):
// \Mux18~3_combout  = (\Mux18~2_combout  & (((\register[30][13]~q ) # (!Selector3)))) # (!\Mux18~2_combout  & (\register[22][13]~q  & ((Selector3))))

	.dataa(\register[22][13]~q ),
	.datab(\Mux18~2_combout ),
	.datac(\register[30][13]~q ),
	.datad(Selector3),
	.cin(gnd),
	.combout(\Mux18~3_combout ),
	.cout());
// synopsys translate_off
defparam \Mux18~3 .lut_mask = 16'hE2CC;
defparam \Mux18~3 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X65_Y38_N11
dffeas \register[28][13] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\register~82_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~57_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\register[28][13]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \register[28][13] .is_wysiwyg = "true";
defparam \register[28][13] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X65_Y34_N24
cycloneive_lcell_comb \Mux18~4 (
// Equation(s):
// \Mux18~4_combout  = (Selector2 & ((Selector3) # ((\register[24][13]~q )))) # (!Selector2 & (!Selector3 & (\register[16][13]~q )))

	.dataa(Selector2),
	.datab(Selector3),
	.datac(\register[16][13]~q ),
	.datad(\register[24][13]~q ),
	.cin(gnd),
	.combout(\Mux18~4_combout ),
	.cout());
// synopsys translate_off
defparam \Mux18~4 .lut_mask = 16'hBA98;
defparam \Mux18~4 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X65_Y38_N10
cycloneive_lcell_comb \Mux18~5 (
// Equation(s):
// \Mux18~5_combout  = (Selector3 & ((\Mux18~4_combout  & ((\register[28][13]~q ))) # (!\Mux18~4_combout  & (\register[20][13]~q )))) # (!Selector3 & (((\Mux18~4_combout ))))

	.dataa(Selector3),
	.datab(\register[20][13]~q ),
	.datac(\register[28][13]~q ),
	.datad(\Mux18~4_combout ),
	.cin(gnd),
	.combout(\Mux18~5_combout ),
	.cout());
// synopsys translate_off
defparam \Mux18~5 .lut_mask = 16'hF588;
defparam \Mux18~5 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X63_Y38_N20
cycloneive_lcell_comb \Mux18~6 (
// Equation(s):
// \Mux18~6_combout  = (Selector5 & (Selector41)) # (!Selector5 & ((Selector41 & (\Mux18~3_combout )) # (!Selector41 & ((\Mux18~5_combout )))))

	.dataa(Selector5),
	.datab(Selector41),
	.datac(\Mux18~3_combout ),
	.datad(\Mux18~5_combout ),
	.cin(gnd),
	.combout(\Mux18~6_combout ),
	.cout());
// synopsys translate_off
defparam \Mux18~6 .lut_mask = 16'hD9C8;
defparam \Mux18~6 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X63_Y38_N8
cycloneive_lcell_comb \register[25][13]~feeder (
// Equation(s):
// \register[25][13]~feeder_combout  = \register~82_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(\register~82_combout ),
	.cin(gnd),
	.combout(\register[25][13]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \register[25][13]~feeder .lut_mask = 16'hFF00;
defparam \register[25][13]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X63_Y38_N9
dffeas \register[25][13] (
	.clk(!CLK),
	.d(\register[25][13]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~24_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\register[25][13]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \register[25][13] .is_wysiwyg = "true";
defparam \register[25][13] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X63_Y38_N24
cycloneive_lcell_comb \Mux18~0 (
// Equation(s):
// \Mux18~0_combout  = (Selector2 & (((Selector3)))) # (!Selector2 & ((Selector3 & (\register[21][13]~q )) # (!Selector3 & ((\register[17][13]~q )))))

	.dataa(\register[21][13]~q ),
	.datab(\register[17][13]~q ),
	.datac(Selector2),
	.datad(Selector3),
	.cin(gnd),
	.combout(\Mux18~0_combout ),
	.cout());
// synopsys translate_off
defparam \Mux18~0 .lut_mask = 16'hFA0C;
defparam \Mux18~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X63_Y38_N14
cycloneive_lcell_comb \Mux18~1 (
// Equation(s):
// \Mux18~1_combout  = (Selector2 & ((\Mux18~0_combout  & (\register[29][13]~q )) # (!\Mux18~0_combout  & ((\register[25][13]~q ))))) # (!Selector2 & (((\Mux18~0_combout ))))

	.dataa(\register[29][13]~q ),
	.datab(Selector2),
	.datac(\register[25][13]~q ),
	.datad(\Mux18~0_combout ),
	.cin(gnd),
	.combout(\Mux18~1_combout ),
	.cout());
// synopsys translate_off
defparam \Mux18~1 .lut_mask = 16'hBBC0;
defparam \Mux18~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X62_Y40_N27
dffeas \register[8][13] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\register~82_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~46_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\register[8][13]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \register[8][13] .is_wysiwyg = "true";
defparam \register[8][13] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X62_Y40_N26
cycloneive_lcell_comb \Mux18~10 (
// Equation(s):
// \Mux18~10_combout  = (Selector41 & ((\register[10][13]~q ) # ((Selector5)))) # (!Selector41 & (((\register[8][13]~q  & !Selector5))))

	.dataa(Selector41),
	.datab(\register[10][13]~q ),
	.datac(\register[8][13]~q ),
	.datad(Selector5),
	.cin(gnd),
	.combout(\Mux18~10_combout ),
	.cout());
// synopsys translate_off
defparam \Mux18~10 .lut_mask = 16'hAAD8;
defparam \Mux18~10 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X63_Y40_N23
dffeas \register[11][13] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\register~82_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~47_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\register[11][13]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \register[11][13] .is_wysiwyg = "true";
defparam \register[11][13] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X63_Y40_N22
cycloneive_lcell_comb \Mux18~11 (
// Equation(s):
// \Mux18~11_combout  = (\Mux18~10_combout  & (((\register[11][13]~q ) # (!Selector5)))) # (!\Mux18~10_combout  & (\register[9][13]~q  & ((Selector5))))

	.dataa(\Mux18~10_combout ),
	.datab(\register[9][13]~q ),
	.datac(\register[11][13]~q ),
	.datad(Selector5),
	.cin(gnd),
	.combout(\Mux18~11_combout ),
	.cout());
// synopsys translate_off
defparam \Mux18~11 .lut_mask = 16'hE4AA;
defparam \Mux18~11 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X59_Y36_N27
dffeas \register[13][13] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\register~82_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~62_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\register[13][13]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \register[13][13] .is_wysiwyg = "true";
defparam \register[13][13] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X59_Y36_N26
cycloneive_lcell_comb \Mux18~17 (
// Equation(s):
// \Mux18~17_combout  = (Selector41 & (Selector5)) # (!Selector41 & ((Selector5 & (\register[13][13]~q )) # (!Selector5 & ((\register[12][13]~q )))))

	.dataa(Selector41),
	.datab(Selector5),
	.datac(\register[13][13]~q ),
	.datad(\register[12][13]~q ),
	.cin(gnd),
	.combout(\Mux18~17_combout ),
	.cout());
// synopsys translate_off
defparam \Mux18~17 .lut_mask = 16'hD9C8;
defparam \Mux18~17 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y36_N16
cycloneive_lcell_comb \Mux18~18 (
// Equation(s):
// \Mux18~18_combout  = (\Mux18~17_combout  & ((\register[15][13]~q ) # ((!Selector41)))) # (!\Mux18~17_combout  & (((\register[14][13]~q  & Selector41))))

	.dataa(\Mux18~17_combout ),
	.datab(\register[15][13]~q ),
	.datac(\register[14][13]~q ),
	.datad(Selector41),
	.cin(gnd),
	.combout(\Mux18~18_combout ),
	.cout());
// synopsys translate_off
defparam \Mux18~18 .lut_mask = 16'hD8AA;
defparam \Mux18~18 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X69_Y32_N23
dffeas \register[4][13] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\register~82_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~60_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\register[4][13]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \register[4][13] .is_wysiwyg = "true";
defparam \register[4][13] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X69_Y32_N22
cycloneive_lcell_comb \Mux18~12 (
// Equation(s):
// \Mux18~12_combout  = (Selector41 & (Selector5)) # (!Selector41 & ((Selector5 & ((\register[5][13]~q ))) # (!Selector5 & (\register[4][13]~q ))))

	.dataa(Selector41),
	.datab(Selector5),
	.datac(\register[4][13]~q ),
	.datad(\register[5][13]~q ),
	.cin(gnd),
	.combout(\Mux18~12_combout ),
	.cout());
// synopsys translate_off
defparam \Mux18~12 .lut_mask = 16'hDC98;
defparam \Mux18~12 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X68_Y32_N26
cycloneive_lcell_comb \Mux18~13 (
// Equation(s):
// \Mux18~13_combout  = (Selector41 & ((\Mux18~12_combout  & ((\register[7][13]~q ))) # (!\Mux18~12_combout  & (\register[6][13]~q )))) # (!Selector41 & (((\Mux18~12_combout ))))

	.dataa(Selector41),
	.datab(\register[6][13]~q ),
	.datac(\register[7][13]~q ),
	.datad(\Mux18~12_combout ),
	.cin(gnd),
	.combout(\Mux18~13_combout ),
	.cout());
// synopsys translate_off
defparam \Mux18~13 .lut_mask = 16'hF588;
defparam \Mux18~13 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X65_Y36_N13
dffeas \register[3][13] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\register~82_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~48_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\register[3][13]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \register[3][13] .is_wysiwyg = "true";
defparam \register[3][13] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X65_Y36_N12
cycloneive_lcell_comb \Mux18~14 (
// Equation(s):
// \Mux18~14_combout  = (Selector4 & ((plif_ifidinstr_l_22 & (\register[3][13]~q )) # (!plif_ifidinstr_l_22 & ((\register[1][13]~q ))))) # (!Selector4 & (((\register[1][13]~q ))))

	.dataa(Selector4),
	.datab(plif_ifidinstr_l_22),
	.datac(\register[3][13]~q ),
	.datad(\register[1][13]~q ),
	.cin(gnd),
	.combout(\Mux18~14_combout ),
	.cout());
// synopsys translate_off
defparam \Mux18~14 .lut_mask = 16'hF780;
defparam \Mux18~14 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X66_Y34_N16
cycloneive_lcell_comb \Mux18~15 (
// Equation(s):
// \Mux18~15_combout  = (Selector5 & (((\Mux18~14_combout )))) # (!Selector5 & (Selector41 & (\register[2][13]~q )))

	.dataa(Selector41),
	.datab(Selector5),
	.datac(\register[2][13]~q ),
	.datad(\Mux18~14_combout ),
	.cin(gnd),
	.combout(\Mux18~15_combout ),
	.cout());
// synopsys translate_off
defparam \Mux18~15 .lut_mask = 16'hEC20;
defparam \Mux18~15 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X63_Y38_N10
cycloneive_lcell_comb \Mux18~16 (
// Equation(s):
// \Mux18~16_combout  = (Selector3 & ((Selector2) # ((\Mux18~13_combout )))) # (!Selector3 & (!Selector2 & ((\Mux18~15_combout ))))

	.dataa(Selector3),
	.datab(Selector2),
	.datac(\Mux18~13_combout ),
	.datad(\Mux18~15_combout ),
	.cin(gnd),
	.combout(\Mux18~16_combout ),
	.cout());
// synopsys translate_off
defparam \Mux18~16 .lut_mask = 16'hB9A8;
defparam \Mux18~16 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y34_N30
cycloneive_lcell_comb \Mux19~0 (
// Equation(s):
// \Mux19~0_combout  = (Selector3 & (((Selector2)))) # (!Selector3 & ((Selector2 & ((\register[25][12]~q ))) # (!Selector2 & (\register[17][12]~q ))))

	.dataa(\register[17][12]~q ),
	.datab(Selector3),
	.datac(\register[25][12]~q ),
	.datad(Selector2),
	.cin(gnd),
	.combout(\Mux19~0_combout ),
	.cout());
// synopsys translate_off
defparam \Mux19~0 .lut_mask = 16'hFC22;
defparam \Mux19~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X63_Y33_N14
cycloneive_lcell_comb \Mux19~1 (
// Equation(s):
// \Mux19~1_combout  = (\Mux19~0_combout  & (((\register[29][12]~q ) # (!Selector3)))) # (!\Mux19~0_combout  & (\register[21][12]~q  & ((Selector3))))

	.dataa(\register[21][12]~q ),
	.datab(\register[29][12]~q ),
	.datac(\Mux19~0_combout ),
	.datad(Selector3),
	.cin(gnd),
	.combout(\Mux19~1_combout ),
	.cout());
// synopsys translate_off
defparam \Mux19~1 .lut_mask = 16'hCAF0;
defparam \Mux19~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y37_N14
cycloneive_lcell_comb \Mux19~7 (
// Equation(s):
// \Mux19~7_combout  = (Selector3 & (Selector2)) # (!Selector3 & ((Selector2 & ((\register[27][12]~q ))) # (!Selector2 & (\register[19][12]~q ))))

	.dataa(Selector3),
	.datab(Selector2),
	.datac(\register[19][12]~q ),
	.datad(\register[27][12]~q ),
	.cin(gnd),
	.combout(\Mux19~7_combout ),
	.cout());
// synopsys translate_off
defparam \Mux19~7 .lut_mask = 16'hDC98;
defparam \Mux19~7 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y30_N30
cycloneive_lcell_comb \Mux19~8 (
// Equation(s):
// \Mux19~8_combout  = (Selector3 & ((\Mux19~7_combout  & (\register[31][12]~q )) # (!\Mux19~7_combout  & ((\register[23][12]~q ))))) # (!Selector3 & (((\Mux19~7_combout ))))

	.dataa(Selector3),
	.datab(\register[31][12]~q ),
	.datac(\register[23][12]~q ),
	.datad(\Mux19~7_combout ),
	.cin(gnd),
	.combout(\Mux19~8_combout ),
	.cout());
// synopsys translate_off
defparam \Mux19~8 .lut_mask = 16'hDDA0;
defparam \Mux19~8 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X69_Y38_N24
cycloneive_lcell_comb \Mux19~4 (
// Equation(s):
// \Mux19~4_combout  = (Selector2 & (((Selector3)))) # (!Selector2 & ((Selector3 & (\register[20][12]~q )) # (!Selector3 & ((\register[16][12]~q )))))

	.dataa(\register[20][12]~q ),
	.datab(Selector2),
	.datac(\register[16][12]~q ),
	.datad(Selector3),
	.cin(gnd),
	.combout(\Mux19~4_combout ),
	.cout());
// synopsys translate_off
defparam \Mux19~4 .lut_mask = 16'hEE30;
defparam \Mux19~4 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X69_Y36_N30
cycloneive_lcell_comb \Mux19~5 (
// Equation(s):
// \Mux19~5_combout  = (Selector2 & ((\Mux19~4_combout  & (\register[28][12]~q )) # (!\Mux19~4_combout  & ((\register[24][12]~q ))))) # (!Selector2 & (((\Mux19~4_combout ))))

	.dataa(Selector2),
	.datab(\register[28][12]~q ),
	.datac(\Mux19~4_combout ),
	.datad(\register[24][12]~q ),
	.cin(gnd),
	.combout(\Mux19~5_combout ),
	.cout());
// synopsys translate_off
defparam \Mux19~5 .lut_mask = 16'hDAD0;
defparam \Mux19~5 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X69_Y37_N2
cycloneive_lcell_comb \Mux19~3 (
// Equation(s):
// \Mux19~3_combout  = (\Mux19~2_combout  & (((\register[30][12]~q ) # (!Selector2)))) # (!\Mux19~2_combout  & (\register[26][12]~q  & (Selector2)))

	.dataa(\Mux19~2_combout ),
	.datab(\register[26][12]~q ),
	.datac(Selector2),
	.datad(\register[30][12]~q ),
	.cin(gnd),
	.combout(\Mux19~3_combout ),
	.cout());
// synopsys translate_off
defparam \Mux19~3 .lut_mask = 16'hEA4A;
defparam \Mux19~3 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y30_N0
cycloneive_lcell_comb \Mux19~6 (
// Equation(s):
// \Mux19~6_combout  = (Selector41 & ((Selector5) # ((\Mux19~3_combout )))) # (!Selector41 & (!Selector5 & (\Mux19~5_combout )))

	.dataa(Selector41),
	.datab(Selector5),
	.datac(\Mux19~5_combout ),
	.datad(\Mux19~3_combout ),
	.cin(gnd),
	.combout(\Mux19~6_combout ),
	.cout());
// synopsys translate_off
defparam \Mux19~6 .lut_mask = 16'hBA98;
defparam \Mux19~6 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y33_N0
cycloneive_lcell_comb \Mux19~17 (
// Equation(s):
// \Mux19~17_combout  = (Selector41 & (((Selector5)))) # (!Selector41 & ((Selector5 & ((\register[13][12]~q ))) # (!Selector5 & (\register[12][12]~q ))))

	.dataa(\register[12][12]~q ),
	.datab(Selector41),
	.datac(\register[13][12]~q ),
	.datad(Selector5),
	.cin(gnd),
	.combout(\Mux19~17_combout ),
	.cout());
// synopsys translate_off
defparam \Mux19~17 .lut_mask = 16'hFC22;
defparam \Mux19~17 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y34_N20
cycloneive_lcell_comb \Mux19~18 (
// Equation(s):
// \Mux19~18_combout  = (Selector41 & ((\Mux19~17_combout  & (\register[15][12]~q )) # (!\Mux19~17_combout  & ((\register[14][12]~q ))))) # (!Selector41 & (((\Mux19~17_combout ))))

	.dataa(\register[15][12]~q ),
	.datab(Selector41),
	.datac(\register[14][12]~q ),
	.datad(\Mux19~17_combout ),
	.cin(gnd),
	.combout(\Mux19~18_combout ),
	.cout());
// synopsys translate_off
defparam \Mux19~18 .lut_mask = 16'hBBC0;
defparam \Mux19~18 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X69_Y32_N27
dffeas \register[4][12] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\register~83_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~60_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\register[4][12]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \register[4][12] .is_wysiwyg = "true";
defparam \register[4][12] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X69_Y32_N26
cycloneive_lcell_comb \Mux19~10 (
// Equation(s):
// \Mux19~10_combout  = (Selector41 & (Selector5)) # (!Selector41 & ((Selector5 & ((\register[5][12]~q ))) # (!Selector5 & (\register[4][12]~q ))))

	.dataa(Selector41),
	.datab(Selector5),
	.datac(\register[4][12]~q ),
	.datad(\register[5][12]~q ),
	.cin(gnd),
	.combout(\Mux19~10_combout ),
	.cout());
// synopsys translate_off
defparam \Mux19~10 .lut_mask = 16'hDC98;
defparam \Mux19~10 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X69_Y34_N8
cycloneive_lcell_comb \Mux19~11 (
// Equation(s):
// \Mux19~11_combout  = (\Mux19~10_combout  & ((\register[7][12]~q ) # ((!Selector41)))) # (!\Mux19~10_combout  & (((\register[6][12]~q  & Selector41))))

	.dataa(\Mux19~10_combout ),
	.datab(\register[7][12]~q ),
	.datac(\register[6][12]~q ),
	.datad(Selector41),
	.cin(gnd),
	.combout(\Mux19~11_combout ),
	.cout());
// synopsys translate_off
defparam \Mux19~11 .lut_mask = 16'hD8AA;
defparam \Mux19~11 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X65_Y33_N28
cycloneive_lcell_comb \Mux19~14 (
// Equation(s):
// \Mux19~14_combout  = (Selector5 & ((Selector41 & ((\register[3][12]~q ))) # (!Selector41 & (\register[1][12]~q ))))

	.dataa(\register[1][12]~q ),
	.datab(Selector41),
	.datac(\register[3][12]~q ),
	.datad(Selector5),
	.cin(gnd),
	.combout(\Mux19~14_combout ),
	.cout());
// synopsys translate_off
defparam \Mux19~14 .lut_mask = 16'hE200;
defparam \Mux19~14 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X69_Y34_N26
cycloneive_lcell_comb \Mux19~15 (
// Equation(s):
// \Mux19~15_combout  = (\Mux19~14_combout ) # ((\register[2][12]~q  & (!Selector5 & Selector41)))

	.dataa(\register[2][12]~q ),
	.datab(Selector5),
	.datac(\Mux19~14_combout ),
	.datad(Selector41),
	.cin(gnd),
	.combout(\Mux19~15_combout ),
	.cout());
// synopsys translate_off
defparam \Mux19~15 .lut_mask = 16'hF2F0;
defparam \Mux19~15 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y40_N28
cycloneive_lcell_comb \Mux19~12 (
// Equation(s):
// \Mux19~12_combout  = (Selector41 & ((Selector5) # ((\register[10][12]~q )))) # (!Selector41 & (!Selector5 & ((\register[8][12]~q ))))

	.dataa(Selector41),
	.datab(Selector5),
	.datac(\register[10][12]~q ),
	.datad(\register[8][12]~q ),
	.cin(gnd),
	.combout(\Mux19~12_combout ),
	.cout());
// synopsys translate_off
defparam \Mux19~12 .lut_mask = 16'hB9A8;
defparam \Mux19~12 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X63_Y40_N16
cycloneive_lcell_comb \Mux19~13 (
// Equation(s):
// \Mux19~13_combout  = (Selector5 & ((\Mux19~12_combout  & (\register[11][12]~q )) # (!\Mux19~12_combout  & ((\register[9][12]~q ))))) # (!Selector5 & (((\Mux19~12_combout ))))

	.dataa(\register[11][12]~q ),
	.datab(Selector5),
	.datac(\register[9][12]~q ),
	.datad(\Mux19~12_combout ),
	.cin(gnd),
	.combout(\Mux19~13_combout ),
	.cout());
// synopsys translate_off
defparam \Mux19~13 .lut_mask = 16'hBBC0;
defparam \Mux19~13 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X69_Y34_N24
cycloneive_lcell_comb \Mux19~16 (
// Equation(s):
// \Mux19~16_combout  = (Selector3 & (Selector2)) # (!Selector3 & ((Selector2 & ((\Mux19~13_combout ))) # (!Selector2 & (\Mux19~15_combout ))))

	.dataa(Selector3),
	.datab(Selector2),
	.datac(\Mux19~15_combout ),
	.datad(\Mux19~13_combout ),
	.cin(gnd),
	.combout(\Mux19~16_combout ),
	.cout());
// synopsys translate_off
defparam \Mux19~16 .lut_mask = 16'hDC98;
defparam \Mux19~16 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y40_N20
cycloneive_lcell_comb \Mux20~7 (
// Equation(s):
// \Mux20~7_combout  = (Selector3 & ((Selector2) # ((\register[23][11]~q )))) # (!Selector3 & (!Selector2 & ((\register[19][11]~q ))))

	.dataa(Selector3),
	.datab(Selector2),
	.datac(\register[23][11]~q ),
	.datad(\register[19][11]~q ),
	.cin(gnd),
	.combout(\Mux20~7_combout ),
	.cout());
// synopsys translate_off
defparam \Mux20~7 .lut_mask = 16'hB9A8;
defparam \Mux20~7 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y38_N6
cycloneive_lcell_comb \Mux20~8 (
// Equation(s):
// \Mux20~8_combout  = (\Mux20~7_combout  & (((\register[31][11]~q )) # (!Selector2))) # (!\Mux20~7_combout  & (Selector2 & (\register[27][11]~q )))

	.dataa(\Mux20~7_combout ),
	.datab(Selector2),
	.datac(\register[27][11]~q ),
	.datad(\register[31][11]~q ),
	.cin(gnd),
	.combout(\Mux20~8_combout ),
	.cout());
// synopsys translate_off
defparam \Mux20~8 .lut_mask = 16'hEA62;
defparam \Mux20~8 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y33_N20
cycloneive_lcell_comb \Mux20~0 (
// Equation(s):
// \Mux20~0_combout  = (Selector2 & (((Selector3)))) # (!Selector2 & ((Selector3 & ((\register[21][11]~q ))) # (!Selector3 & (\register[17][11]~q ))))

	.dataa(Selector2),
	.datab(\register[17][11]~q ),
	.datac(Selector3),
	.datad(\register[21][11]~q ),
	.cin(gnd),
	.combout(\Mux20~0_combout ),
	.cout());
// synopsys translate_off
defparam \Mux20~0 .lut_mask = 16'hF4A4;
defparam \Mux20~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X63_Y38_N30
cycloneive_lcell_comb \Mux20~1 (
// Equation(s):
// \Mux20~1_combout  = (\Mux20~0_combout  & (((\register[29][11]~q ) # (!Selector2)))) # (!\Mux20~0_combout  & (\register[25][11]~q  & ((Selector2))))

	.dataa(\register[25][11]~q ),
	.datab(\Mux20~0_combout ),
	.datac(\register[29][11]~q ),
	.datad(Selector2),
	.cin(gnd),
	.combout(\Mux20~1_combout ),
	.cout());
// synopsys translate_off
defparam \Mux20~1 .lut_mask = 16'hE2CC;
defparam \Mux20~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X61_Y40_N13
dffeas \register[24][11] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\register~84_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~34_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\register[24][11]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \register[24][11] .is_wysiwyg = "true";
defparam \register[24][11] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X61_Y40_N12
cycloneive_lcell_comb \Mux20~4 (
// Equation(s):
// \Mux20~4_combout  = (Selector3 & (((Selector2)))) # (!Selector3 & ((Selector2 & ((\register[24][11]~q ))) # (!Selector2 & (\register[16][11]~q ))))

	.dataa(Selector3),
	.datab(\register[16][11]~q ),
	.datac(\register[24][11]~q ),
	.datad(Selector2),
	.cin(gnd),
	.combout(\Mux20~4_combout ),
	.cout());
// synopsys translate_off
defparam \Mux20~4 .lut_mask = 16'hFA44;
defparam \Mux20~4 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y38_N26
cycloneive_lcell_comb \Mux20~5 (
// Equation(s):
// \Mux20~5_combout  = (Selector3 & ((\Mux20~4_combout  & (\register[28][11]~q )) # (!\Mux20~4_combout  & ((\register[20][11]~q ))))) # (!Selector3 & (((\Mux20~4_combout ))))

	.dataa(\register[28][11]~q ),
	.datab(Selector3),
	.datac(\register[20][11]~q ),
	.datad(\Mux20~4_combout ),
	.cin(gnd),
	.combout(\Mux20~5_combout ),
	.cout());
// synopsys translate_off
defparam \Mux20~5 .lut_mask = 16'hBBC0;
defparam \Mux20~5 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X68_Y39_N30
cycloneive_lcell_comb \register[22][11]~feeder (
// Equation(s):
// \register[22][11]~feeder_combout  = \register~84_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(\register~84_combout ),
	.datad(gnd),
	.cin(gnd),
	.combout(\register[22][11]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \register[22][11]~feeder .lut_mask = 16'hF0F0;
defparam \register[22][11]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X68_Y39_N31
dffeas \register[22][11] (
	.clk(!CLK),
	.d(\register[22][11]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~55_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\register[22][11]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \register[22][11] .is_wysiwyg = "true";
defparam \register[22][11] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X68_Y38_N4
cycloneive_lcell_comb \Mux20~2 (
// Equation(s):
// \Mux20~2_combout  = (Selector3 & (((Selector2)))) # (!Selector3 & ((Selector2 & ((\register[26][11]~q ))) # (!Selector2 & (\register[18][11]~q ))))

	.dataa(Selector3),
	.datab(\register[18][11]~q ),
	.datac(\register[26][11]~q ),
	.datad(Selector2),
	.cin(gnd),
	.combout(\Mux20~2_combout ),
	.cout());
// synopsys translate_off
defparam \Mux20~2 .lut_mask = 16'hFA44;
defparam \Mux20~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X68_Y39_N4
cycloneive_lcell_comb \Mux20~3 (
// Equation(s):
// \Mux20~3_combout  = (Selector3 & ((\Mux20~2_combout  & ((\register[30][11]~q ))) # (!\Mux20~2_combout  & (\register[22][11]~q )))) # (!Selector3 & (((\Mux20~2_combout ))))

	.dataa(Selector3),
	.datab(\register[22][11]~q ),
	.datac(\register[30][11]~q ),
	.datad(\Mux20~2_combout ),
	.cin(gnd),
	.combout(\Mux20~3_combout ),
	.cout());
// synopsys translate_off
defparam \Mux20~3 .lut_mask = 16'hF588;
defparam \Mux20~3 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X63_Y38_N28
cycloneive_lcell_comb \Mux20~6 (
// Equation(s):
// \Mux20~6_combout  = (Selector5 & (Selector41)) # (!Selector5 & ((Selector41 & ((\Mux20~3_combout ))) # (!Selector41 & (\Mux20~5_combout ))))

	.dataa(Selector5),
	.datab(Selector41),
	.datac(\Mux20~5_combout ),
	.datad(\Mux20~3_combout ),
	.cin(gnd),
	.combout(\Mux20~6_combout ),
	.cout());
// synopsys translate_off
defparam \Mux20~6 .lut_mask = 16'hDC98;
defparam \Mux20~6 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X63_Y30_N10
cycloneive_lcell_comb \Mux20~17 (
// Equation(s):
// \Mux20~17_combout  = (Selector5 & ((Selector41) # ((\register[13][11]~q )))) # (!Selector5 & (!Selector41 & (\register[12][11]~q )))

	.dataa(Selector5),
	.datab(Selector41),
	.datac(\register[12][11]~q ),
	.datad(\register[13][11]~q ),
	.cin(gnd),
	.combout(\Mux20~17_combout ),
	.cout());
// synopsys translate_off
defparam \Mux20~17 .lut_mask = 16'hBA98;
defparam \Mux20~17 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y33_N26
cycloneive_lcell_comb \Mux20~18 (
// Equation(s):
// \Mux20~18_combout  = (Selector41 & ((\Mux20~17_combout  & (\register[15][11]~q )) # (!\Mux20~17_combout  & ((\register[14][11]~q ))))) # (!Selector41 & (\Mux20~17_combout ))

	.dataa(Selector41),
	.datab(\Mux20~17_combout ),
	.datac(\register[15][11]~q ),
	.datad(\register[14][11]~q ),
	.cin(gnd),
	.combout(\Mux20~18_combout ),
	.cout());
// synopsys translate_off
defparam \Mux20~18 .lut_mask = 16'hE6C4;
defparam \Mux20~18 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X65_Y36_N14
cycloneive_lcell_comb \Mux20~14 (
// Equation(s):
// \Mux20~14_combout  = (Selector4 & ((plif_ifidinstr_l_22 & (\register[3][11]~q )) # (!plif_ifidinstr_l_22 & ((\register[1][11]~q ))))) # (!Selector4 & (((\register[1][11]~q ))))

	.dataa(Selector4),
	.datab(\register[3][11]~q ),
	.datac(\register[1][11]~q ),
	.datad(plif_ifidinstr_l_22),
	.cin(gnd),
	.combout(\Mux20~14_combout ),
	.cout());
// synopsys translate_off
defparam \Mux20~14 .lut_mask = 16'hD8F0;
defparam \Mux20~14 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X66_Y34_N30
cycloneive_lcell_comb \Mux20~15 (
// Equation(s):
// \Mux20~15_combout  = (Selector5 & (((\Mux20~14_combout )))) # (!Selector5 & (Selector41 & (\register[2][11]~q )))

	.dataa(Selector41),
	.datab(Selector5),
	.datac(\register[2][11]~q ),
	.datad(\Mux20~14_combout ),
	.cin(gnd),
	.combout(\Mux20~15_combout ),
	.cout());
// synopsys translate_off
defparam \Mux20~15 .lut_mask = 16'hEC20;
defparam \Mux20~15 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X69_Y32_N18
cycloneive_lcell_comb \Mux20~12 (
// Equation(s):
// \Mux20~12_combout  = (Selector41 & (((Selector5)))) # (!Selector41 & ((Selector5 & (\register[5][11]~q )) # (!Selector5 & ((\register[4][11]~q )))))

	.dataa(Selector41),
	.datab(\register[5][11]~q ),
	.datac(\register[4][11]~q ),
	.datad(Selector5),
	.cin(gnd),
	.combout(\Mux20~12_combout ),
	.cout());
// synopsys translate_off
defparam \Mux20~12 .lut_mask = 16'hEE50;
defparam \Mux20~12 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X68_Y32_N22
cycloneive_lcell_comb \Mux20~13 (
// Equation(s):
// \Mux20~13_combout  = (Selector41 & ((\Mux20~12_combout  & ((\register[7][11]~q ))) # (!\Mux20~12_combout  & (\register[6][11]~q )))) # (!Selector41 & (((\Mux20~12_combout ))))

	.dataa(Selector41),
	.datab(\register[6][11]~q ),
	.datac(\register[7][11]~q ),
	.datad(\Mux20~12_combout ),
	.cin(gnd),
	.combout(\Mux20~13_combout ),
	.cout());
// synopsys translate_off
defparam \Mux20~13 .lut_mask = 16'hF588;
defparam \Mux20~13 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X63_Y38_N0
cycloneive_lcell_comb \Mux20~16 (
// Equation(s):
// \Mux20~16_combout  = (Selector3 & ((Selector2) # ((\Mux20~13_combout )))) # (!Selector3 & (!Selector2 & (\Mux20~15_combout )))

	.dataa(Selector3),
	.datab(Selector2),
	.datac(\Mux20~15_combout ),
	.datad(\Mux20~13_combout ),
	.cin(gnd),
	.combout(\Mux20~16_combout ),
	.cout());
// synopsys translate_off
defparam \Mux20~16 .lut_mask = 16'hBA98;
defparam \Mux20~16 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y40_N6
cycloneive_lcell_comb \Mux20~10 (
// Equation(s):
// \Mux20~10_combout  = (Selector41 & ((Selector5) # ((\register[10][11]~q )))) # (!Selector41 & (!Selector5 & (\register[8][11]~q )))

	.dataa(Selector41),
	.datab(Selector5),
	.datac(\register[8][11]~q ),
	.datad(\register[10][11]~q ),
	.cin(gnd),
	.combout(\Mux20~10_combout ),
	.cout());
// synopsys translate_off
defparam \Mux20~10 .lut_mask = 16'hBA98;
defparam \Mux20~10 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X63_Y40_N11
dffeas \register[11][11] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\register~84_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~47_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\register[11][11]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \register[11][11] .is_wysiwyg = "true";
defparam \register[11][11] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X63_Y40_N10
cycloneive_lcell_comb \Mux20~11 (
// Equation(s):
// \Mux20~11_combout  = (\Mux20~10_combout  & (((\register[11][11]~q ) # (!Selector5)))) # (!\Mux20~10_combout  & (\register[9][11]~q  & ((Selector5))))

	.dataa(\Mux20~10_combout ),
	.datab(\register[9][11]~q ),
	.datac(\register[11][11]~q ),
	.datad(Selector5),
	.cin(gnd),
	.combout(\Mux20~11_combout ),
	.cout());
// synopsys translate_off
defparam \Mux20~11 .lut_mask = 16'hE4AA;
defparam \Mux20~11 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X60_Y37_N21
dffeas \register[17][10] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\register~85_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~26_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\register[17][10]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \register[17][10] .is_wysiwyg = "true";
defparam \register[17][10] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X60_Y37_N20
cycloneive_lcell_comb \Mux21~0 (
// Equation(s):
// \Mux21~0_combout  = (Selector3 & (Selector2)) # (!Selector3 & ((Selector2 & ((\register[25][10]~q ))) # (!Selector2 & (\register[17][10]~q ))))

	.dataa(Selector3),
	.datab(Selector2),
	.datac(\register[17][10]~q ),
	.datad(\register[25][10]~q ),
	.cin(gnd),
	.combout(\Mux21~0_combout ),
	.cout());
// synopsys translate_off
defparam \Mux21~0 .lut_mask = 16'hDC98;
defparam \Mux21~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y34_N18
cycloneive_lcell_comb \Mux21~1 (
// Equation(s):
// \Mux21~1_combout  = (\Mux21~0_combout  & (((\register[29][10]~q )) # (!Selector3))) # (!\Mux21~0_combout  & (Selector3 & ((\register[21][10]~q ))))

	.dataa(\Mux21~0_combout ),
	.datab(Selector3),
	.datac(\register[29][10]~q ),
	.datad(\register[21][10]~q ),
	.cin(gnd),
	.combout(\Mux21~1_combout ),
	.cout());
// synopsys translate_off
defparam \Mux21~1 .lut_mask = 16'hE6A2;
defparam \Mux21~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X69_Y35_N1
dffeas \register[22][10] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\register~85_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~55_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\register[22][10]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \register[22][10] .is_wysiwyg = "true";
defparam \register[22][10] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X69_Y35_N0
cycloneive_lcell_comb \Mux21~2 (
// Equation(s):
// \Mux21~2_combout  = (Selector3 & (((\register[22][10]~q ) # (Selector2)))) # (!Selector3 & (\register[18][10]~q  & ((!Selector2))))

	.dataa(\register[18][10]~q ),
	.datab(Selector3),
	.datac(\register[22][10]~q ),
	.datad(Selector2),
	.cin(gnd),
	.combout(\Mux21~2_combout ),
	.cout());
// synopsys translate_off
defparam \Mux21~2 .lut_mask = 16'hCCE2;
defparam \Mux21~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X68_Y39_N6
cycloneive_lcell_comb \Mux21~3 (
// Equation(s):
// \Mux21~3_combout  = (Selector2 & ((\Mux21~2_combout  & ((\register[30][10]~q ))) # (!\Mux21~2_combout  & (\register[26][10]~q )))) # (!Selector2 & (((\Mux21~2_combout ))))

	.dataa(Selector2),
	.datab(\register[26][10]~q ),
	.datac(\register[30][10]~q ),
	.datad(\Mux21~2_combout ),
	.cin(gnd),
	.combout(\Mux21~3_combout ),
	.cout());
// synopsys translate_off
defparam \Mux21~3 .lut_mask = 16'hF588;
defparam \Mux21~3 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X66_Y36_N30
cycloneive_lcell_comb \register[20][10]~feeder (
// Equation(s):
// \register[20][10]~feeder_combout  = \register~85_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(\register~85_combout ),
	.datad(gnd),
	.cin(gnd),
	.combout(\register[20][10]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \register[20][10]~feeder .lut_mask = 16'hF0F0;
defparam \register[20][10]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X66_Y36_N31
dffeas \register[20][10] (
	.clk(!CLK),
	.d(\register[20][10]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~35_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\register[20][10]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \register[20][10] .is_wysiwyg = "true";
defparam \register[20][10] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X66_Y36_N22
cycloneive_lcell_comb \Mux21~4 (
// Equation(s):
// \Mux21~4_combout  = (Selector2 & (((Selector3)))) # (!Selector2 & ((Selector3 & ((\register[20][10]~q ))) # (!Selector3 & (\register[16][10]~q ))))

	.dataa(\register[16][10]~q ),
	.datab(Selector2),
	.datac(\register[20][10]~q ),
	.datad(Selector3),
	.cin(gnd),
	.combout(\Mux21~4_combout ),
	.cout());
// synopsys translate_off
defparam \Mux21~4 .lut_mask = 16'hFC22;
defparam \Mux21~4 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X66_Y36_N12
cycloneive_lcell_comb \Mux21~5 (
// Equation(s):
// \Mux21~5_combout  = (Selector2 & ((\Mux21~4_combout  & (\register[28][10]~q )) # (!\Mux21~4_combout  & ((\register[24][10]~q ))))) # (!Selector2 & (((\Mux21~4_combout ))))

	.dataa(\register[28][10]~q ),
	.datab(Selector2),
	.datac(\Mux21~4_combout ),
	.datad(\register[24][10]~q ),
	.cin(gnd),
	.combout(\Mux21~5_combout ),
	.cout());
// synopsys translate_off
defparam \Mux21~5 .lut_mask = 16'hBCB0;
defparam \Mux21~5 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X66_Y36_N14
cycloneive_lcell_comb \Mux21~6 (
// Equation(s):
// \Mux21~6_combout  = (Selector5 & (Selector41)) # (!Selector5 & ((Selector41 & (\Mux21~3_combout )) # (!Selector41 & ((\Mux21~5_combout )))))

	.dataa(Selector5),
	.datab(Selector41),
	.datac(\Mux21~3_combout ),
	.datad(\Mux21~5_combout ),
	.cin(gnd),
	.combout(\Mux21~6_combout ),
	.cout());
// synopsys translate_off
defparam \Mux21~6 .lut_mask = 16'hD9C8;
defparam \Mux21~6 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y39_N8
cycloneive_lcell_comb \Mux21~7 (
// Equation(s):
// \Mux21~7_combout  = (Selector3 & (((Selector2)))) # (!Selector3 & ((Selector2 & ((\register[27][10]~q ))) # (!Selector2 & (\register[19][10]~q ))))

	.dataa(Selector3),
	.datab(\register[19][10]~q ),
	.datac(\register[27][10]~q ),
	.datad(Selector2),
	.cin(gnd),
	.combout(\Mux21~7_combout ),
	.cout());
// synopsys translate_off
defparam \Mux21~7 .lut_mask = 16'hFA44;
defparam \Mux21~7 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y38_N28
cycloneive_lcell_comb \Mux21~8 (
// Equation(s):
// \Mux21~8_combout  = (Selector3 & ((\Mux21~7_combout  & (\register[31][10]~q )) # (!\Mux21~7_combout  & ((\register[23][10]~q ))))) # (!Selector3 & (((\Mux21~7_combout ))))

	.dataa(\register[31][10]~q ),
	.datab(Selector3),
	.datac(\register[23][10]~q ),
	.datad(\Mux21~7_combout ),
	.cin(gnd),
	.combout(\Mux21~8_combout ),
	.cout());
// synopsys translate_off
defparam \Mux21~8 .lut_mask = 16'hBBC0;
defparam \Mux21~8 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X67_Y33_N12
cycloneive_lcell_comb \register[6][10]~feeder (
// Equation(s):
// \register[6][10]~feeder_combout  = \register~85_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(\register~85_combout ),
	.cin(gnd),
	.combout(\register[6][10]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \register[6][10]~feeder .lut_mask = 16'hFF00;
defparam \register[6][10]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X67_Y33_N13
dffeas \register[6][10] (
	.clk(!CLK),
	.d(\register[6][10]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~58_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\register[6][10]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \register[6][10] .is_wysiwyg = "true";
defparam \register[6][10] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X67_Y32_N0
cycloneive_lcell_comb \Mux21~10 (
// Equation(s):
// \Mux21~10_combout  = (Selector41 & (Selector5)) # (!Selector41 & ((Selector5 & (\register[5][10]~q )) # (!Selector5 & ((\register[4][10]~q )))))

	.dataa(Selector41),
	.datab(Selector5),
	.datac(\register[5][10]~q ),
	.datad(\register[4][10]~q ),
	.cin(gnd),
	.combout(\Mux21~10_combout ),
	.cout());
// synopsys translate_off
defparam \Mux21~10 .lut_mask = 16'hD9C8;
defparam \Mux21~10 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X67_Y33_N28
cycloneive_lcell_comb \Mux21~11 (
// Equation(s):
// \Mux21~11_combout  = (\Mux21~10_combout  & (((\register[7][10]~q ) # (!Selector41)))) # (!\Mux21~10_combout  & (\register[6][10]~q  & (Selector41)))

	.dataa(\register[6][10]~q ),
	.datab(\Mux21~10_combout ),
	.datac(Selector41),
	.datad(\register[7][10]~q ),
	.cin(gnd),
	.combout(\Mux21~11_combout ),
	.cout());
// synopsys translate_off
defparam \Mux21~11 .lut_mask = 16'hEC2C;
defparam \Mux21~11 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y33_N28
cycloneive_lcell_comb \Mux21~17 (
// Equation(s):
// \Mux21~17_combout  = (Selector41 & (((Selector5)))) # (!Selector41 & ((Selector5 & ((\register[13][10]~q ))) # (!Selector5 & (\register[12][10]~q ))))

	.dataa(\register[12][10]~q ),
	.datab(Selector41),
	.datac(\register[13][10]~q ),
	.datad(Selector5),
	.cin(gnd),
	.combout(\Mux21~17_combout ),
	.cout());
// synopsys translate_off
defparam \Mux21~17 .lut_mask = 16'hFC22;
defparam \Mux21~17 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X65_Y35_N6
cycloneive_lcell_comb \Mux21~18 (
// Equation(s):
// \Mux21~18_combout  = (Selector41 & ((\Mux21~17_combout  & ((\register[15][10]~q ))) # (!\Mux21~17_combout  & (\register[14][10]~q )))) # (!Selector41 & (((\Mux21~17_combout ))))

	.dataa(Selector41),
	.datab(\register[14][10]~q ),
	.datac(\register[15][10]~q ),
	.datad(\Mux21~17_combout ),
	.cin(gnd),
	.combout(\Mux21~18_combout ),
	.cout());
// synopsys translate_off
defparam \Mux21~18 .lut_mask = 16'hF588;
defparam \Mux21~18 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X63_Y40_N2
cycloneive_lcell_comb \Mux21~13 (
// Equation(s):
// \Mux21~13_combout  = (\Mux21~12_combout  & (((\register[11][10]~q ) # (!Selector5)))) # (!\Mux21~12_combout  & (\register[9][10]~q  & ((Selector5))))

	.dataa(\Mux21~12_combout ),
	.datab(\register[9][10]~q ),
	.datac(\register[11][10]~q ),
	.datad(Selector5),
	.cin(gnd),
	.combout(\Mux21~13_combout ),
	.cout());
// synopsys translate_off
defparam \Mux21~13 .lut_mask = 16'hE4AA;
defparam \Mux21~13 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X65_Y33_N18
cycloneive_lcell_comb \Mux21~14 (
// Equation(s):
// \Mux21~14_combout  = (Selector5 & ((Selector41 & (\register[3][10]~q )) # (!Selector41 & ((\register[1][10]~q )))))

	.dataa(Selector41),
	.datab(\register[3][10]~q ),
	.datac(\register[1][10]~q ),
	.datad(Selector5),
	.cin(gnd),
	.combout(\Mux21~14_combout ),
	.cout());
// synopsys translate_off
defparam \Mux21~14 .lut_mask = 16'hD800;
defparam \Mux21~14 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X66_Y36_N18
cycloneive_lcell_comb \Mux21~15 (
// Equation(s):
// \Mux21~15_combout  = (\Mux21~14_combout ) # ((!Selector5 & (\register[2][10]~q  & Selector41)))

	.dataa(Selector5),
	.datab(\register[2][10]~q ),
	.datac(\Mux21~14_combout ),
	.datad(Selector41),
	.cin(gnd),
	.combout(\Mux21~15_combout ),
	.cout());
// synopsys translate_off
defparam \Mux21~15 .lut_mask = 16'hF4F0;
defparam \Mux21~15 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X66_Y36_N20
cycloneive_lcell_comb \Mux21~16 (
// Equation(s):
// \Mux21~16_combout  = (Selector3 & (Selector2)) # (!Selector3 & ((Selector2 & (\Mux21~13_combout )) # (!Selector2 & ((\Mux21~15_combout )))))

	.dataa(Selector3),
	.datab(Selector2),
	.datac(\Mux21~13_combout ),
	.datad(\Mux21~15_combout ),
	.cin(gnd),
	.combout(\Mux21~16_combout ),
	.cout());
// synopsys translate_off
defparam \Mux21~16 .lut_mask = 16'hD9C8;
defparam \Mux21~16 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y35_N26
cycloneive_lcell_comb \Mux22~7 (
// Equation(s):
// \Mux22~7_combout  = (Selector2 & (Selector3)) # (!Selector2 & ((Selector3 & (\register[23][9]~q )) # (!Selector3 & ((\register[19][9]~q )))))

	.dataa(Selector2),
	.datab(Selector3),
	.datac(\register[23][9]~q ),
	.datad(\register[19][9]~q ),
	.cin(gnd),
	.combout(\Mux22~7_combout ),
	.cout());
// synopsys translate_off
defparam \Mux22~7 .lut_mask = 16'hD9C8;
defparam \Mux22~7 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y41_N26
cycloneive_lcell_comb \Mux22~8 (
// Equation(s):
// \Mux22~8_combout  = (Selector2 & ((\Mux22~7_combout  & (\register[31][9]~q )) # (!\Mux22~7_combout  & ((\register[27][9]~q ))))) # (!Selector2 & (((\Mux22~7_combout ))))

	.dataa(Selector2),
	.datab(\register[31][9]~q ),
	.datac(\register[27][9]~q ),
	.datad(\Mux22~7_combout ),
	.cin(gnd),
	.combout(\Mux22~8_combout ),
	.cout());
// synopsys translate_off
defparam \Mux22~8 .lut_mask = 16'hDDA0;
defparam \Mux22~8 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X60_Y37_N3
dffeas \register[17][9] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\register~86_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~26_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\register[17][9]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \register[17][9] .is_wysiwyg = "true";
defparam \register[17][9] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X60_Y37_N2
cycloneive_lcell_comb \Mux22~0 (
// Equation(s):
// \Mux22~0_combout  = (Selector3 & ((Selector2) # ((\register[21][9]~q )))) # (!Selector3 & (!Selector2 & (\register[17][9]~q )))

	.dataa(Selector3),
	.datab(Selector2),
	.datac(\register[17][9]~q ),
	.datad(\register[21][9]~q ),
	.cin(gnd),
	.combout(\Mux22~0_combout ),
	.cout());
// synopsys translate_off
defparam \Mux22~0 .lut_mask = 16'hBA98;
defparam \Mux22~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y34_N30
cycloneive_lcell_comb \Mux22~1 (
// Equation(s):
// \Mux22~1_combout  = (Selector2 & ((\Mux22~0_combout  & ((\register[29][9]~q ))) # (!\Mux22~0_combout  & (\register[25][9]~q )))) # (!Selector2 & (((\Mux22~0_combout ))))

	.dataa(Selector2),
	.datab(\register[25][9]~q ),
	.datac(\register[29][9]~q ),
	.datad(\Mux22~0_combout ),
	.cin(gnd),
	.combout(\Mux22~1_combout ),
	.cout());
// synopsys translate_off
defparam \Mux22~1 .lut_mask = 16'hF588;
defparam \Mux22~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y40_N6
cycloneive_lcell_comb \register[24][9]~feeder (
// Equation(s):
// \register[24][9]~feeder_combout  = \register~86_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(\register~86_combout ),
	.datad(gnd),
	.cin(gnd),
	.combout(\register[24][9]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \register[24][9]~feeder .lut_mask = 16'hF0F0;
defparam \register[24][9]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X61_Y40_N7
dffeas \register[24][9] (
	.clk(!CLK),
	.d(\register[24][9]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~34_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\register[24][9]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \register[24][9] .is_wysiwyg = "true";
defparam \register[24][9] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X65_Y39_N12
cycloneive_lcell_comb \Mux22~4 (
// Equation(s):
// \Mux22~4_combout  = (Selector2 & ((\register[24][9]~q ) # ((Selector3)))) # (!Selector2 & (((\register[16][9]~q  & !Selector3))))

	.dataa(Selector2),
	.datab(\register[24][9]~q ),
	.datac(\register[16][9]~q ),
	.datad(Selector3),
	.cin(gnd),
	.combout(\Mux22~4_combout ),
	.cout());
// synopsys translate_off
defparam \Mux22~4 .lut_mask = 16'hAAD8;
defparam \Mux22~4 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y41_N10
cycloneive_lcell_comb \Mux22~5 (
// Equation(s):
// \Mux22~5_combout  = (\Mux22~4_combout  & (((\register[28][9]~q ) # (!Selector3)))) # (!\Mux22~4_combout  & (\register[20][9]~q  & (Selector3)))

	.dataa(\register[20][9]~q ),
	.datab(\Mux22~4_combout ),
	.datac(Selector3),
	.datad(\register[28][9]~q ),
	.cin(gnd),
	.combout(\Mux22~5_combout ),
	.cout());
// synopsys translate_off
defparam \Mux22~5 .lut_mask = 16'hEC2C;
defparam \Mux22~5 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X69_Y37_N23
dffeas \register[22][9] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\register~86_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~55_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\register[22][9]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \register[22][9] .is_wysiwyg = "true";
defparam \register[22][9] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X69_Y36_N6
cycloneive_lcell_comb \register[30][9]~feeder (
// Equation(s):
// \register[30][9]~feeder_combout  = \register~86_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(\register~86_combout ),
	.cin(gnd),
	.combout(\register[30][9]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \register[30][9]~feeder .lut_mask = 16'hFF00;
defparam \register[30][9]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X69_Y36_N7
dffeas \register[30][9] (
	.clk(!CLK),
	.d(\register[30][9]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~56_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\register[30][9]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \register[30][9] .is_wysiwyg = "true";
defparam \register[30][9] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X69_Y37_N22
cycloneive_lcell_comb \Mux22~3 (
// Equation(s):
// \Mux22~3_combout  = (\Mux22~2_combout  & (((\register[30][9]~q )) # (!Selector3))) # (!\Mux22~2_combout  & (Selector3 & (\register[22][9]~q )))

	.dataa(\Mux22~2_combout ),
	.datab(Selector3),
	.datac(\register[22][9]~q ),
	.datad(\register[30][9]~q ),
	.cin(gnd),
	.combout(\Mux22~3_combout ),
	.cout());
// synopsys translate_off
defparam \Mux22~3 .lut_mask = 16'hEA62;
defparam \Mux22~3 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y41_N16
cycloneive_lcell_comb \Mux22~6 (
// Equation(s):
// \Mux22~6_combout  = (Selector5 & (((Selector41)))) # (!Selector5 & ((Selector41 & ((\Mux22~3_combout ))) # (!Selector41 & (\Mux22~5_combout ))))

	.dataa(\Mux22~5_combout ),
	.datab(Selector5),
	.datac(\Mux22~3_combout ),
	.datad(Selector41),
	.cin(gnd),
	.combout(\Mux22~6_combout ),
	.cout());
// synopsys translate_off
defparam \Mux22~6 .lut_mask = 16'hFC22;
defparam \Mux22~6 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y33_N24
cycloneive_lcell_comb \Mux22~17 (
// Equation(s):
// \Mux22~17_combout  = (Selector5 & (((\register[13][9]~q ) # (Selector41)))) # (!Selector5 & (\register[12][9]~q  & ((!Selector41))))

	.dataa(Selector5),
	.datab(\register[12][9]~q ),
	.datac(\register[13][9]~q ),
	.datad(Selector41),
	.cin(gnd),
	.combout(\Mux22~17_combout ),
	.cout());
// synopsys translate_off
defparam \Mux22~17 .lut_mask = 16'hAAE4;
defparam \Mux22~17 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y41_N24
cycloneive_lcell_comb \Mux22~18 (
// Equation(s):
// \Mux22~18_combout  = (\Mux22~17_combout  & ((\register[15][9]~q ) # ((!Selector41)))) # (!\Mux22~17_combout  & (((\register[14][9]~q  & Selector41))))

	.dataa(\register[15][9]~q ),
	.datab(\register[14][9]~q ),
	.datac(\Mux22~17_combout ),
	.datad(Selector41),
	.cin(gnd),
	.combout(\Mux22~18_combout ),
	.cout());
// synopsys translate_off
defparam \Mux22~18 .lut_mask = 16'hACF0;
defparam \Mux22~18 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y41_N28
cycloneive_lcell_comb \Mux22~10 (
// Equation(s):
// \Mux22~10_combout  = (Selector41 & ((Selector5) # ((\register[10][9]~q )))) # (!Selector41 & (!Selector5 & ((\register[8][9]~q ))))

	.dataa(Selector41),
	.datab(Selector5),
	.datac(\register[10][9]~q ),
	.datad(\register[8][9]~q ),
	.cin(gnd),
	.combout(\Mux22~10_combout ),
	.cout());
// synopsys translate_off
defparam \Mux22~10 .lut_mask = 16'hB9A8;
defparam \Mux22~10 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X65_Y41_N20
cycloneive_lcell_comb \Mux22~11 (
// Equation(s):
// \Mux22~11_combout  = (\Mux22~10_combout  & ((\register[11][9]~q ) # ((!Selector5)))) # (!\Mux22~10_combout  & (((\register[9][9]~q  & Selector5))))

	.dataa(\register[11][9]~q ),
	.datab(\Mux22~10_combout ),
	.datac(\register[9][9]~q ),
	.datad(Selector5),
	.cin(gnd),
	.combout(\Mux22~11_combout ),
	.cout());
// synopsys translate_off
defparam \Mux22~11 .lut_mask = 16'hB8CC;
defparam \Mux22~11 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X69_Y33_N28
cycloneive_lcell_comb \Mux22~14 (
// Equation(s):
// \Mux22~14_combout  = (plif_ifidinstr_l_22 & ((Selector4 & ((\register[3][9]~q ))) # (!Selector4 & (\register[1][9]~q )))) # (!plif_ifidinstr_l_22 & (\register[1][9]~q ))

	.dataa(\register[1][9]~q ),
	.datab(plif_ifidinstr_l_22),
	.datac(\register[3][9]~q ),
	.datad(Selector4),
	.cin(gnd),
	.combout(\Mux22~14_combout ),
	.cout());
// synopsys translate_off
defparam \Mux22~14 .lut_mask = 16'hE2AA;
defparam \Mux22~14 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y41_N18
cycloneive_lcell_comb \Mux22~15 (
// Equation(s):
// \Mux22~15_combout  = (Selector5 & (((\Mux22~14_combout )))) # (!Selector5 & (\register[2][9]~q  & (Selector41)))

	.dataa(\register[2][9]~q ),
	.datab(Selector41),
	.datac(Selector5),
	.datad(\Mux22~14_combout ),
	.cin(gnd),
	.combout(\Mux22~15_combout ),
	.cout());
// synopsys translate_off
defparam \Mux22~15 .lut_mask = 16'hF808;
defparam \Mux22~15 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X67_Y32_N24
cycloneive_lcell_comb \Mux22~12 (
// Equation(s):
// \Mux22~12_combout  = (Selector41 & (((Selector5)))) # (!Selector41 & ((Selector5 & ((\register[5][9]~q ))) # (!Selector5 & (\register[4][9]~q ))))

	.dataa(\register[4][9]~q ),
	.datab(Selector41),
	.datac(\register[5][9]~q ),
	.datad(Selector5),
	.cin(gnd),
	.combout(\Mux22~12_combout ),
	.cout());
// synopsys translate_off
defparam \Mux22~12 .lut_mask = 16'hFC22;
defparam \Mux22~12 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X68_Y33_N18
cycloneive_lcell_comb \Mux22~13 (
// Equation(s):
// \Mux22~13_combout  = (Selector41 & ((\Mux22~12_combout  & ((\register[7][9]~q ))) # (!\Mux22~12_combout  & (\register[6][9]~q )))) # (!Selector41 & (((\Mux22~12_combout ))))

	.dataa(Selector41),
	.datab(\register[6][9]~q ),
	.datac(\register[7][9]~q ),
	.datad(\Mux22~12_combout ),
	.cin(gnd),
	.combout(\Mux22~13_combout ),
	.cout());
// synopsys translate_off
defparam \Mux22~13 .lut_mask = 16'hF588;
defparam \Mux22~13 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y41_N0
cycloneive_lcell_comb \Mux22~16 (
// Equation(s):
// \Mux22~16_combout  = (Selector2 & (((Selector3)))) # (!Selector2 & ((Selector3 & ((\Mux22~13_combout ))) # (!Selector3 & (\Mux22~15_combout ))))

	.dataa(Selector2),
	.datab(\Mux22~15_combout ),
	.datac(Selector3),
	.datad(\Mux22~13_combout ),
	.cin(gnd),
	.combout(\Mux22~16_combout ),
	.cout());
// synopsys translate_off
defparam \Mux22~16 .lut_mask = 16'hF4A4;
defparam \Mux22~16 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y37_N22
cycloneive_lcell_comb \register[17][4]~feeder (
// Equation(s):
// \register[17][4]~feeder_combout  = \register~94_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(\register~94_combout ),
	.datad(gnd),
	.cin(gnd),
	.combout(\register[17][4]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \register[17][4]~feeder .lut_mask = 16'hF0F0;
defparam \register[17][4]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X60_Y37_N23
dffeas \register[17][4] (
	.clk(!CLK),
	.d(\register[17][4]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~26_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\register[17][4]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \register[17][4] .is_wysiwyg = "true";
defparam \register[17][4] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X60_Y37_N26
cycloneive_lcell_comb \Mux59~0 (
// Equation(s):
// \Mux59~0_combout  = (Selector8 & ((\register[21][4]~q ) # ((Selector7)))) # (!Selector8 & (((!Selector7 & \register[17][4]~q ))))

	.dataa(Selector8),
	.datab(\register[21][4]~q ),
	.datac(Selector7),
	.datad(\register[17][4]~q ),
	.cin(gnd),
	.combout(\Mux59~0_combout ),
	.cout());
// synopsys translate_off
defparam \Mux59~0 .lut_mask = 16'hADA8;
defparam \Mux59~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y41_N28
cycloneive_lcell_comb \Mux59~1 (
// Equation(s):
// \Mux59~1_combout  = (Selector7 & ((\Mux59~0_combout  & ((\register[29][4]~q ))) # (!\Mux59~0_combout  & (\register[25][4]~q )))) # (!Selector7 & (((\Mux59~0_combout ))))

	.dataa(\register[25][4]~q ),
	.datab(\register[29][4]~q ),
	.datac(Selector7),
	.datad(\Mux59~0_combout ),
	.cin(gnd),
	.combout(\Mux59~1_combout ),
	.cout());
// synopsys translate_off
defparam \Mux59~1 .lut_mask = 16'hCFA0;
defparam \Mux59~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y37_N16
cycloneive_lcell_comb \Mux59~7 (
// Equation(s):
// \Mux59~7_combout  = (Selector8 & ((Selector7) # ((\register[23][4]~q )))) # (!Selector8 & (!Selector7 & (\register[19][4]~q )))

	.dataa(Selector8),
	.datab(Selector7),
	.datac(\register[19][4]~q ),
	.datad(\register[23][4]~q ),
	.cin(gnd),
	.combout(\Mux59~7_combout ),
	.cout());
// synopsys translate_off
defparam \Mux59~7 .lut_mask = 16'hBA98;
defparam \Mux59~7 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y41_N14
cycloneive_lcell_comb \Mux59~8 (
// Equation(s):
// \Mux59~8_combout  = (Selector7 & ((\Mux59~7_combout  & (\register[31][4]~q )) # (!\Mux59~7_combout  & ((\register[27][4]~q ))))) # (!Selector7 & (((\Mux59~7_combout ))))

	.dataa(\register[31][4]~q ),
	.datab(Selector7),
	.datac(\Mux59~7_combout ),
	.datad(\register[27][4]~q ),
	.cin(gnd),
	.combout(\Mux59~8_combout ),
	.cout());
// synopsys translate_off
defparam \Mux59~8 .lut_mask = 16'hBCB0;
defparam \Mux59~8 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X68_Y37_N8
cycloneive_lcell_comb \Mux59~2 (
// Equation(s):
// \Mux59~2_combout  = (Selector8 & (((Selector7)))) # (!Selector8 & ((Selector7 & ((\register[26][4]~q ))) # (!Selector7 & (\register[18][4]~q ))))

	.dataa(\register[18][4]~q ),
	.datab(Selector8),
	.datac(\register[26][4]~q ),
	.datad(Selector7),
	.cin(gnd),
	.combout(\Mux59~2_combout ),
	.cout());
// synopsys translate_off
defparam \Mux59~2 .lut_mask = 16'hFC22;
defparam \Mux59~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X67_Y37_N23
dffeas \register[22][4] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\register~94_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~55_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\register[22][4]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \register[22][4] .is_wysiwyg = "true";
defparam \register[22][4] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X67_Y37_N22
cycloneive_lcell_comb \Mux59~3 (
// Equation(s):
// \Mux59~3_combout  = (Selector8 & ((\Mux59~2_combout  & ((\register[30][4]~q ))) # (!\Mux59~2_combout  & (\register[22][4]~q )))) # (!Selector8 & (\Mux59~2_combout ))

	.dataa(Selector8),
	.datab(\Mux59~2_combout ),
	.datac(\register[22][4]~q ),
	.datad(\register[30][4]~q ),
	.cin(gnd),
	.combout(\Mux59~3_combout ),
	.cout());
// synopsys translate_off
defparam \Mux59~3 .lut_mask = 16'hEC64;
defparam \Mux59~3 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X65_Y37_N28
cycloneive_lcell_comb \Mux59~4 (
// Equation(s):
// \Mux59~4_combout  = (Selector8 & (Selector7)) # (!Selector8 & ((Selector7 & ((\register[24][4]~q ))) # (!Selector7 & (\register[16][4]~q ))))

	.dataa(Selector8),
	.datab(Selector7),
	.datac(\register[16][4]~q ),
	.datad(\register[24][4]~q ),
	.cin(gnd),
	.combout(\Mux59~4_combout ),
	.cout());
// synopsys translate_off
defparam \Mux59~4 .lut_mask = 16'hDC98;
defparam \Mux59~4 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X66_Y33_N30
cycloneive_lcell_comb \Mux59~5 (
// Equation(s):
// \Mux59~5_combout  = (Selector8 & ((\Mux59~4_combout  & (\register[28][4]~q )) # (!\Mux59~4_combout  & ((\register[20][4]~q ))))) # (!Selector8 & (((\Mux59~4_combout ))))

	.dataa(\register[28][4]~q ),
	.datab(\register[20][4]~q ),
	.datac(Selector8),
	.datad(\Mux59~4_combout ),
	.cin(gnd),
	.combout(\Mux59~5_combout ),
	.cout());
// synopsys translate_off
defparam \Mux59~5 .lut_mask = 16'hAFC0;
defparam \Mux59~5 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y41_N6
cycloneive_lcell_comb \Mux59~6 (
// Equation(s):
// \Mux59~6_combout  = (Selector10 & (((Selector91)))) # (!Selector10 & ((Selector91 & (\Mux59~3_combout )) # (!Selector91 & ((\Mux59~5_combout )))))

	.dataa(Selector10),
	.datab(\Mux59~3_combout ),
	.datac(Selector91),
	.datad(\Mux59~5_combout ),
	.cin(gnd),
	.combout(\Mux59~6_combout ),
	.cout());
// synopsys translate_off
defparam \Mux59~6 .lut_mask = 16'hE5E0;
defparam \Mux59~6 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X67_Y31_N4
cycloneive_lcell_comb \Mux59~12 (
// Equation(s):
// \Mux59~12_combout  = (Selector10 & ((Selector91) # ((\register[5][4]~q )))) # (!Selector10 & (!Selector91 & ((\register[4][4]~q ))))

	.dataa(Selector10),
	.datab(Selector91),
	.datac(\register[5][4]~q ),
	.datad(\register[4][4]~q ),
	.cin(gnd),
	.combout(\Mux59~12_combout ),
	.cout());
// synopsys translate_off
defparam \Mux59~12 .lut_mask = 16'hB9A8;
defparam \Mux59~12 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X66_Y31_N10
cycloneive_lcell_comb \Mux59~13 (
// Equation(s):
// \Mux59~13_combout  = (Selector91 & ((\Mux59~12_combout  & ((\register[7][4]~q ))) # (!\Mux59~12_combout  & (\register[6][4]~q )))) # (!Selector91 & (((\Mux59~12_combout ))))

	.dataa(Selector91),
	.datab(\register[6][4]~q ),
	.datac(\register[7][4]~q ),
	.datad(\Mux59~12_combout ),
	.cin(gnd),
	.combout(\Mux59~13_combout ),
	.cout());
// synopsys translate_off
defparam \Mux59~13 .lut_mask = 16'hF588;
defparam \Mux59~13 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X67_Y34_N31
dffeas \register[2][4] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\register~94_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~50_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\register[2][4]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \register[2][4] .is_wysiwyg = "true";
defparam \register[2][4] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X67_Y34_N30
cycloneive_lcell_comb \Mux59~15 (
// Equation(s):
// \Mux59~15_combout  = (\Mux59~14_combout ) # ((!Selector10 & (\register[2][4]~q  & Selector91)))

	.dataa(\Mux59~14_combout ),
	.datab(Selector10),
	.datac(\register[2][4]~q ),
	.datad(Selector91),
	.cin(gnd),
	.combout(\Mux59~15_combout ),
	.cout());
// synopsys translate_off
defparam \Mux59~15 .lut_mask = 16'hBAAA;
defparam \Mux59~15 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y41_N10
cycloneive_lcell_comb \Mux59~16 (
// Equation(s):
// \Mux59~16_combout  = (Selector7 & (Selector8)) # (!Selector7 & ((Selector8 & (\Mux59~13_combout )) # (!Selector8 & ((\Mux59~15_combout )))))

	.dataa(Selector7),
	.datab(Selector8),
	.datac(\Mux59~13_combout ),
	.datad(\Mux59~15_combout ),
	.cin(gnd),
	.combout(\Mux59~16_combout ),
	.cout());
// synopsys translate_off
defparam \Mux59~16 .lut_mask = 16'hD9C8;
defparam \Mux59~16 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y33_N2
cycloneive_lcell_comb \Mux59~17 (
// Equation(s):
// \Mux59~17_combout  = (Selector10 & ((\register[13][4]~q ) # ((Selector91)))) # (!Selector10 & (((\register[12][4]~q  & !Selector91))))

	.dataa(\register[13][4]~q ),
	.datab(Selector10),
	.datac(\register[12][4]~q ),
	.datad(Selector91),
	.cin(gnd),
	.combout(\Mux59~17_combout ),
	.cout());
// synopsys translate_off
defparam \Mux59~17 .lut_mask = 16'hCCB8;
defparam \Mux59~17 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y34_N22
cycloneive_lcell_comb \Mux59~18 (
// Equation(s):
// \Mux59~18_combout  = (Selector91 & ((\Mux59~17_combout  & (\register[15][4]~q )) # (!\Mux59~17_combout  & ((\register[14][4]~q ))))) # (!Selector91 & (((\Mux59~17_combout ))))

	.dataa(\register[15][4]~q ),
	.datab(Selector91),
	.datac(\register[14][4]~q ),
	.datad(\Mux59~17_combout ),
	.cin(gnd),
	.combout(\Mux59~18_combout ),
	.cout());
// synopsys translate_off
defparam \Mux59~18 .lut_mask = 16'hBBC0;
defparam \Mux59~18 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X67_Y38_N8
cycloneive_lcell_comb \Mux59~10 (
// Equation(s):
// \Mux59~10_combout  = (Selector10 & (((Selector91)))) # (!Selector10 & ((Selector91 & ((\register[10][4]~q ))) # (!Selector91 & (\register[8][4]~q ))))

	.dataa(Selector10),
	.datab(\register[8][4]~q ),
	.datac(\register[10][4]~q ),
	.datad(Selector91),
	.cin(gnd),
	.combout(\Mux59~10_combout ),
	.cout());
// synopsys translate_off
defparam \Mux59~10 .lut_mask = 16'hFA44;
defparam \Mux59~10 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X63_Y34_N26
cycloneive_lcell_comb \Mux59~11 (
// Equation(s):
// \Mux59~11_combout  = (Selector10 & ((\Mux59~10_combout  & (\register[11][4]~q )) # (!\Mux59~10_combout  & ((\register[9][4]~q ))))) # (!Selector10 & (((\Mux59~10_combout ))))

	.dataa(\register[11][4]~q ),
	.datab(Selector10),
	.datac(\register[9][4]~q ),
	.datad(\Mux59~10_combout ),
	.cin(gnd),
	.combout(\Mux59~11_combout ),
	.cout());
// synopsys translate_off
defparam \Mux59~11 .lut_mask = 16'hBBC0;
defparam \Mux59~11 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y35_N2
cycloneive_lcell_comb \Mux0~7 (
// Equation(s):
// \Mux0~7_combout  = (Selector3 & (((\register[23][31]~q ) # (Selector2)))) # (!Selector3 & (\register[19][31]~q  & ((!Selector2))))

	.dataa(\register[19][31]~q ),
	.datab(\register[23][31]~q ),
	.datac(Selector3),
	.datad(Selector2),
	.cin(gnd),
	.combout(\Mux0~7_combout ),
	.cout());
// synopsys translate_off
defparam \Mux0~7 .lut_mask = 16'hF0CA;
defparam \Mux0~7 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y33_N14
cycloneive_lcell_comb \Mux0~8 (
// Equation(s):
// \Mux0~8_combout  = (\Mux0~7_combout  & (((\register[31][31]~q ) # (!Selector2)))) # (!\Mux0~7_combout  & (\register[27][31]~q  & ((Selector2))))

	.dataa(\Mux0~7_combout ),
	.datab(\register[27][31]~q ),
	.datac(\register[31][31]~q ),
	.datad(Selector2),
	.cin(gnd),
	.combout(\Mux0~8_combout ),
	.cout());
// synopsys translate_off
defparam \Mux0~8 .lut_mask = 16'hE4AA;
defparam \Mux0~8 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X62_Y35_N17
dffeas \register[17][31] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\register~64_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~26_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\register[17][31]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \register[17][31] .is_wysiwyg = "true";
defparam \register[17][31] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X62_Y35_N16
cycloneive_lcell_comb \Mux0~0 (
// Equation(s):
// \Mux0~0_combout  = (Selector2 & (Selector3)) # (!Selector2 & ((Selector3 & ((\register[21][31]~q ))) # (!Selector3 & (\register[17][31]~q ))))

	.dataa(Selector2),
	.datab(Selector3),
	.datac(\register[17][31]~q ),
	.datad(\register[21][31]~q ),
	.cin(gnd),
	.combout(\Mux0~0_combout ),
	.cout());
// synopsys translate_off
defparam \Mux0~0 .lut_mask = 16'hDC98;
defparam \Mux0~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y37_N12
cycloneive_lcell_comb \Mux0~1 (
// Equation(s):
// \Mux0~1_combout  = (Selector2 & ((\Mux0~0_combout  & (\register[29][31]~q )) # (!\Mux0~0_combout  & ((\register[25][31]~q ))))) # (!Selector2 & (\Mux0~0_combout ))

	.dataa(Selector2),
	.datab(\Mux0~0_combout ),
	.datac(\register[29][31]~q ),
	.datad(\register[25][31]~q ),
	.cin(gnd),
	.combout(\Mux0~1_combout ),
	.cout());
// synopsys translate_off
defparam \Mux0~1 .lut_mask = 16'hE6C4;
defparam \Mux0~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X65_Y39_N9
dffeas \register[20][31] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\register~64_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~35_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\register[20][31]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \register[20][31] .is_wysiwyg = "true";
defparam \register[20][31] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X65_Y35_N16
cycloneive_lcell_comb \Mux0~4 (
// Equation(s):
// \Mux0~4_combout  = (Selector2 & (((\register[24][31]~q ) # (Selector3)))) # (!Selector2 & (\register[16][31]~q  & ((!Selector3))))

	.dataa(\register[16][31]~q ),
	.datab(Selector2),
	.datac(\register[24][31]~q ),
	.datad(Selector3),
	.cin(gnd),
	.combout(\Mux0~4_combout ),
	.cout());
// synopsys translate_off
defparam \Mux0~4 .lut_mask = 16'hCCE2;
defparam \Mux0~4 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X65_Y39_N8
cycloneive_lcell_comb \Mux0~5 (
// Equation(s):
// \Mux0~5_combout  = (Selector3 & ((\Mux0~4_combout  & (\register[28][31]~q )) # (!\Mux0~4_combout  & ((\register[20][31]~q ))))) # (!Selector3 & (((\Mux0~4_combout ))))

	.dataa(Selector3),
	.datab(\register[28][31]~q ),
	.datac(\register[20][31]~q ),
	.datad(\Mux0~4_combout ),
	.cin(gnd),
	.combout(\Mux0~5_combout ),
	.cout());
// synopsys translate_off
defparam \Mux0~5 .lut_mask = 16'hDDA0;
defparam \Mux0~5 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X69_Y35_N18
cycloneive_lcell_comb \Mux0~2 (
// Equation(s):
// \Mux0~2_combout  = (Selector2 & ((Selector3) # ((\register[26][31]~q )))) # (!Selector2 & (!Selector3 & (\register[18][31]~q )))

	.dataa(Selector2),
	.datab(Selector3),
	.datac(\register[18][31]~q ),
	.datad(\register[26][31]~q ),
	.cin(gnd),
	.combout(\Mux0~2_combout ),
	.cout());
// synopsys translate_off
defparam \Mux0~2 .lut_mask = 16'hBA98;
defparam \Mux0~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X69_Y39_N6
cycloneive_lcell_comb \Mux0~3 (
// Equation(s):
// \Mux0~3_combout  = (Selector3 & ((\Mux0~2_combout  & ((\register[30][31]~q ))) # (!\Mux0~2_combout  & (\register[22][31]~q )))) # (!Selector3 & (((\Mux0~2_combout ))))

	.dataa(Selector3),
	.datab(\register[22][31]~q ),
	.datac(\register[30][31]~q ),
	.datad(\Mux0~2_combout ),
	.cin(gnd),
	.combout(\Mux0~3_combout ),
	.cout());
// synopsys translate_off
defparam \Mux0~3 .lut_mask = 16'hF588;
defparam \Mux0~3 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y33_N6
cycloneive_lcell_comb \Mux0~6 (
// Equation(s):
// \Mux0~6_combout  = (Selector41 & ((Selector5) # ((\Mux0~3_combout )))) # (!Selector41 & (!Selector5 & (\Mux0~5_combout )))

	.dataa(Selector41),
	.datab(Selector5),
	.datac(\Mux0~5_combout ),
	.datad(\Mux0~3_combout ),
	.cin(gnd),
	.combout(\Mux0~6_combout ),
	.cout());
// synopsys translate_off
defparam \Mux0~6 .lut_mask = 16'hBA98;
defparam \Mux0~6 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X69_Y31_N23
dffeas \register[4][31] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\register~64_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~60_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\register[4][31]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \register[4][31] .is_wysiwyg = "true";
defparam \register[4][31] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X69_Y31_N22
cycloneive_lcell_comb \Mux0~12 (
// Equation(s):
// \Mux0~12_combout  = (Selector5 & ((Selector41) # ((\register[5][31]~q )))) # (!Selector5 & (!Selector41 & (\register[4][31]~q )))

	.dataa(Selector5),
	.datab(Selector41),
	.datac(\register[4][31]~q ),
	.datad(\register[5][31]~q ),
	.cin(gnd),
	.combout(\Mux0~12_combout ),
	.cout());
// synopsys translate_off
defparam \Mux0~12 .lut_mask = 16'hBA98;
defparam \Mux0~12 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X68_Y31_N26
cycloneive_lcell_comb \Mux0~13 (
// Equation(s):
// \Mux0~13_combout  = (Selector41 & ((\Mux0~12_combout  & ((\register[7][31]~q ))) # (!\Mux0~12_combout  & (\register[6][31]~q )))) # (!Selector41 & (((\Mux0~12_combout ))))

	.dataa(Selector41),
	.datab(\register[6][31]~q ),
	.datac(\register[7][31]~q ),
	.datad(\Mux0~12_combout ),
	.cin(gnd),
	.combout(\Mux0~13_combout ),
	.cout());
// synopsys translate_off
defparam \Mux0~13 .lut_mask = 16'hF588;
defparam \Mux0~13 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X65_Y33_N8
cycloneive_lcell_comb \Mux0~14 (
// Equation(s):
// \Mux0~14_combout  = (plif_ifidinstr_l_22 & ((Selector4 & (\register[3][31]~q )) # (!Selector4 & ((\register[1][31]~q ))))) # (!plif_ifidinstr_l_22 & (((\register[1][31]~q ))))

	.dataa(plif_ifidinstr_l_22),
	.datab(Selector4),
	.datac(\register[3][31]~q ),
	.datad(\register[1][31]~q ),
	.cin(gnd),
	.combout(\Mux0~14_combout ),
	.cout());
// synopsys translate_off
defparam \Mux0~14 .lut_mask = 16'hF780;
defparam \Mux0~14 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X67_Y34_N4
cycloneive_lcell_comb \Mux0~15 (
// Equation(s):
// \Mux0~15_combout  = (Selector5 & (((\Mux0~14_combout )))) # (!Selector5 & (Selector41 & (\register[2][31]~q )))

	.dataa(Selector41),
	.datab(Selector5),
	.datac(\register[2][31]~q ),
	.datad(\Mux0~14_combout ),
	.cin(gnd),
	.combout(\Mux0~15_combout ),
	.cout());
// synopsys translate_off
defparam \Mux0~15 .lut_mask = 16'hEC20;
defparam \Mux0~15 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y33_N10
cycloneive_lcell_comb \Mux0~16 (
// Equation(s):
// \Mux0~16_combout  = (Selector3 & ((Selector2) # ((\Mux0~13_combout )))) # (!Selector3 & (!Selector2 & ((\Mux0~15_combout ))))

	.dataa(Selector3),
	.datab(Selector2),
	.datac(\Mux0~13_combout ),
	.datad(\Mux0~15_combout ),
	.cin(gnd),
	.combout(\Mux0~16_combout ),
	.cout());
// synopsys translate_off
defparam \Mux0~16 .lut_mask = 16'hB9A8;
defparam \Mux0~16 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X67_Y34_N12
cycloneive_lcell_comb \register[11][31]~feeder (
// Equation(s):
// \register[11][31]~feeder_combout  = \register~64_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(\register~64_combout ),
	.datad(gnd),
	.cin(gnd),
	.combout(\register[11][31]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \register[11][31]~feeder .lut_mask = 16'hF0F0;
defparam \register[11][31]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X67_Y34_N13
dffeas \register[11][31] (
	.clk(!CLK),
	.d(\register[11][31]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~47_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\register[11][31]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \register[11][31] .is_wysiwyg = "true";
defparam \register[11][31] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X62_Y41_N16
cycloneive_lcell_comb \Mux0~10 (
// Equation(s):
// \Mux0~10_combout  = (Selector41 & (((\register[10][31]~q ) # (Selector5)))) # (!Selector41 & (\register[8][31]~q  & ((!Selector5))))

	.dataa(\register[8][31]~q ),
	.datab(Selector41),
	.datac(\register[10][31]~q ),
	.datad(Selector5),
	.cin(gnd),
	.combout(\Mux0~10_combout ),
	.cout());
// synopsys translate_off
defparam \Mux0~10 .lut_mask = 16'hCCE2;
defparam \Mux0~10 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X66_Y38_N28
cycloneive_lcell_comb \Mux0~11 (
// Equation(s):
// \Mux0~11_combout  = (Selector5 & ((\Mux0~10_combout  & (\register[11][31]~q )) # (!\Mux0~10_combout  & ((\register[9][31]~q ))))) # (!Selector5 & (((\Mux0~10_combout ))))

	.dataa(Selector5),
	.datab(\register[11][31]~q ),
	.datac(\register[9][31]~q ),
	.datad(\Mux0~10_combout ),
	.cin(gnd),
	.combout(\Mux0~11_combout ),
	.cout());
// synopsys translate_off
defparam \Mux0~11 .lut_mask = 16'hDDA0;
defparam \Mux0~11 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X62_Y30_N31
dffeas \register[12][31] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\register~64_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~52_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\register[12][31]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \register[12][31] .is_wysiwyg = "true";
defparam \register[12][31] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X62_Y30_N30
cycloneive_lcell_comb \Mux0~17 (
// Equation(s):
// \Mux0~17_combout  = (Selector5 & ((Selector41) # ((\register[13][31]~q )))) # (!Selector5 & (!Selector41 & (\register[12][31]~q )))

	.dataa(Selector5),
	.datab(Selector41),
	.datac(\register[12][31]~q ),
	.datad(\register[13][31]~q ),
	.cin(gnd),
	.combout(\Mux0~17_combout ),
	.cout());
// synopsys translate_off
defparam \Mux0~17 .lut_mask = 16'hBA98;
defparam \Mux0~17 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y32_N20
cycloneive_lcell_comb \Mux0~18 (
// Equation(s):
// \Mux0~18_combout  = (\Mux0~17_combout  & ((\register[15][31]~q ) # ((!Selector41)))) # (!\Mux0~17_combout  & (((Selector41 & \register[14][31]~q ))))

	.dataa(\Mux0~17_combout ),
	.datab(\register[15][31]~q ),
	.datac(Selector41),
	.datad(\register[14][31]~q ),
	.cin(gnd),
	.combout(\Mux0~18_combout ),
	.cout());
// synopsys translate_off
defparam \Mux0~18 .lut_mask = 16'hDA8A;
defparam \Mux0~18 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y35_N4
cycloneive_lcell_comb \Mux2~0 (
// Equation(s):
// \Mux2~0_combout  = (Selector3 & ((\register[21][29]~q ) # ((Selector2)))) # (!Selector3 & (((\register[17][29]~q  & !Selector2))))

	.dataa(\register[21][29]~q ),
	.datab(Selector3),
	.datac(\register[17][29]~q ),
	.datad(Selector2),
	.cin(gnd),
	.combout(\Mux2~0_combout ),
	.cout());
// synopsys translate_off
defparam \Mux2~0 .lut_mask = 16'hCCB8;
defparam \Mux2~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y31_N14
cycloneive_lcell_comb \Mux2~1 (
// Equation(s):
// \Mux2~1_combout  = (Selector2 & ((\Mux2~0_combout  & (\register[29][29]~q )) # (!\Mux2~0_combout  & ((\register[25][29]~q ))))) # (!Selector2 & (((\Mux2~0_combout ))))

	.dataa(\register[29][29]~q ),
	.datab(Selector2),
	.datac(\Mux2~0_combout ),
	.datad(\register[25][29]~q ),
	.cin(gnd),
	.combout(\Mux2~1_combout ),
	.cout());
// synopsys translate_off
defparam \Mux2~1 .lut_mask = 16'hBCB0;
defparam \Mux2~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X68_Y35_N31
dffeas \register[30][29] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\register~66_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~56_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\register[30][29]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \register[30][29] .is_wysiwyg = "true";
defparam \register[30][29] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X68_Y35_N30
cycloneive_lcell_comb \Mux2~3 (
// Equation(s):
// \Mux2~3_combout  = (\Mux2~2_combout  & (((\register[30][29]~q ) # (!Selector3)))) # (!\Mux2~2_combout  & (\register[22][29]~q  & ((Selector3))))

	.dataa(\Mux2~2_combout ),
	.datab(\register[22][29]~q ),
	.datac(\register[30][29]~q ),
	.datad(Selector3),
	.cin(gnd),
	.combout(\Mux2~3_combout ),
	.cout());
// synopsys translate_off
defparam \Mux2~3 .lut_mask = 16'hE4AA;
defparam \Mux2~3 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X65_Y35_N9
dffeas \register[24][29] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\register~66_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~34_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\register[24][29]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \register[24][29] .is_wysiwyg = "true";
defparam \register[24][29] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X65_Y35_N8
cycloneive_lcell_comb \Mux2~4 (
// Equation(s):
// \Mux2~4_combout  = (Selector2 & (((\register[24][29]~q ) # (Selector3)))) # (!Selector2 & (\register[16][29]~q  & ((!Selector3))))

	.dataa(\register[16][29]~q ),
	.datab(Selector2),
	.datac(\register[24][29]~q ),
	.datad(Selector3),
	.cin(gnd),
	.combout(\Mux2~4_combout ),
	.cout());
// synopsys translate_off
defparam \Mux2~4 .lut_mask = 16'hCCE2;
defparam \Mux2~4 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X66_Y35_N20
cycloneive_lcell_comb \Mux2~5 (
// Equation(s):
// \Mux2~5_combout  = (Selector3 & ((\Mux2~4_combout  & ((\register[28][29]~q ))) # (!\Mux2~4_combout  & (\register[20][29]~q )))) # (!Selector3 & (((\Mux2~4_combout ))))

	.dataa(Selector3),
	.datab(\register[20][29]~q ),
	.datac(\register[28][29]~q ),
	.datad(\Mux2~4_combout ),
	.cin(gnd),
	.combout(\Mux2~5_combout ),
	.cout());
// synopsys translate_off
defparam \Mux2~5 .lut_mask = 16'hF588;
defparam \Mux2~5 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y33_N22
cycloneive_lcell_comb \Mux2~6 (
// Equation(s):
// \Mux2~6_combout  = (Selector41 & ((Selector5) # ((\Mux2~3_combout )))) # (!Selector41 & (!Selector5 & ((\Mux2~5_combout ))))

	.dataa(Selector41),
	.datab(Selector5),
	.datac(\Mux2~3_combout ),
	.datad(\Mux2~5_combout ),
	.cin(gnd),
	.combout(\Mux2~6_combout ),
	.cout());
// synopsys translate_off
defparam \Mux2~6 .lut_mask = 16'hB9A8;
defparam \Mux2~6 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y38_N8
cycloneive_lcell_comb \Mux2~7 (
// Equation(s):
// \Mux2~7_combout  = (Selector3 & ((Selector2) # ((\register[23][29]~q )))) # (!Selector3 & (!Selector2 & (\register[19][29]~q )))

	.dataa(Selector3),
	.datab(Selector2),
	.datac(\register[19][29]~q ),
	.datad(\register[23][29]~q ),
	.cin(gnd),
	.combout(\Mux2~7_combout ),
	.cout());
// synopsys translate_off
defparam \Mux2~7 .lut_mask = 16'hBA98;
defparam \Mux2~7 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y33_N12
cycloneive_lcell_comb \Mux2~8 (
// Equation(s):
// \Mux2~8_combout  = (\Mux2~7_combout  & (((\register[31][29]~q )) # (!Selector2))) # (!\Mux2~7_combout  & (Selector2 & ((\register[27][29]~q ))))

	.dataa(\Mux2~7_combout ),
	.datab(Selector2),
	.datac(\register[31][29]~q ),
	.datad(\register[27][29]~q ),
	.cin(gnd),
	.combout(\Mux2~8_combout ),
	.cout());
// synopsys translate_off
defparam \Mux2~8 .lut_mask = 16'hE6A2;
defparam \Mux2~8 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y36_N16
cycloneive_lcell_comb \Mux2~17 (
// Equation(s):
// \Mux2~17_combout  = (Selector41 & (((Selector5)))) # (!Selector41 & ((Selector5 & ((\register[13][29]~q ))) # (!Selector5 & (\register[12][29]~q ))))

	.dataa(\register[12][29]~q ),
	.datab(\register[13][29]~q ),
	.datac(Selector41),
	.datad(Selector5),
	.cin(gnd),
	.combout(\Mux2~17_combout ),
	.cout());
// synopsys translate_off
defparam \Mux2~17 .lut_mask = 16'hFC0A;
defparam \Mux2~17 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y36_N8
cycloneive_lcell_comb \Mux2~18 (
// Equation(s):
// \Mux2~18_combout  = (\Mux2~17_combout  & ((\register[15][29]~q ) # ((!Selector41)))) # (!\Mux2~17_combout  & (((\register[14][29]~q  & Selector41))))

	.dataa(\Mux2~17_combout ),
	.datab(\register[15][29]~q ),
	.datac(\register[14][29]~q ),
	.datad(Selector41),
	.cin(gnd),
	.combout(\Mux2~18_combout ),
	.cout());
// synopsys translate_off
defparam \Mux2~18 .lut_mask = 16'hD8AA;
defparam \Mux2~18 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X62_Y41_N31
dffeas \register[8][29] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\register~66_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~46_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\register[8][29]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \register[8][29] .is_wysiwyg = "true";
defparam \register[8][29] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X62_Y41_N30
cycloneive_lcell_comb \Mux2~10 (
// Equation(s):
// \Mux2~10_combout  = (Selector41 & ((\register[10][29]~q ) # ((Selector5)))) # (!Selector41 & (((\register[8][29]~q  & !Selector5))))

	.dataa(Selector41),
	.datab(\register[10][29]~q ),
	.datac(\register[8][29]~q ),
	.datad(Selector5),
	.cin(gnd),
	.combout(\Mux2~10_combout ),
	.cout());
// synopsys translate_off
defparam \Mux2~10 .lut_mask = 16'hAAD8;
defparam \Mux2~10 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X65_Y40_N0
cycloneive_lcell_comb \Mux2~11 (
// Equation(s):
// \Mux2~11_combout  = (Selector5 & ((\Mux2~10_combout  & (\register[11][29]~q )) # (!\Mux2~10_combout  & ((\register[9][29]~q ))))) # (!Selector5 & (((\Mux2~10_combout ))))

	.dataa(\register[11][29]~q ),
	.datab(Selector5),
	.datac(\register[9][29]~q ),
	.datad(\Mux2~10_combout ),
	.cin(gnd),
	.combout(\Mux2~11_combout ),
	.cout());
// synopsys translate_off
defparam \Mux2~11 .lut_mask = 16'hBBC0;
defparam \Mux2~11 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X69_Y33_N3
dffeas \register[1][29] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\register~66_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~49_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\register[1][29]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \register[1][29] .is_wysiwyg = "true";
defparam \register[1][29] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X69_Y33_N2
cycloneive_lcell_comb \Mux2~14 (
// Equation(s):
// \Mux2~14_combout  = (Selector5 & ((Selector41 & (\register[3][29]~q )) # (!Selector41 & ((\register[1][29]~q )))))

	.dataa(\register[3][29]~q ),
	.datab(Selector5),
	.datac(\register[1][29]~q ),
	.datad(Selector41),
	.cin(gnd),
	.combout(\Mux2~14_combout ),
	.cout());
// synopsys translate_off
defparam \Mux2~14 .lut_mask = 16'h88C0;
defparam \Mux2~14 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y33_N30
cycloneive_lcell_comb \Mux2~15 (
// Equation(s):
// \Mux2~15_combout  = (\Mux2~14_combout ) # ((Selector41 & (!Selector5 & \register[2][29]~q )))

	.dataa(Selector41),
	.datab(Selector5),
	.datac(\Mux2~14_combout ),
	.datad(\register[2][29]~q ),
	.cin(gnd),
	.combout(\Mux2~15_combout ),
	.cout());
// synopsys translate_off
defparam \Mux2~15 .lut_mask = 16'hF2F0;
defparam \Mux2~15 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X66_Y31_N26
cycloneive_lcell_comb \Mux2~13 (
// Equation(s):
// \Mux2~13_combout  = (\Mux2~12_combout  & (((\register[7][29]~q ) # (!Selector41)))) # (!\Mux2~12_combout  & (\register[6][29]~q  & ((Selector41))))

	.dataa(\Mux2~12_combout ),
	.datab(\register[6][29]~q ),
	.datac(\register[7][29]~q ),
	.datad(Selector41),
	.cin(gnd),
	.combout(\Mux2~13_combout ),
	.cout());
// synopsys translate_off
defparam \Mux2~13 .lut_mask = 16'hE4AA;
defparam \Mux2~13 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y33_N20
cycloneive_lcell_comb \Mux2~16 (
// Equation(s):
// \Mux2~16_combout  = (Selector3 & ((Selector2) # ((\Mux2~13_combout )))) # (!Selector3 & (!Selector2 & (\Mux2~15_combout )))

	.dataa(Selector3),
	.datab(Selector2),
	.datac(\Mux2~15_combout ),
	.datad(\Mux2~13_combout ),
	.cin(gnd),
	.combout(\Mux2~16_combout ),
	.cout());
// synopsys translate_off
defparam \Mux2~16 .lut_mask = 16'hBA98;
defparam \Mux2~16 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X65_Y35_N5
dffeas \register[24][30] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\register~65_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~34_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\register[24][30]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \register[24][30] .is_wysiwyg = "true";
defparam \register[24][30] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X65_Y39_N22
cycloneive_lcell_comb \Mux1~4 (
// Equation(s):
// \Mux1~4_combout  = (Selector2 & (Selector3)) # (!Selector2 & ((Selector3 & (\register[20][30]~q )) # (!Selector3 & ((\register[16][30]~q )))))

	.dataa(Selector2),
	.datab(Selector3),
	.datac(\register[20][30]~q ),
	.datad(\register[16][30]~q ),
	.cin(gnd),
	.combout(\Mux1~4_combout ),
	.cout());
// synopsys translate_off
defparam \Mux1~4 .lut_mask = 16'hD9C8;
defparam \Mux1~4 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X65_Y35_N4
cycloneive_lcell_comb \Mux1~5 (
// Equation(s):
// \Mux1~5_combout  = (Selector2 & ((\Mux1~4_combout  & (\register[28][30]~q )) # (!\Mux1~4_combout  & ((\register[24][30]~q ))))) # (!Selector2 & (((\Mux1~4_combout ))))

	.dataa(\register[28][30]~q ),
	.datab(Selector2),
	.datac(\register[24][30]~q ),
	.datad(\Mux1~4_combout ),
	.cin(gnd),
	.combout(\Mux1~5_combout ),
	.cout());
// synopsys translate_off
defparam \Mux1~5 .lut_mask = 16'hBBC0;
defparam \Mux1~5 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X69_Y35_N13
dffeas \register[22][30] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\register~65_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~55_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\register[22][30]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \register[22][30] .is_wysiwyg = "true";
defparam \register[22][30] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X69_Y35_N12
cycloneive_lcell_comb \Mux1~2 (
// Equation(s):
// \Mux1~2_combout  = (Selector3 & (((\register[22][30]~q ) # (Selector2)))) # (!Selector3 & (\register[18][30]~q  & ((!Selector2))))

	.dataa(\register[18][30]~q ),
	.datab(Selector3),
	.datac(\register[22][30]~q ),
	.datad(Selector2),
	.cin(gnd),
	.combout(\Mux1~2_combout ),
	.cout());
// synopsys translate_off
defparam \Mux1~2 .lut_mask = 16'hCCE2;
defparam \Mux1~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X68_Y35_N15
dffeas \register[26][30] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\register~65_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~54_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\register[26][30]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \register[26][30] .is_wysiwyg = "true";
defparam \register[26][30] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X68_Y35_N14
cycloneive_lcell_comb \Mux1~3 (
// Equation(s):
// \Mux1~3_combout  = (Selector2 & ((\Mux1~2_combout  & ((\register[30][30]~q ))) # (!\Mux1~2_combout  & (\register[26][30]~q )))) # (!Selector2 & (\Mux1~2_combout ))

	.dataa(Selector2),
	.datab(\Mux1~2_combout ),
	.datac(\register[26][30]~q ),
	.datad(\register[30][30]~q ),
	.cin(gnd),
	.combout(\Mux1~3_combout ),
	.cout());
// synopsys translate_off
defparam \Mux1~3 .lut_mask = 16'hEC64;
defparam \Mux1~3 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X65_Y35_N24
cycloneive_lcell_comb \Mux1~6 (
// Equation(s):
// \Mux1~6_combout  = (Selector5 & (((Selector41)))) # (!Selector5 & ((Selector41 & ((\Mux1~3_combout ))) # (!Selector41 & (\Mux1~5_combout ))))

	.dataa(Selector5),
	.datab(\Mux1~5_combout ),
	.datac(Selector41),
	.datad(\Mux1~3_combout ),
	.cin(gnd),
	.combout(\Mux1~6_combout ),
	.cout());
// synopsys translate_off
defparam \Mux1~6 .lut_mask = 16'hF4A4;
defparam \Mux1~6 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X62_Y35_N15
dffeas \register[17][30] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\register~65_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~26_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\register[17][30]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \register[17][30] .is_wysiwyg = "true";
defparam \register[17][30] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X62_Y35_N14
cycloneive_lcell_comb \Mux1~0 (
// Equation(s):
// \Mux1~0_combout  = (Selector2 & ((Selector3) # ((\register[25][30]~q )))) # (!Selector2 & (!Selector3 & (\register[17][30]~q )))

	.dataa(Selector2),
	.datab(Selector3),
	.datac(\register[17][30]~q ),
	.datad(\register[25][30]~q ),
	.cin(gnd),
	.combout(\Mux1~0_combout ),
	.cout());
// synopsys translate_off
defparam \Mux1~0 .lut_mask = 16'hBA98;
defparam \Mux1~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X63_Y33_N2
cycloneive_lcell_comb \Mux1~1 (
// Equation(s):
// \Mux1~1_combout  = (\Mux1~0_combout  & (((\register[29][30]~q ) # (!Selector3)))) # (!\Mux1~0_combout  & (\register[21][30]~q  & ((Selector3))))

	.dataa(\Mux1~0_combout ),
	.datab(\register[21][30]~q ),
	.datac(\register[29][30]~q ),
	.datad(Selector3),
	.cin(gnd),
	.combout(\Mux1~1_combout ),
	.cout());
// synopsys translate_off
defparam \Mux1~1 .lut_mask = 16'hE4AA;
defparam \Mux1~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y39_N6
cycloneive_lcell_comb \Mux1~7 (
// Equation(s):
// \Mux1~7_combout  = (Selector3 & (((Selector2)))) # (!Selector3 & ((Selector2 & ((\register[27][30]~q ))) # (!Selector2 & (\register[19][30]~q ))))

	.dataa(Selector3),
	.datab(\register[19][30]~q ),
	.datac(\register[27][30]~q ),
	.datad(Selector2),
	.cin(gnd),
	.combout(\Mux1~7_combout ),
	.cout());
// synopsys translate_off
defparam \Mux1~7 .lut_mask = 16'hFA44;
defparam \Mux1~7 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y39_N16
cycloneive_lcell_comb \Mux1~8 (
// Equation(s):
// \Mux1~8_combout  = (Selector3 & ((\Mux1~7_combout  & ((\register[31][30]~q ))) # (!\Mux1~7_combout  & (\register[23][30]~q )))) # (!Selector3 & (((\Mux1~7_combout ))))

	.dataa(Selector3),
	.datab(\register[23][30]~q ),
	.datac(\register[31][30]~q ),
	.datad(\Mux1~7_combout ),
	.cin(gnd),
	.combout(\Mux1~8_combout ),
	.cout());
// synopsys translate_off
defparam \Mux1~8 .lut_mask = 16'hF588;
defparam \Mux1~8 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X69_Y31_N11
dffeas \register[4][30] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\register~65_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~60_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\register[4][30]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \register[4][30] .is_wysiwyg = "true";
defparam \register[4][30] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X69_Y31_N10
cycloneive_lcell_comb \Mux1~10 (
// Equation(s):
// \Mux1~10_combout  = (Selector5 & ((\register[5][30]~q ) # ((Selector41)))) # (!Selector5 & (((\register[4][30]~q  & !Selector41))))

	.dataa(Selector5),
	.datab(\register[5][30]~q ),
	.datac(\register[4][30]~q ),
	.datad(Selector41),
	.cin(gnd),
	.combout(\Mux1~10_combout ),
	.cout());
// synopsys translate_off
defparam \Mux1~10 .lut_mask = 16'hAAD8;
defparam \Mux1~10 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X68_Y31_N20
cycloneive_lcell_comb \Mux1~11 (
// Equation(s):
// \Mux1~11_combout  = (Selector41 & ((\Mux1~10_combout  & ((\register[7][30]~q ))) # (!\Mux1~10_combout  & (\register[6][30]~q )))) # (!Selector41 & (\Mux1~10_combout ))

	.dataa(Selector41),
	.datab(\Mux1~10_combout ),
	.datac(\register[6][30]~q ),
	.datad(\register[7][30]~q ),
	.cin(gnd),
	.combout(\Mux1~11_combout ),
	.cout());
// synopsys translate_off
defparam \Mux1~11 .lut_mask = 16'hEC64;
defparam \Mux1~11 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y30_N8
cycloneive_lcell_comb \Mux1~17 (
// Equation(s):
// \Mux1~17_combout  = (Selector5 & ((Selector41) # ((\register[13][30]~q )))) # (!Selector5 & (!Selector41 & ((\register[12][30]~q ))))

	.dataa(Selector5),
	.datab(Selector41),
	.datac(\register[13][30]~q ),
	.datad(\register[12][30]~q ),
	.cin(gnd),
	.combout(\Mux1~17_combout ),
	.cout());
// synopsys translate_off
defparam \Mux1~17 .lut_mask = 16'hB9A8;
defparam \Mux1~17 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y32_N2
cycloneive_lcell_comb \Mux1~18 (
// Equation(s):
// \Mux1~18_combout  = (Selector41 & ((\Mux1~17_combout  & (\register[15][30]~q )) # (!\Mux1~17_combout  & ((\register[14][30]~q ))))) # (!Selector41 & (((\Mux1~17_combout ))))

	.dataa(\register[15][30]~q ),
	.datab(Selector41),
	.datac(\register[14][30]~q ),
	.datad(\Mux1~17_combout ),
	.cin(gnd),
	.combout(\Mux1~18_combout ),
	.cout());
// synopsys translate_off
defparam \Mux1~18 .lut_mask = 16'hBBC0;
defparam \Mux1~18 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X65_Y33_N16
cycloneive_lcell_comb \Mux1~14 (
// Equation(s):
// \Mux1~14_combout  = (Selector4 & ((plif_ifidinstr_l_22 & ((\register[3][30]~q ))) # (!plif_ifidinstr_l_22 & (\register[1][30]~q )))) # (!Selector4 & (\register[1][30]~q ))

	.dataa(\register[1][30]~q ),
	.datab(Selector4),
	.datac(\register[3][30]~q ),
	.datad(plif_ifidinstr_l_22),
	.cin(gnd),
	.combout(\Mux1~14_combout ),
	.cout());
// synopsys translate_off
defparam \Mux1~14 .lut_mask = 16'hE2AA;
defparam \Mux1~14 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X66_Y34_N12
cycloneive_lcell_comb \Mux1~15 (
// Equation(s):
// \Mux1~15_combout  = (Selector5 & (((\Mux1~14_combout )))) # (!Selector5 & (Selector41 & (\register[2][30]~q )))

	.dataa(Selector41),
	.datab(Selector5),
	.datac(\register[2][30]~q ),
	.datad(\Mux1~14_combout ),
	.cin(gnd),
	.combout(\Mux1~15_combout ),
	.cout());
// synopsys translate_off
defparam \Mux1~15 .lut_mask = 16'hEC20;
defparam \Mux1~15 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y41_N8
cycloneive_lcell_comb \Mux1~12 (
// Equation(s):
// \Mux1~12_combout  = (Selector41 & (((\register[10][30]~q ) # (Selector5)))) # (!Selector41 & (\register[8][30]~q  & ((!Selector5))))

	.dataa(Selector41),
	.datab(\register[8][30]~q ),
	.datac(\register[10][30]~q ),
	.datad(Selector5),
	.cin(gnd),
	.combout(\Mux1~12_combout ),
	.cout());
// synopsys translate_off
defparam \Mux1~12 .lut_mask = 16'hAAE4;
defparam \Mux1~12 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X66_Y38_N24
cycloneive_lcell_comb \Mux1~13 (
// Equation(s):
// \Mux1~13_combout  = (\Mux1~12_combout  & (((\register[11][30]~q ) # (!Selector5)))) # (!\Mux1~12_combout  & (\register[9][30]~q  & ((Selector5))))

	.dataa(\register[9][30]~q ),
	.datab(\Mux1~12_combout ),
	.datac(\register[11][30]~q ),
	.datad(Selector5),
	.cin(gnd),
	.combout(\Mux1~13_combout ),
	.cout());
// synopsys translate_off
defparam \Mux1~13 .lut_mask = 16'hE2CC;
defparam \Mux1~13 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X65_Y37_N6
cycloneive_lcell_comb \Mux1~16 (
// Equation(s):
// \Mux1~16_combout  = (Selector3 & (Selector2)) # (!Selector3 & ((Selector2 & ((\Mux1~13_combout ))) # (!Selector2 & (\Mux1~15_combout ))))

	.dataa(Selector3),
	.datab(Selector2),
	.datac(\Mux1~15_combout ),
	.datad(\Mux1~13_combout ),
	.cin(gnd),
	.combout(\Mux1~16_combout ),
	.cout());
// synopsys translate_off
defparam \Mux1~16 .lut_mask = 16'hDC98;
defparam \Mux1~16 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y35_N26
cycloneive_lcell_comb \register[17][28]~feeder (
// Equation(s):
// \register[17][28]~feeder_combout  = \register~67_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(\register~67_combout ),
	.cin(gnd),
	.combout(\register[17][28]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \register[17][28]~feeder .lut_mask = 16'hFF00;
defparam \register[17][28]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X62_Y35_N27
dffeas \register[17][28] (
	.clk(!CLK),
	.d(\register[17][28]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~26_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\register[17][28]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \register[17][28] .is_wysiwyg = "true";
defparam \register[17][28] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X62_Y35_N30
cycloneive_lcell_comb \Mux3~0 (
// Equation(s):
// \Mux3~0_combout  = (Selector2 & ((Selector3) # ((\register[25][28]~q )))) # (!Selector2 & (!Selector3 & (\register[17][28]~q )))

	.dataa(Selector2),
	.datab(Selector3),
	.datac(\register[17][28]~q ),
	.datad(\register[25][28]~q ),
	.cin(gnd),
	.combout(\Mux3~0_combout ),
	.cout());
// synopsys translate_off
defparam \Mux3~0 .lut_mask = 16'hBA98;
defparam \Mux3~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X63_Y39_N30
cycloneive_lcell_comb \Mux3~1 (
// Equation(s):
// \Mux3~1_combout  = (Selector3 & ((\Mux3~0_combout  & (\register[29][28]~q )) # (!\Mux3~0_combout  & ((\register[21][28]~q ))))) # (!Selector3 & (((\Mux3~0_combout ))))

	.dataa(\register[29][28]~q ),
	.datab(Selector3),
	.datac(\register[21][28]~q ),
	.datad(\Mux3~0_combout ),
	.cin(gnd),
	.combout(\Mux3~1_combout ),
	.cout());
// synopsys translate_off
defparam \Mux3~1 .lut_mask = 16'hBBC0;
defparam \Mux3~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y35_N28
cycloneive_lcell_comb \Mux3~7 (
// Equation(s):
// \Mux3~7_combout  = (Selector2 & ((Selector3) # ((\register[27][28]~q )))) # (!Selector2 & (!Selector3 & (\register[19][28]~q )))

	.dataa(Selector2),
	.datab(Selector3),
	.datac(\register[19][28]~q ),
	.datad(\register[27][28]~q ),
	.cin(gnd),
	.combout(\Mux3~7_combout ),
	.cout());
// synopsys translate_off
defparam \Mux3~7 .lut_mask = 16'hBA98;
defparam \Mux3~7 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y35_N24
cycloneive_lcell_comb \Mux3~8 (
// Equation(s):
// \Mux3~8_combout  = (Selector3 & ((\Mux3~7_combout  & ((\register[31][28]~q ))) # (!\Mux3~7_combout  & (\register[23][28]~q )))) # (!Selector3 & (((\Mux3~7_combout ))))

	.dataa(\register[23][28]~q ),
	.datab(\register[31][28]~q ),
	.datac(Selector3),
	.datad(\Mux3~7_combout ),
	.cin(gnd),
	.combout(\Mux3~8_combout ),
	.cout());
// synopsys translate_off
defparam \Mux3~8 .lut_mask = 16'hCFA0;
defparam \Mux3~8 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X69_Y39_N2
cycloneive_lcell_comb \Mux3~2 (
// Equation(s):
// \Mux3~2_combout  = (Selector2 & (((Selector3)))) # (!Selector2 & ((Selector3 & (\register[22][28]~q )) # (!Selector3 & ((\register[18][28]~q )))))

	.dataa(\register[22][28]~q ),
	.datab(Selector2),
	.datac(\register[18][28]~q ),
	.datad(Selector3),
	.cin(gnd),
	.combout(\Mux3~2_combout ),
	.cout());
// synopsys translate_off
defparam \Mux3~2 .lut_mask = 16'hEE30;
defparam \Mux3~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X67_Y39_N26
cycloneive_lcell_comb \Mux3~3 (
// Equation(s):
// \Mux3~3_combout  = (\Mux3~2_combout  & ((\register[30][28]~q ) # ((!Selector2)))) # (!\Mux3~2_combout  & (((\register[26][28]~q  & Selector2))))

	.dataa(\register[30][28]~q ),
	.datab(\Mux3~2_combout ),
	.datac(\register[26][28]~q ),
	.datad(Selector2),
	.cin(gnd),
	.combout(\Mux3~3_combout ),
	.cout());
// synopsys translate_off
defparam \Mux3~3 .lut_mask = 16'hB8CC;
defparam \Mux3~3 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X65_Y39_N17
dffeas \register[16][28] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\register~67_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~36_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\register[16][28]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \register[16][28] .is_wysiwyg = "true";
defparam \register[16][28] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X65_Y39_N10
cycloneive_lcell_comb \Mux3~4 (
// Equation(s):
// \Mux3~4_combout  = (Selector2 & (((Selector3)))) # (!Selector2 & ((Selector3 & ((\register[20][28]~q ))) # (!Selector3 & (\register[16][28]~q ))))

	.dataa(Selector2),
	.datab(\register[16][28]~q ),
	.datac(\register[20][28]~q ),
	.datad(Selector3),
	.cin(gnd),
	.combout(\Mux3~4_combout ),
	.cout());
// synopsys translate_off
defparam \Mux3~4 .lut_mask = 16'hFA44;
defparam \Mux3~4 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X67_Y39_N8
cycloneive_lcell_comb \Mux3~5 (
// Equation(s):
// \Mux3~5_combout  = (Selector2 & ((\Mux3~4_combout  & ((\register[28][28]~q ))) # (!\Mux3~4_combout  & (\register[24][28]~q )))) # (!Selector2 & (((\Mux3~4_combout ))))

	.dataa(\register[24][28]~q ),
	.datab(\register[28][28]~q ),
	.datac(Selector2),
	.datad(\Mux3~4_combout ),
	.cin(gnd),
	.combout(\Mux3~5_combout ),
	.cout());
// synopsys translate_off
defparam \Mux3~5 .lut_mask = 16'hCFA0;
defparam \Mux3~5 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X63_Y39_N12
cycloneive_lcell_comb \Mux3~6 (
// Equation(s):
// \Mux3~6_combout  = (Selector5 & (((Selector41)))) # (!Selector5 & ((Selector41 & (\Mux3~3_combout )) # (!Selector41 & ((\Mux3~5_combout )))))

	.dataa(\Mux3~3_combout ),
	.datab(Selector5),
	.datac(Selector41),
	.datad(\Mux3~5_combout ),
	.cin(gnd),
	.combout(\Mux3~6_combout ),
	.cout());
// synopsys translate_off
defparam \Mux3~6 .lut_mask = 16'hE3E0;
defparam \Mux3~6 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y41_N2
cycloneive_lcell_comb \Mux3~12 (
// Equation(s):
// \Mux3~12_combout  = (Selector41 & ((\register[10][28]~q ) # ((Selector5)))) # (!Selector41 & (((\register[8][28]~q  & !Selector5))))

	.dataa(Selector41),
	.datab(\register[10][28]~q ),
	.datac(\register[8][28]~q ),
	.datad(Selector5),
	.cin(gnd),
	.combout(\Mux3~12_combout ),
	.cout());
// synopsys translate_off
defparam \Mux3~12 .lut_mask = 16'hAAD8;
defparam \Mux3~12 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X65_Y40_N18
cycloneive_lcell_comb \Mux3~13 (
// Equation(s):
// \Mux3~13_combout  = (Selector5 & ((\Mux3~12_combout  & ((\register[11][28]~q ))) # (!\Mux3~12_combout  & (\register[9][28]~q )))) # (!Selector5 & (((\Mux3~12_combout ))))

	.dataa(Selector5),
	.datab(\register[9][28]~q ),
	.datac(\register[11][28]~q ),
	.datad(\Mux3~12_combout ),
	.cin(gnd),
	.combout(\Mux3~13_combout ),
	.cout());
// synopsys translate_off
defparam \Mux3~13 .lut_mask = 16'hF588;
defparam \Mux3~13 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X63_Y39_N24
cycloneive_lcell_comb \Mux3~15 (
// Equation(s):
// \Mux3~15_combout  = (\Mux3~14_combout ) # ((!Selector5 & (Selector41 & \register[2][28]~q )))

	.dataa(\Mux3~14_combout ),
	.datab(Selector5),
	.datac(Selector41),
	.datad(\register[2][28]~q ),
	.cin(gnd),
	.combout(\Mux3~15_combout ),
	.cout());
// synopsys translate_off
defparam \Mux3~15 .lut_mask = 16'hBAAA;
defparam \Mux3~15 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X63_Y39_N10
cycloneive_lcell_comb \Mux3~16 (
// Equation(s):
// \Mux3~16_combout  = (Selector2 & ((Selector3) # ((\Mux3~13_combout )))) # (!Selector2 & (!Selector3 & ((\Mux3~15_combout ))))

	.dataa(Selector2),
	.datab(Selector3),
	.datac(\Mux3~13_combout ),
	.datad(\Mux3~15_combout ),
	.cin(gnd),
	.combout(\Mux3~16_combout ),
	.cout());
// synopsys translate_off
defparam \Mux3~16 .lut_mask = 16'hB9A8;
defparam \Mux3~16 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X59_Y36_N15
dffeas \register[13][28] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\register~67_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~62_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\register[13][28]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \register[13][28] .is_wysiwyg = "true";
defparam \register[13][28] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X59_Y36_N14
cycloneive_lcell_comb \Mux3~17 (
// Equation(s):
// \Mux3~17_combout  = (Selector41 & (Selector5)) # (!Selector41 & ((Selector5 & (\register[13][28]~q )) # (!Selector5 & ((\register[12][28]~q )))))

	.dataa(Selector41),
	.datab(Selector5),
	.datac(\register[13][28]~q ),
	.datad(\register[12][28]~q ),
	.cin(gnd),
	.combout(\Mux3~17_combout ),
	.cout());
// synopsys translate_off
defparam \Mux3~17 .lut_mask = 16'hD9C8;
defparam \Mux3~17 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X63_Y37_N30
cycloneive_lcell_comb \Mux3~18 (
// Equation(s):
// \Mux3~18_combout  = (Selector41 & ((\Mux3~17_combout  & (\register[15][28]~q )) # (!\Mux3~17_combout  & ((\register[14][28]~q ))))) # (!Selector41 & (((\Mux3~17_combout ))))

	.dataa(\register[15][28]~q ),
	.datab(\register[14][28]~q ),
	.datac(Selector41),
	.datad(\Mux3~17_combout ),
	.cin(gnd),
	.combout(\Mux3~18_combout ),
	.cout());
// synopsys translate_off
defparam \Mux3~18 .lut_mask = 16'hAFC0;
defparam \Mux3~18 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X66_Y31_N21
dffeas \register[6][28] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\register~67_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~58_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\register[6][28]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \register[6][28] .is_wysiwyg = "true";
defparam \register[6][28] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X69_Y31_N20
cycloneive_lcell_comb \Mux3~10 (
// Equation(s):
// \Mux3~10_combout  = (Selector5 & ((Selector41) # ((\register[5][28]~q )))) # (!Selector5 & (!Selector41 & ((\register[4][28]~q ))))

	.dataa(Selector5),
	.datab(Selector41),
	.datac(\register[5][28]~q ),
	.datad(\register[4][28]~q ),
	.cin(gnd),
	.combout(\Mux3~10_combout ),
	.cout());
// synopsys translate_off
defparam \Mux3~10 .lut_mask = 16'hB9A8;
defparam \Mux3~10 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X66_Y31_N20
cycloneive_lcell_comb \Mux3~11 (
// Equation(s):
// \Mux3~11_combout  = (Selector41 & ((\Mux3~10_combout  & (\register[7][28]~q )) # (!\Mux3~10_combout  & ((\register[6][28]~q ))))) # (!Selector41 & (((\Mux3~10_combout ))))

	.dataa(Selector41),
	.datab(\register[7][28]~q ),
	.datac(\register[6][28]~q ),
	.datad(\Mux3~10_combout ),
	.cin(gnd),
	.combout(\Mux3~11_combout ),
	.cout());
// synopsys translate_off
defparam \Mux3~11 .lut_mask = 16'hDDA0;
defparam \Mux3~11 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X60_Y38_N27
dffeas \register[19][27] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\register~68_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~39_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\register[19][27]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \register[19][27] .is_wysiwyg = "true";
defparam \register[19][27] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X60_Y38_N26
cycloneive_lcell_comb \Mux4~7 (
// Equation(s):
// \Mux4~7_combout  = (Selector3 & ((Selector2) # ((\register[23][27]~q )))) # (!Selector3 & (!Selector2 & (\register[19][27]~q )))

	.dataa(Selector3),
	.datab(Selector2),
	.datac(\register[19][27]~q ),
	.datad(\register[23][27]~q ),
	.cin(gnd),
	.combout(\Mux4~7_combout ),
	.cout());
// synopsys translate_off
defparam \Mux4~7 .lut_mask = 16'hBA98;
defparam \Mux4~7 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y39_N0
cycloneive_lcell_comb \Mux4~8 (
// Equation(s):
// \Mux4~8_combout  = (\Mux4~7_combout  & (((\register[31][27]~q ) # (!Selector2)))) # (!\Mux4~7_combout  & (\register[27][27]~q  & ((Selector2))))

	.dataa(\Mux4~7_combout ),
	.datab(\register[27][27]~q ),
	.datac(\register[31][27]~q ),
	.datad(Selector2),
	.cin(gnd),
	.combout(\Mux4~8_combout ),
	.cout());
// synopsys translate_off
defparam \Mux4~8 .lut_mask = 16'hE4AA;
defparam \Mux4~8 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y35_N22
cycloneive_lcell_comb \Mux4~0 (
// Equation(s):
// \Mux4~0_combout  = (Selector2 & (((Selector3)))) # (!Selector2 & ((Selector3 & (\register[21][27]~q )) # (!Selector3 & ((\register[17][27]~q )))))

	.dataa(\register[21][27]~q ),
	.datab(Selector2),
	.datac(Selector3),
	.datad(\register[17][27]~q ),
	.cin(gnd),
	.combout(\Mux4~0_combout ),
	.cout());
// synopsys translate_off
defparam \Mux4~0 .lut_mask = 16'hE3E0;
defparam \Mux4~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X63_Y39_N22
cycloneive_lcell_comb \Mux4~1 (
// Equation(s):
// \Mux4~1_combout  = (Selector2 & ((\Mux4~0_combout  & (\register[29][27]~q )) # (!\Mux4~0_combout  & ((\register[25][27]~q ))))) # (!Selector2 & (((\Mux4~0_combout ))))

	.dataa(Selector2),
	.datab(\register[29][27]~q ),
	.datac(\register[25][27]~q ),
	.datad(\Mux4~0_combout ),
	.cin(gnd),
	.combout(\Mux4~1_combout ),
	.cout());
// synopsys translate_off
defparam \Mux4~1 .lut_mask = 16'hDDA0;
defparam \Mux4~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X65_Y39_N24
cycloneive_lcell_comb \Mux4~4 (
// Equation(s):
// \Mux4~4_combout  = (Selector2 & ((Selector3) # ((\register[24][27]~q )))) # (!Selector2 & (!Selector3 & (\register[16][27]~q )))

	.dataa(Selector2),
	.datab(Selector3),
	.datac(\register[16][27]~q ),
	.datad(\register[24][27]~q ),
	.cin(gnd),
	.combout(\Mux4~4_combout ),
	.cout());
// synopsys translate_off
defparam \Mux4~4 .lut_mask = 16'hBA98;
defparam \Mux4~4 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X66_Y39_N18
cycloneive_lcell_comb \Mux4~5 (
// Equation(s):
// \Mux4~5_combout  = (Selector3 & ((\Mux4~4_combout  & (\register[28][27]~q )) # (!\Mux4~4_combout  & ((\register[20][27]~q ))))) # (!Selector3 & (((\Mux4~4_combout ))))

	.dataa(Selector3),
	.datab(\register[28][27]~q ),
	.datac(\register[20][27]~q ),
	.datad(\Mux4~4_combout ),
	.cin(gnd),
	.combout(\Mux4~5_combout ),
	.cout());
// synopsys translate_off
defparam \Mux4~5 .lut_mask = 16'hDDA0;
defparam \Mux4~5 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X68_Y35_N0
cycloneive_lcell_comb \Mux4~2 (
// Equation(s):
// \Mux4~2_combout  = (Selector2 & ((Selector3) # ((\register[26][27]~q )))) # (!Selector2 & (!Selector3 & ((\register[18][27]~q ))))

	.dataa(Selector2),
	.datab(Selector3),
	.datac(\register[26][27]~q ),
	.datad(\register[18][27]~q ),
	.cin(gnd),
	.combout(\Mux4~2_combout ),
	.cout());
// synopsys translate_off
defparam \Mux4~2 .lut_mask = 16'hB9A8;
defparam \Mux4~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X68_Y35_N18
cycloneive_lcell_comb \Mux4~3 (
// Equation(s):
// \Mux4~3_combout  = (Selector3 & ((\Mux4~2_combout  & ((\register[30][27]~q ))) # (!\Mux4~2_combout  & (\register[22][27]~q )))) # (!Selector3 & (((\Mux4~2_combout ))))

	.dataa(\register[22][27]~q ),
	.datab(Selector3),
	.datac(\register[30][27]~q ),
	.datad(\Mux4~2_combout ),
	.cin(gnd),
	.combout(\Mux4~3_combout ),
	.cout());
// synopsys translate_off
defparam \Mux4~3 .lut_mask = 16'hF388;
defparam \Mux4~3 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X63_Y39_N0
cycloneive_lcell_comb \Mux4~6 (
// Equation(s):
// \Mux4~6_combout  = (Selector5 & (((Selector41)))) # (!Selector5 & ((Selector41 & ((\Mux4~3_combout ))) # (!Selector41 & (\Mux4~5_combout ))))

	.dataa(\Mux4~5_combout ),
	.datab(Selector5),
	.datac(Selector41),
	.datad(\Mux4~3_combout ),
	.cin(gnd),
	.combout(\Mux4~6_combout ),
	.cout());
// synopsys translate_off
defparam \Mux4~6 .lut_mask = 16'hF2C2;
defparam \Mux4~6 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X69_Y31_N7
dffeas \register[4][27] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\register~68_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~60_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\register[4][27]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \register[4][27] .is_wysiwyg = "true";
defparam \register[4][27] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X69_Y31_N6
cycloneive_lcell_comb \Mux4~12 (
// Equation(s):
// \Mux4~12_combout  = (Selector5 & ((\register[5][27]~q ) # ((Selector41)))) # (!Selector5 & (((\register[4][27]~q  & !Selector41))))

	.dataa(Selector5),
	.datab(\register[5][27]~q ),
	.datac(\register[4][27]~q ),
	.datad(Selector41),
	.cin(gnd),
	.combout(\Mux4~12_combout ),
	.cout());
// synopsys translate_off
defparam \Mux4~12 .lut_mask = 16'hAAD8;
defparam \Mux4~12 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X68_Y31_N2
cycloneive_lcell_comb \Mux4~13 (
// Equation(s):
// \Mux4~13_combout  = (Selector41 & ((\Mux4~12_combout  & ((\register[7][27]~q ))) # (!\Mux4~12_combout  & (\register[6][27]~q )))) # (!Selector41 & (((\Mux4~12_combout ))))

	.dataa(Selector41),
	.datab(\register[6][27]~q ),
	.datac(\register[7][27]~q ),
	.datad(\Mux4~12_combout ),
	.cin(gnd),
	.combout(\Mux4~13_combout ),
	.cout());
// synopsys translate_off
defparam \Mux4~13 .lut_mask = 16'hF588;
defparam \Mux4~13 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X67_Y34_N9
dffeas \register[2][27] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\register~68_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~50_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\register[2][27]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \register[2][27] .is_wysiwyg = "true";
defparam \register[2][27] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X69_Y33_N0
cycloneive_lcell_comb \Mux4~14 (
// Equation(s):
// \Mux4~14_combout  = (plif_ifidinstr_l_22 & ((Selector4 & ((\register[3][27]~q ))) # (!Selector4 & (\register[1][27]~q )))) # (!plif_ifidinstr_l_22 & (\register[1][27]~q ))

	.dataa(\register[1][27]~q ),
	.datab(plif_ifidinstr_l_22),
	.datac(\register[3][27]~q ),
	.datad(Selector4),
	.cin(gnd),
	.combout(\Mux4~14_combout ),
	.cout());
// synopsys translate_off
defparam \Mux4~14 .lut_mask = 16'hE2AA;
defparam \Mux4~14 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X67_Y34_N8
cycloneive_lcell_comb \Mux4~15 (
// Equation(s):
// \Mux4~15_combout  = (Selector5 & (((\Mux4~14_combout )))) # (!Selector5 & (Selector41 & (\register[2][27]~q )))

	.dataa(Selector41),
	.datab(Selector5),
	.datac(\register[2][27]~q ),
	.datad(\Mux4~14_combout ),
	.cin(gnd),
	.combout(\Mux4~15_combout ),
	.cout());
// synopsys translate_off
defparam \Mux4~15 .lut_mask = 16'hEC20;
defparam \Mux4~15 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X63_Y39_N28
cycloneive_lcell_comb \Mux4~16 (
// Equation(s):
// \Mux4~16_combout  = (Selector2 & (Selector3)) # (!Selector2 & ((Selector3 & (\Mux4~13_combout )) # (!Selector3 & ((\Mux4~15_combout )))))

	.dataa(Selector2),
	.datab(Selector3),
	.datac(\Mux4~13_combout ),
	.datad(\Mux4~15_combout ),
	.cin(gnd),
	.combout(\Mux4~16_combout ),
	.cout());
// synopsys translate_off
defparam \Mux4~16 .lut_mask = 16'hD9C8;
defparam \Mux4~16 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y41_N10
cycloneive_lcell_comb \Mux4~10 (
// Equation(s):
// \Mux4~10_combout  = (Selector41 & ((Selector5) # ((\register[10][27]~q )))) # (!Selector41 & (!Selector5 & (\register[8][27]~q )))

	.dataa(Selector41),
	.datab(Selector5),
	.datac(\register[8][27]~q ),
	.datad(\register[10][27]~q ),
	.cin(gnd),
	.combout(\Mux4~10_combout ),
	.cout());
// synopsys translate_off
defparam \Mux4~10 .lut_mask = 16'hBA98;
defparam \Mux4~10 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X66_Y38_N22
cycloneive_lcell_comb \Mux4~11 (
// Equation(s):
// \Mux4~11_combout  = (\Mux4~10_combout  & ((\register[11][27]~q ) # ((!Selector5)))) # (!\Mux4~10_combout  & (((\register[9][27]~q  & Selector5))))

	.dataa(\Mux4~10_combout ),
	.datab(\register[11][27]~q ),
	.datac(\register[9][27]~q ),
	.datad(Selector5),
	.cin(gnd),
	.combout(\Mux4~11_combout ),
	.cout());
// synopsys translate_off
defparam \Mux4~11 .lut_mask = 16'hD8AA;
defparam \Mux4~11 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X62_Y30_N23
dffeas \register[12][27] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\register~68_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~52_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\register[12][27]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \register[12][27] .is_wysiwyg = "true";
defparam \register[12][27] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X62_Y30_N22
cycloneive_lcell_comb \Mux4~17 (
// Equation(s):
// \Mux4~17_combout  = (Selector5 & ((Selector41) # ((\register[13][27]~q )))) # (!Selector5 & (!Selector41 & (\register[12][27]~q )))

	.dataa(Selector5),
	.datab(Selector41),
	.datac(\register[12][27]~q ),
	.datad(\register[13][27]~q ),
	.cin(gnd),
	.combout(\Mux4~17_combout ),
	.cout());
// synopsys translate_off
defparam \Mux4~17 .lut_mask = 16'hBA98;
defparam \Mux4~17 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y32_N14
cycloneive_lcell_comb \Mux4~18 (
// Equation(s):
// \Mux4~18_combout  = (\Mux4~17_combout  & (((\register[15][27]~q )) # (!Selector41))) # (!\Mux4~17_combout  & (Selector41 & (\register[14][27]~q )))

	.dataa(\Mux4~17_combout ),
	.datab(Selector41),
	.datac(\register[14][27]~q ),
	.datad(\register[15][27]~q ),
	.cin(gnd),
	.combout(\Mux4~18_combout ),
	.cout());
// synopsys translate_off
defparam \Mux4~18 .lut_mask = 16'hEA62;
defparam \Mux4~18 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y35_N4
cycloneive_lcell_comb \Mux5~7 (
// Equation(s):
// \Mux5~7_combout  = (Selector3 & (((Selector2)))) # (!Selector3 & ((Selector2 & (\register[27][26]~q )) # (!Selector2 & ((\register[19][26]~q )))))

	.dataa(\register[27][26]~q ),
	.datab(Selector3),
	.datac(\register[19][26]~q ),
	.datad(Selector2),
	.cin(gnd),
	.combout(\Mux5~7_combout ),
	.cout());
// synopsys translate_off
defparam \Mux5~7 .lut_mask = 16'hEE30;
defparam \Mux5~7 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X63_Y32_N12
cycloneive_lcell_comb \Mux5~8 (
// Equation(s):
// \Mux5~8_combout  = (Selector3 & ((\Mux5~7_combout  & ((\register[31][26]~q ))) # (!\Mux5~7_combout  & (\register[23][26]~q )))) # (!Selector3 & (((\Mux5~7_combout ))))

	.dataa(\register[23][26]~q ),
	.datab(Selector3),
	.datac(\Mux5~7_combout ),
	.datad(\register[31][26]~q ),
	.cin(gnd),
	.combout(\Mux5~8_combout ),
	.cout());
// synopsys translate_off
defparam \Mux5~8 .lut_mask = 16'hF838;
defparam \Mux5~8 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y37_N24
cycloneive_lcell_comb \Mux5~0 (
// Equation(s):
// \Mux5~0_combout  = (Selector2 & ((\register[25][26]~q ) # ((Selector3)))) # (!Selector2 & (((\register[17][26]~q  & !Selector3))))

	.dataa(\register[25][26]~q ),
	.datab(Selector2),
	.datac(\register[17][26]~q ),
	.datad(Selector3),
	.cin(gnd),
	.combout(\Mux5~0_combout ),
	.cout());
// synopsys translate_off
defparam \Mux5~0 .lut_mask = 16'hCCB8;
defparam \Mux5~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X63_Y32_N8
cycloneive_lcell_comb \Mux5~1 (
// Equation(s):
// \Mux5~1_combout  = (Selector3 & ((\Mux5~0_combout  & ((\register[29][26]~q ))) # (!\Mux5~0_combout  & (\register[21][26]~q )))) # (!Selector3 & (((\Mux5~0_combout ))))

	.dataa(\register[21][26]~q ),
	.datab(\register[29][26]~q ),
	.datac(Selector3),
	.datad(\Mux5~0_combout ),
	.cin(gnd),
	.combout(\Mux5~1_combout ),
	.cout());
// synopsys translate_off
defparam \Mux5~1 .lut_mask = 16'hCFA0;
defparam \Mux5~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X69_Y35_N16
cycloneive_lcell_comb \Mux5~2 (
// Equation(s):
// \Mux5~2_combout  = (Selector2 & (((Selector3)))) # (!Selector2 & ((Selector3 & (\register[22][26]~q )) # (!Selector3 & ((\register[18][26]~q )))))

	.dataa(Selector2),
	.datab(\register[22][26]~q ),
	.datac(\register[18][26]~q ),
	.datad(Selector3),
	.cin(gnd),
	.combout(\Mux5~2_combout ),
	.cout());
// synopsys translate_off
defparam \Mux5~2 .lut_mask = 16'hEE50;
defparam \Mux5~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X68_Y34_N6
cycloneive_lcell_comb \Mux5~3 (
// Equation(s):
// \Mux5~3_combout  = (Selector2 & ((\Mux5~2_combout  & (\register[30][26]~q )) # (!\Mux5~2_combout  & ((\register[26][26]~q ))))) # (!Selector2 & (((\Mux5~2_combout ))))

	.dataa(Selector2),
	.datab(\register[30][26]~q ),
	.datac(\Mux5~2_combout ),
	.datad(\register[26][26]~q ),
	.cin(gnd),
	.combout(\Mux5~3_combout ),
	.cout());
// synopsys translate_off
defparam \Mux5~3 .lut_mask = 16'hDAD0;
defparam \Mux5~3 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X65_Y35_N13
dffeas \register[16][26] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\register~69_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~36_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\register[16][26]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \register[16][26] .is_wysiwyg = "true";
defparam \register[16][26] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X65_Y35_N12
cycloneive_lcell_comb \Mux5~4 (
// Equation(s):
// \Mux5~4_combout  = (Selector2 & (((Selector3)))) # (!Selector2 & ((Selector3 & (\register[20][26]~q )) # (!Selector3 & ((\register[16][26]~q )))))

	.dataa(\register[20][26]~q ),
	.datab(Selector2),
	.datac(\register[16][26]~q ),
	.datad(Selector3),
	.cin(gnd),
	.combout(\Mux5~4_combout ),
	.cout());
// synopsys translate_off
defparam \Mux5~4 .lut_mask = 16'hEE30;
defparam \Mux5~4 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X66_Y35_N22
cycloneive_lcell_comb \Mux5~5 (
// Equation(s):
// \Mux5~5_combout  = (Selector2 & ((\Mux5~4_combout  & (\register[28][26]~q )) # (!\Mux5~4_combout  & ((\register[24][26]~q ))))) # (!Selector2 & (((\Mux5~4_combout ))))

	.dataa(\register[28][26]~q ),
	.datab(\register[24][26]~q ),
	.datac(Selector2),
	.datad(\Mux5~4_combout ),
	.cin(gnd),
	.combout(\Mux5~5_combout ),
	.cout());
// synopsys translate_off
defparam \Mux5~5 .lut_mask = 16'hAFC0;
defparam \Mux5~5 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X63_Y32_N10
cycloneive_lcell_comb \Mux5~6 (
// Equation(s):
// \Mux5~6_combout  = (Selector5 & (((Selector41)))) # (!Selector5 & ((Selector41 & (\Mux5~3_combout )) # (!Selector41 & ((\Mux5~5_combout )))))

	.dataa(\Mux5~3_combout ),
	.datab(Selector5),
	.datac(Selector41),
	.datad(\Mux5~5_combout ),
	.cin(gnd),
	.combout(\Mux5~6_combout ),
	.cout());
// synopsys translate_off
defparam \Mux5~6 .lut_mask = 16'hE3E0;
defparam \Mux5~6 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y30_N18
cycloneive_lcell_comb \Mux5~17 (
// Equation(s):
// \Mux5~17_combout  = (Selector5 & ((\register[13][26]~q ) # ((Selector41)))) # (!Selector5 & (((\register[12][26]~q  & !Selector41))))

	.dataa(Selector5),
	.datab(\register[13][26]~q ),
	.datac(\register[12][26]~q ),
	.datad(Selector41),
	.cin(gnd),
	.combout(\Mux5~17_combout ),
	.cout());
// synopsys translate_off
defparam \Mux5~17 .lut_mask = 16'hAAD8;
defparam \Mux5~17 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y32_N0
cycloneive_lcell_comb \Mux5~18 (
// Equation(s):
// \Mux5~18_combout  = (Selector41 & ((\Mux5~17_combout  & ((\register[15][26]~q ))) # (!\Mux5~17_combout  & (\register[14][26]~q )))) # (!Selector41 & (((\Mux5~17_combout ))))

	.dataa(\register[14][26]~q ),
	.datab(Selector41),
	.datac(\register[15][26]~q ),
	.datad(\Mux5~17_combout ),
	.cin(gnd),
	.combout(\Mux5~18_combout ),
	.cout());
// synopsys translate_off
defparam \Mux5~18 .lut_mask = 16'hF388;
defparam \Mux5~18 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X69_Y31_N28
cycloneive_lcell_comb \Mux5~10 (
// Equation(s):
// \Mux5~10_combout  = (Selector41 & (((Selector5)))) # (!Selector41 & ((Selector5 & ((\register[5][26]~q ))) # (!Selector5 & (\register[4][26]~q ))))

	.dataa(\register[4][26]~q ),
	.datab(Selector41),
	.datac(\register[5][26]~q ),
	.datad(Selector5),
	.cin(gnd),
	.combout(\Mux5~10_combout ),
	.cout());
// synopsys translate_off
defparam \Mux5~10 .lut_mask = 16'hFC22;
defparam \Mux5~10 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X68_Y31_N0
cycloneive_lcell_comb \Mux5~11 (
// Equation(s):
// \Mux5~11_combout  = (Selector41 & ((\Mux5~10_combout  & (\register[7][26]~q )) # (!\Mux5~10_combout  & ((\register[6][26]~q ))))) # (!Selector41 & (((\Mux5~10_combout ))))

	.dataa(Selector41),
	.datab(\register[7][26]~q ),
	.datac(\register[6][26]~q ),
	.datad(\Mux5~10_combout ),
	.cin(gnd),
	.combout(\Mux5~11_combout ),
	.cout());
// synopsys translate_off
defparam \Mux5~11 .lut_mask = 16'hDDA0;
defparam \Mux5~11 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X66_Y34_N8
cycloneive_lcell_comb \register[2][26]~feeder (
// Equation(s):
// \register[2][26]~feeder_combout  = \register~69_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(\register~69_combout ),
	.cin(gnd),
	.combout(\register[2][26]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \register[2][26]~feeder .lut_mask = 16'hFF00;
defparam \register[2][26]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X66_Y34_N9
dffeas \register[2][26] (
	.clk(!CLK),
	.d(\register[2][26]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~50_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\register[2][26]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \register[2][26] .is_wysiwyg = "true";
defparam \register[2][26] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X69_Y33_N20
cycloneive_lcell_comb \Mux5~14 (
// Equation(s):
// \Mux5~14_combout  = (Selector5 & ((Selector41 & (\register[3][26]~q )) # (!Selector41 & ((\register[1][26]~q )))))

	.dataa(Selector41),
	.datab(Selector5),
	.datac(\register[3][26]~q ),
	.datad(\register[1][26]~q ),
	.cin(gnd),
	.combout(\Mux5~14_combout ),
	.cout());
// synopsys translate_off
defparam \Mux5~14 .lut_mask = 16'hC480;
defparam \Mux5~14 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X66_Y34_N6
cycloneive_lcell_comb \Mux5~15 (
// Equation(s):
// \Mux5~15_combout  = (\Mux5~14_combout ) # ((!Selector5 & (\register[2][26]~q  & Selector41)))

	.dataa(Selector5),
	.datab(\register[2][26]~q ),
	.datac(\Mux5~14_combout ),
	.datad(Selector41),
	.cin(gnd),
	.combout(\Mux5~15_combout ),
	.cout());
// synopsys translate_off
defparam \Mux5~15 .lut_mask = 16'hF4F0;
defparam \Mux5~15 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X66_Y40_N2
cycloneive_lcell_comb \Mux5~12 (
// Equation(s):
// \Mux5~12_combout  = (Selector41 & ((\register[10][26]~q ) # ((Selector5)))) # (!Selector41 & (((\register[8][26]~q  & !Selector5))))

	.dataa(\register[10][26]~q ),
	.datab(Selector41),
	.datac(\register[8][26]~q ),
	.datad(Selector5),
	.cin(gnd),
	.combout(\Mux5~12_combout ),
	.cout());
// synopsys translate_off
defparam \Mux5~12 .lut_mask = 16'hCCB8;
defparam \Mux5~12 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X63_Y34_N0
cycloneive_lcell_comb \Mux5~13 (
// Equation(s):
// \Mux5~13_combout  = (Selector5 & ((\Mux5~12_combout  & (\register[11][26]~q )) # (!\Mux5~12_combout  & ((\register[9][26]~q ))))) # (!Selector5 & (((\Mux5~12_combout ))))

	.dataa(\register[11][26]~q ),
	.datab(Selector5),
	.datac(\register[9][26]~q ),
	.datad(\Mux5~12_combout ),
	.cin(gnd),
	.combout(\Mux5~13_combout ),
	.cout());
// synopsys translate_off
defparam \Mux5~13 .lut_mask = 16'hBBC0;
defparam \Mux5~13 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X63_Y32_N28
cycloneive_lcell_comb \Mux5~16 (
// Equation(s):
// \Mux5~16_combout  = (Selector2 & (((Selector3) # (\Mux5~13_combout )))) # (!Selector2 & (\Mux5~15_combout  & (!Selector3)))

	.dataa(\Mux5~15_combout ),
	.datab(Selector2),
	.datac(Selector3),
	.datad(\Mux5~13_combout ),
	.cin(gnd),
	.combout(\Mux5~16_combout ),
	.cout());
// synopsys translate_off
defparam \Mux5~16 .lut_mask = 16'hCEC2;
defparam \Mux5~16 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y35_N12
cycloneive_lcell_comb \Mux6~0 (
// Equation(s):
// \Mux6~0_combout  = (Selector2 & (Selector3)) # (!Selector2 & ((Selector3 & ((\register[21][25]~q ))) # (!Selector3 & (\register[17][25]~q ))))

	.dataa(Selector2),
	.datab(Selector3),
	.datac(\register[17][25]~q ),
	.datad(\register[21][25]~q ),
	.cin(gnd),
	.combout(\Mux6~0_combout ),
	.cout());
// synopsys translate_off
defparam \Mux6~0 .lut_mask = 16'hDC98;
defparam \Mux6~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y31_N16
cycloneive_lcell_comb \Mux6~1 (
// Equation(s):
// \Mux6~1_combout  = (Selector2 & ((\Mux6~0_combout  & ((\register[29][25]~q ))) # (!\Mux6~0_combout  & (\register[25][25]~q )))) # (!Selector2 & (((\Mux6~0_combout ))))

	.dataa(\register[25][25]~q ),
	.datab(Selector2),
	.datac(\Mux6~0_combout ),
	.datad(\register[29][25]~q ),
	.cin(gnd),
	.combout(\Mux6~1_combout ),
	.cout());
// synopsys translate_off
defparam \Mux6~1 .lut_mask = 16'hF838;
defparam \Mux6~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y38_N14
cycloneive_lcell_comb \Mux6~7 (
// Equation(s):
// \Mux6~7_combout  = (Selector3 & ((Selector2) # ((\register[23][25]~q )))) # (!Selector3 & (!Selector2 & (\register[19][25]~q )))

	.dataa(Selector3),
	.datab(Selector2),
	.datac(\register[19][25]~q ),
	.datad(\register[23][25]~q ),
	.cin(gnd),
	.combout(\Mux6~7_combout ),
	.cout());
// synopsys translate_off
defparam \Mux6~7 .lut_mask = 16'hBA98;
defparam \Mux6~7 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X65_Y31_N30
cycloneive_lcell_comb \Mux6~8 (
// Equation(s):
// \Mux6~8_combout  = (Selector2 & ((\Mux6~7_combout  & ((\register[31][25]~q ))) # (!\Mux6~7_combout  & (\register[27][25]~q )))) # (!Selector2 & (((\Mux6~7_combout ))))

	.dataa(\register[27][25]~q ),
	.datab(\register[31][25]~q ),
	.datac(Selector2),
	.datad(\Mux6~7_combout ),
	.cin(gnd),
	.combout(\Mux6~8_combout ),
	.cout());
// synopsys translate_off
defparam \Mux6~8 .lut_mask = 16'hCFA0;
defparam \Mux6~8 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X69_Y35_N26
cycloneive_lcell_comb \Mux6~2 (
// Equation(s):
// \Mux6~2_combout  = (Selector2 & ((Selector3) # ((\register[26][25]~q )))) # (!Selector2 & (!Selector3 & (\register[18][25]~q )))

	.dataa(Selector2),
	.datab(Selector3),
	.datac(\register[18][25]~q ),
	.datad(\register[26][25]~q ),
	.cin(gnd),
	.combout(\Mux6~2_combout ),
	.cout());
// synopsys translate_off
defparam \Mux6~2 .lut_mask = 16'hBA98;
defparam \Mux6~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X65_Y31_N6
cycloneive_lcell_comb \Mux6~3 (
// Equation(s):
// \Mux6~3_combout  = (Selector3 & ((\Mux6~2_combout  & ((\register[30][25]~q ))) # (!\Mux6~2_combout  & (\register[22][25]~q )))) # (!Selector3 & (((\Mux6~2_combout ))))

	.dataa(Selector3),
	.datab(\register[22][25]~q ),
	.datac(\register[30][25]~q ),
	.datad(\Mux6~2_combout ),
	.cin(gnd),
	.combout(\Mux6~3_combout ),
	.cout());
// synopsys translate_off
defparam \Mux6~3 .lut_mask = 16'hF588;
defparam \Mux6~3 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X66_Y39_N7
dffeas \register[24][25] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\register~70_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~34_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\register[24][25]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \register[24][25] .is_wysiwyg = "true";
defparam \register[24][25] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X69_Y38_N26
cycloneive_lcell_comb \register[16][25]~feeder (
// Equation(s):
// \register[16][25]~feeder_combout  = \register~70_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(\register~70_combout ),
	.datad(gnd),
	.cin(gnd),
	.combout(\register[16][25]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \register[16][25]~feeder .lut_mask = 16'hF0F0;
defparam \register[16][25]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X69_Y38_N27
dffeas \register[16][25] (
	.clk(!CLK),
	.d(\register[16][25]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~36_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\register[16][25]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \register[16][25] .is_wysiwyg = "true";
defparam \register[16][25] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X66_Y39_N6
cycloneive_lcell_comb \Mux6~4 (
// Equation(s):
// \Mux6~4_combout  = (Selector3 & (Selector2)) # (!Selector3 & ((Selector2 & (\register[24][25]~q )) # (!Selector2 & ((\register[16][25]~q )))))

	.dataa(Selector3),
	.datab(Selector2),
	.datac(\register[24][25]~q ),
	.datad(\register[16][25]~q ),
	.cin(gnd),
	.combout(\Mux6~4_combout ),
	.cout());
// synopsys translate_off
defparam \Mux6~4 .lut_mask = 16'hD9C8;
defparam \Mux6~4 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X66_Y39_N16
cycloneive_lcell_comb \Mux6~5 (
// Equation(s):
// \Mux6~5_combout  = (Selector3 & ((\Mux6~4_combout  & ((\register[28][25]~q ))) # (!\Mux6~4_combout  & (\register[20][25]~q )))) # (!Selector3 & (((\Mux6~4_combout ))))

	.dataa(Selector3),
	.datab(\register[20][25]~q ),
	.datac(\register[28][25]~q ),
	.datad(\Mux6~4_combout ),
	.cin(gnd),
	.combout(\Mux6~5_combout ),
	.cout());
// synopsys translate_off
defparam \Mux6~5 .lut_mask = 16'hF588;
defparam \Mux6~5 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X65_Y31_N16
cycloneive_lcell_comb \Mux6~6 (
// Equation(s):
// \Mux6~6_combout  = (Selector5 & (((Selector41)))) # (!Selector5 & ((Selector41 & (\Mux6~3_combout )) # (!Selector41 & ((\Mux6~5_combout )))))

	.dataa(\Mux6~3_combout ),
	.datab(Selector5),
	.datac(Selector41),
	.datad(\Mux6~5_combout ),
	.cin(gnd),
	.combout(\Mux6~6_combout ),
	.cout());
// synopsys translate_off
defparam \Mux6~6 .lut_mask = 16'hE3E0;
defparam \Mux6~6 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X66_Y40_N28
cycloneive_lcell_comb \Mux6~10 (
// Equation(s):
// \Mux6~10_combout  = (Selector5 & (((Selector41)))) # (!Selector5 & ((Selector41 & ((\register[10][25]~q ))) # (!Selector41 & (\register[8][25]~q ))))

	.dataa(\register[8][25]~q ),
	.datab(Selector5),
	.datac(\register[10][25]~q ),
	.datad(Selector41),
	.cin(gnd),
	.combout(\Mux6~10_combout ),
	.cout());
// synopsys translate_off
defparam \Mux6~10 .lut_mask = 16'hFC22;
defparam \Mux6~10 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X65_Y40_N28
cycloneive_lcell_comb \Mux6~11 (
// Equation(s):
// \Mux6~11_combout  = (\Mux6~10_combout  & ((\register[11][25]~q ) # ((!Selector5)))) # (!\Mux6~10_combout  & (((\register[9][25]~q  & Selector5))))

	.dataa(\register[11][25]~q ),
	.datab(\Mux6~10_combout ),
	.datac(\register[9][25]~q ),
	.datad(Selector5),
	.cin(gnd),
	.combout(\Mux6~11_combout ),
	.cout());
// synopsys translate_off
defparam \Mux6~11 .lut_mask = 16'hB8CC;
defparam \Mux6~11 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X67_Y31_N27
dffeas \register[4][25] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\register~70_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~60_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\register[4][25]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \register[4][25] .is_wysiwyg = "true";
defparam \register[4][25] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X67_Y31_N26
cycloneive_lcell_comb \Mux6~12 (
// Equation(s):
// \Mux6~12_combout  = (Selector41 & (((Selector5)))) # (!Selector41 & ((Selector5 & (\register[5][25]~q )) # (!Selector5 & ((\register[4][25]~q )))))

	.dataa(Selector41),
	.datab(\register[5][25]~q ),
	.datac(\register[4][25]~q ),
	.datad(Selector5),
	.cin(gnd),
	.combout(\Mux6~12_combout ),
	.cout());
// synopsys translate_off
defparam \Mux6~12 .lut_mask = 16'hEE50;
defparam \Mux6~12 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X66_Y31_N12
cycloneive_lcell_comb \Mux6~13 (
// Equation(s):
// \Mux6~13_combout  = (Selector41 & ((\Mux6~12_combout  & ((\register[7][25]~q ))) # (!\Mux6~12_combout  & (\register[6][25]~q )))) # (!Selector41 & (((\Mux6~12_combout ))))

	.dataa(\register[6][25]~q ),
	.datab(Selector41),
	.datac(\register[7][25]~q ),
	.datad(\Mux6~12_combout ),
	.cin(gnd),
	.combout(\Mux6~13_combout ),
	.cout());
// synopsys translate_off
defparam \Mux6~13 .lut_mask = 16'hF388;
defparam \Mux6~13 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X65_Y31_N10
cycloneive_lcell_comb \Mux6~15 (
// Equation(s):
// \Mux6~15_combout  = (Selector5 & (\Mux6~14_combout )) # (!Selector5 & (((Selector41 & \register[2][25]~q ))))

	.dataa(\Mux6~14_combout ),
	.datab(Selector5),
	.datac(Selector41),
	.datad(\register[2][25]~q ),
	.cin(gnd),
	.combout(\Mux6~15_combout ),
	.cout());
// synopsys translate_off
defparam \Mux6~15 .lut_mask = 16'hB888;
defparam \Mux6~15 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X65_Y31_N28
cycloneive_lcell_comb \Mux6~16 (
// Equation(s):
// \Mux6~16_combout  = (Selector2 & (((Selector3)))) # (!Selector2 & ((Selector3 & (\Mux6~13_combout )) # (!Selector3 & ((\Mux6~15_combout )))))

	.dataa(Selector2),
	.datab(\Mux6~13_combout ),
	.datac(Selector3),
	.datad(\Mux6~15_combout ),
	.cin(gnd),
	.combout(\Mux6~16_combout ),
	.cout());
// synopsys translate_off
defparam \Mux6~16 .lut_mask = 16'hE5E0;
defparam \Mux6~16 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X59_Y36_N9
dffeas \register[13][25] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\register~70_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~62_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\register[13][25]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \register[13][25] .is_wysiwyg = "true";
defparam \register[13][25] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X59_Y36_N8
cycloneive_lcell_comb \Mux6~17 (
// Equation(s):
// \Mux6~17_combout  = (Selector41 & (Selector5)) # (!Selector41 & ((Selector5 & (\register[13][25]~q )) # (!Selector5 & ((\register[12][25]~q )))))

	.dataa(Selector41),
	.datab(Selector5),
	.datac(\register[13][25]~q ),
	.datad(\register[12][25]~q ),
	.cin(gnd),
	.combout(\Mux6~17_combout ),
	.cout());
// synopsys translate_off
defparam \Mux6~17 .lut_mask = 16'hD9C8;
defparam \Mux6~17 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y35_N24
cycloneive_lcell_comb \Mux6~18 (
// Equation(s):
// \Mux6~18_combout  = (\Mux6~17_combout  & (((\register[15][25]~q )) # (!Selector41))) # (!\Mux6~17_combout  & (Selector41 & ((\register[14][25]~q ))))

	.dataa(\Mux6~17_combout ),
	.datab(Selector41),
	.datac(\register[15][25]~q ),
	.datad(\register[14][25]~q ),
	.cin(gnd),
	.combout(\Mux6~18_combout ),
	.cout());
// synopsys translate_off
defparam \Mux6~18 .lut_mask = 16'hE6A2;
defparam \Mux6~18 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y35_N24
cycloneive_lcell_comb \Mux7~7 (
// Equation(s):
// \Mux7~7_combout  = (Selector2 & ((Selector3) # ((\register[27][24]~q )))) # (!Selector2 & (!Selector3 & (\register[19][24]~q )))

	.dataa(Selector2),
	.datab(Selector3),
	.datac(\register[19][24]~q ),
	.datad(\register[27][24]~q ),
	.cin(gnd),
	.combout(\Mux7~7_combout ),
	.cout());
// synopsys translate_off
defparam \Mux7~7 .lut_mask = 16'hBA98;
defparam \Mux7~7 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y34_N8
cycloneive_lcell_comb \Mux7~8 (
// Equation(s):
// \Mux7~8_combout  = (\Mux7~7_combout  & (((\register[31][24]~q ) # (!Selector3)))) # (!\Mux7~7_combout  & (\register[23][24]~q  & (Selector3)))

	.dataa(\Mux7~7_combout ),
	.datab(\register[23][24]~q ),
	.datac(Selector3),
	.datad(\register[31][24]~q ),
	.cin(gnd),
	.combout(\Mux7~8_combout ),
	.cout());
// synopsys translate_off
defparam \Mux7~8 .lut_mask = 16'hEA4A;
defparam \Mux7~8 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X62_Y37_N5
dffeas \register[28][24] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\register~71_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~57_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\register[28][24]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \register[28][24] .is_wysiwyg = "true";
defparam \register[28][24] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X65_Y34_N12
cycloneive_lcell_comb \Mux7~4 (
// Equation(s):
// \Mux7~4_combout  = (Selector2 & (Selector3)) # (!Selector2 & ((Selector3 & (\register[20][24]~q )) # (!Selector3 & ((\register[16][24]~q )))))

	.dataa(Selector2),
	.datab(Selector3),
	.datac(\register[20][24]~q ),
	.datad(\register[16][24]~q ),
	.cin(gnd),
	.combout(\Mux7~4_combout ),
	.cout());
// synopsys translate_off
defparam \Mux7~4 .lut_mask = 16'hD9C8;
defparam \Mux7~4 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y37_N4
cycloneive_lcell_comb \Mux7~5 (
// Equation(s):
// \Mux7~5_combout  = (Selector2 & ((\Mux7~4_combout  & ((\register[28][24]~q ))) # (!\Mux7~4_combout  & (\register[24][24]~q )))) # (!Selector2 & (((\Mux7~4_combout ))))

	.dataa(Selector2),
	.datab(\register[24][24]~q ),
	.datac(\register[28][24]~q ),
	.datad(\Mux7~4_combout ),
	.cin(gnd),
	.combout(\Mux7~5_combout ),
	.cout());
// synopsys translate_off
defparam \Mux7~5 .lut_mask = 16'hF588;
defparam \Mux7~5 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X67_Y37_N31
dffeas \register[18][24] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\register~71_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~33_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\register[18][24]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \register[18][24] .is_wysiwyg = "true";
defparam \register[18][24] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X67_Y37_N30
cycloneive_lcell_comb \Mux7~2 (
// Equation(s):
// \Mux7~2_combout  = (Selector3 & ((\register[22][24]~q ) # ((Selector2)))) # (!Selector3 & (((\register[18][24]~q  & !Selector2))))

	.dataa(Selector3),
	.datab(\register[22][24]~q ),
	.datac(\register[18][24]~q ),
	.datad(Selector2),
	.cin(gnd),
	.combout(\Mux7~2_combout ),
	.cout());
// synopsys translate_off
defparam \Mux7~2 .lut_mask = 16'hAAD8;
defparam \Mux7~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X68_Y37_N14
cycloneive_lcell_comb \Mux7~3 (
// Equation(s):
// \Mux7~3_combout  = (Selector2 & ((\Mux7~2_combout  & (\register[30][24]~q )) # (!\Mux7~2_combout  & ((\register[26][24]~q ))))) # (!Selector2 & (\Mux7~2_combout ))

	.dataa(Selector2),
	.datab(\Mux7~2_combout ),
	.datac(\register[30][24]~q ),
	.datad(\register[26][24]~q ),
	.cin(gnd),
	.combout(\Mux7~3_combout ),
	.cout());
// synopsys translate_off
defparam \Mux7~3 .lut_mask = 16'hE6C4;
defparam \Mux7~3 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y34_N30
cycloneive_lcell_comb \Mux7~6 (
// Equation(s):
// \Mux7~6_combout  = (Selector5 & (Selector41)) # (!Selector5 & ((Selector41 & ((\Mux7~3_combout ))) # (!Selector41 & (\Mux7~5_combout ))))

	.dataa(Selector5),
	.datab(Selector41),
	.datac(\Mux7~5_combout ),
	.datad(\Mux7~3_combout ),
	.cin(gnd),
	.combout(\Mux7~6_combout ),
	.cout());
// synopsys translate_off
defparam \Mux7~6 .lut_mask = 16'hDC98;
defparam \Mux7~6 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y34_N8
cycloneive_lcell_comb \Mux7~0 (
// Equation(s):
// \Mux7~0_combout  = (Selector3 & (((Selector2)))) # (!Selector3 & ((Selector2 & (\register[25][24]~q )) # (!Selector2 & ((\register[17][24]~q )))))

	.dataa(\register[25][24]~q ),
	.datab(Selector3),
	.datac(\register[17][24]~q ),
	.datad(Selector2),
	.cin(gnd),
	.combout(\Mux7~0_combout ),
	.cout());
// synopsys translate_off
defparam \Mux7~0 .lut_mask = 16'hEE30;
defparam \Mux7~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y34_N24
cycloneive_lcell_comb \register[21][24]~feeder (
// Equation(s):
// \register[21][24]~feeder_combout  = \register~71_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(\register~71_combout ),
	.cin(gnd),
	.combout(\register[21][24]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \register[21][24]~feeder .lut_mask = 16'hFF00;
defparam \register[21][24]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X59_Y34_N25
dffeas \register[21][24] (
	.clk(!CLK),
	.d(\register[21][24]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~22_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\register[21][24]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \register[21][24] .is_wysiwyg = "true";
defparam \register[21][24] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X59_Y34_N16
cycloneive_lcell_comb \Mux7~1 (
// Equation(s):
// \Mux7~1_combout  = (\Mux7~0_combout  & (((\register[29][24]~q ) # (!Selector3)))) # (!\Mux7~0_combout  & (\register[21][24]~q  & (Selector3)))

	.dataa(\Mux7~0_combout ),
	.datab(\register[21][24]~q ),
	.datac(Selector3),
	.datad(\register[29][24]~q ),
	.cin(gnd),
	.combout(\Mux7~1_combout ),
	.cout());
// synopsys translate_off
defparam \Mux7~1 .lut_mask = 16'hEA4A;
defparam \Mux7~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X69_Y31_N17
dffeas \register[5][24] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\register~71_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~59_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\register[5][24]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \register[5][24] .is_wysiwyg = "true";
defparam \register[5][24] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X69_Y31_N16
cycloneive_lcell_comb \Mux7~10 (
// Equation(s):
// \Mux7~10_combout  = (Selector41 & (((Selector5)))) # (!Selector41 & ((Selector5 & ((\register[5][24]~q ))) # (!Selector5 & (\register[4][24]~q ))))

	.dataa(\register[4][24]~q ),
	.datab(Selector41),
	.datac(\register[5][24]~q ),
	.datad(Selector5),
	.cin(gnd),
	.combout(\Mux7~10_combout ),
	.cout());
// synopsys translate_off
defparam \Mux7~10 .lut_mask = 16'hFC22;
defparam \Mux7~10 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X68_Y31_N16
cycloneive_lcell_comb \Mux7~11 (
// Equation(s):
// \Mux7~11_combout  = (Selector41 & ((\Mux7~10_combout  & (\register[7][24]~q )) # (!\Mux7~10_combout  & ((\register[6][24]~q ))))) # (!Selector41 & (((\Mux7~10_combout ))))

	.dataa(Selector41),
	.datab(\register[7][24]~q ),
	.datac(\register[6][24]~q ),
	.datad(\Mux7~10_combout ),
	.cin(gnd),
	.combout(\Mux7~11_combout ),
	.cout());
// synopsys translate_off
defparam \Mux7~11 .lut_mask = 16'hDDA0;
defparam \Mux7~11 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y30_N24
cycloneive_lcell_comb \Mux7~17 (
// Equation(s):
// \Mux7~17_combout  = (Selector41 & (((Selector5)))) # (!Selector41 & ((Selector5 & ((\register[13][24]~q ))) # (!Selector5 & (\register[12][24]~q ))))

	.dataa(\register[12][24]~q ),
	.datab(Selector41),
	.datac(\register[13][24]~q ),
	.datad(Selector5),
	.cin(gnd),
	.combout(\Mux7~17_combout ),
	.cout());
// synopsys translate_off
defparam \Mux7~17 .lut_mask = 16'hFC22;
defparam \Mux7~17 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y36_N16
cycloneive_lcell_comb \Mux7~18 (
// Equation(s):
// \Mux7~18_combout  = (Selector41 & ((\Mux7~17_combout  & (\register[15][24]~q )) # (!\Mux7~17_combout  & ((\register[14][24]~q ))))) # (!Selector41 & (((\Mux7~17_combout ))))

	.dataa(Selector41),
	.datab(\register[15][24]~q ),
	.datac(\Mux7~17_combout ),
	.datad(\register[14][24]~q ),
	.cin(gnd),
	.combout(\Mux7~18_combout ),
	.cout());
// synopsys translate_off
defparam \Mux7~18 .lut_mask = 16'hDAD0;
defparam \Mux7~18 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X69_Y33_N24
cycloneive_lcell_comb \Mux7~14 (
// Equation(s):
// \Mux7~14_combout  = (Selector5 & ((Selector41 & ((\register[3][24]~q ))) # (!Selector41 & (\register[1][24]~q ))))

	.dataa(\register[1][24]~q ),
	.datab(Selector5),
	.datac(\register[3][24]~q ),
	.datad(Selector41),
	.cin(gnd),
	.combout(\Mux7~14_combout ),
	.cout());
// synopsys translate_off
defparam \Mux7~14 .lut_mask = 16'hC088;
defparam \Mux7~14 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X66_Y34_N18
cycloneive_lcell_comb \Mux7~15 (
// Equation(s):
// \Mux7~15_combout  = (\Mux7~14_combout ) # ((Selector41 & (!Selector5 & \register[2][24]~q )))

	.dataa(Selector41),
	.datab(Selector5),
	.datac(\register[2][24]~q ),
	.datad(\Mux7~14_combout ),
	.cin(gnd),
	.combout(\Mux7~15_combout ),
	.cout());
// synopsys translate_off
defparam \Mux7~15 .lut_mask = 16'hFF20;
defparam \Mux7~15 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X67_Y38_N2
cycloneive_lcell_comb \Mux7~12 (
// Equation(s):
// \Mux7~12_combout  = (Selector5 & (Selector41)) # (!Selector5 & ((Selector41 & ((\register[10][24]~q ))) # (!Selector41 & (\register[8][24]~q ))))

	.dataa(Selector5),
	.datab(Selector41),
	.datac(\register[8][24]~q ),
	.datad(\register[10][24]~q ),
	.cin(gnd),
	.combout(\Mux7~12_combout ),
	.cout());
// synopsys translate_off
defparam \Mux7~12 .lut_mask = 16'hDC98;
defparam \Mux7~12 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X66_Y34_N20
cycloneive_lcell_comb \Mux7~13 (
// Equation(s):
// \Mux7~13_combout  = (Selector5 & ((\Mux7~12_combout  & ((\register[11][24]~q ))) # (!\Mux7~12_combout  & (\register[9][24]~q )))) # (!Selector5 & (((\Mux7~12_combout ))))

	.dataa(\register[9][24]~q ),
	.datab(\register[11][24]~q ),
	.datac(Selector5),
	.datad(\Mux7~12_combout ),
	.cin(gnd),
	.combout(\Mux7~13_combout ),
	.cout());
// synopsys translate_off
defparam \Mux7~13 .lut_mask = 16'hCFA0;
defparam \Mux7~13 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y34_N20
cycloneive_lcell_comb \Mux7~16 (
// Equation(s):
// \Mux7~16_combout  = (Selector2 & (((Selector3) # (\Mux7~13_combout )))) # (!Selector2 & (\Mux7~15_combout  & (!Selector3)))

	.dataa(\Mux7~15_combout ),
	.datab(Selector2),
	.datac(Selector3),
	.datad(\Mux7~13_combout ),
	.cin(gnd),
	.combout(\Mux7~16_combout ),
	.cout());
// synopsys translate_off
defparam \Mux7~16 .lut_mask = 16'hCEC2;
defparam \Mux7~16 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y31_N24
cycloneive_lcell_comb \Mux8~7 (
// Equation(s):
// \Mux8~7_combout  = (Selector3 & ((Selector2) # ((\register[23][23]~q )))) # (!Selector3 & (!Selector2 & ((\register[19][23]~q ))))

	.dataa(Selector3),
	.datab(Selector2),
	.datac(\register[23][23]~q ),
	.datad(\register[19][23]~q ),
	.cin(gnd),
	.combout(\Mux8~7_combout ),
	.cout());
// synopsys translate_off
defparam \Mux8~7 .lut_mask = 16'hB9A8;
defparam \Mux8~7 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X63_Y31_N4
cycloneive_lcell_comb \Mux8~8 (
// Equation(s):
// \Mux8~8_combout  = (\Mux8~7_combout  & ((\register[31][23]~q ) # ((!Selector2)))) # (!\Mux8~7_combout  & (((Selector2 & \register[27][23]~q ))))

	.dataa(\register[31][23]~q ),
	.datab(\Mux8~7_combout ),
	.datac(Selector2),
	.datad(\register[27][23]~q ),
	.cin(gnd),
	.combout(\Mux8~8_combout ),
	.cout());
// synopsys translate_off
defparam \Mux8~8 .lut_mask = 16'hBC8C;
defparam \Mux8~8 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y34_N24
cycloneive_lcell_comb \register[17][23]~feeder (
// Equation(s):
// \register[17][23]~feeder_combout  = \register~72_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(\register~72_combout ),
	.cin(gnd),
	.combout(\register[17][23]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \register[17][23]~feeder .lut_mask = 16'hFF00;
defparam \register[17][23]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X62_Y34_N25
dffeas \register[17][23] (
	.clk(!CLK),
	.d(\register[17][23]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~26_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\register[17][23]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \register[17][23] .is_wysiwyg = "true";
defparam \register[17][23] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X62_Y33_N28
cycloneive_lcell_comb \Mux8~0 (
// Equation(s):
// \Mux8~0_combout  = (Selector2 & (Selector3)) # (!Selector2 & ((Selector3 & (\register[21][23]~q )) # (!Selector3 & ((\register[17][23]~q )))))

	.dataa(Selector2),
	.datab(Selector3),
	.datac(\register[21][23]~q ),
	.datad(\register[17][23]~q ),
	.cin(gnd),
	.combout(\Mux8~0_combout ),
	.cout());
// synopsys translate_off
defparam \Mux8~0 .lut_mask = 16'hD9C8;
defparam \Mux8~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X70_Y37_N28
cycloneive_lcell_comb \Mux8~1 (
// Equation(s):
// \Mux8~1_combout  = (Selector2 & ((\Mux8~0_combout  & (\register[29][23]~q )) # (!\Mux8~0_combout  & ((\register[25][23]~q ))))) # (!Selector2 & (((\Mux8~0_combout ))))

	.dataa(\register[29][23]~q ),
	.datab(\register[25][23]~q ),
	.datac(Selector2),
	.datad(\Mux8~0_combout ),
	.cin(gnd),
	.combout(\Mux8~1_combout ),
	.cout());
// synopsys translate_off
defparam \Mux8~1 .lut_mask = 16'hAFC0;
defparam \Mux8~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X68_Y38_N22
cycloneive_lcell_comb \register[18][23]~feeder (
// Equation(s):
// \register[18][23]~feeder_combout  = \register~72_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(\register~72_combout ),
	.datad(gnd),
	.cin(gnd),
	.combout(\register[18][23]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \register[18][23]~feeder .lut_mask = 16'hF0F0;
defparam \register[18][23]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X68_Y38_N23
dffeas \register[18][23] (
	.clk(!CLK),
	.d(\register[18][23]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~33_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\register[18][23]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \register[18][23] .is_wysiwyg = "true";
defparam \register[18][23] .power_up = "low";
// synopsys translate_on

// Location: FF_X68_Y38_N17
dffeas \register[26][23] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\register~72_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~54_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\register[26][23]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \register[26][23] .is_wysiwyg = "true";
defparam \register[26][23] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X68_Y38_N16
cycloneive_lcell_comb \Mux8~2 (
// Equation(s):
// \Mux8~2_combout  = (Selector3 & (((Selector2)))) # (!Selector3 & ((Selector2 & ((\register[26][23]~q ))) # (!Selector2 & (\register[18][23]~q ))))

	.dataa(Selector3),
	.datab(\register[18][23]~q ),
	.datac(\register[26][23]~q ),
	.datad(Selector2),
	.cin(gnd),
	.combout(\Mux8~2_combout ),
	.cout());
// synopsys translate_off
defparam \Mux8~2 .lut_mask = 16'hFA44;
defparam \Mux8~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X70_Y37_N14
cycloneive_lcell_comb \Mux8~3 (
// Equation(s):
// \Mux8~3_combout  = (Selector3 & ((\Mux8~2_combout  & (\register[30][23]~q )) # (!\Mux8~2_combout  & ((\register[22][23]~q ))))) # (!Selector3 & (((\Mux8~2_combout ))))

	.dataa(Selector3),
	.datab(\register[30][23]~q ),
	.datac(\Mux8~2_combout ),
	.datad(\register[22][23]~q ),
	.cin(gnd),
	.combout(\Mux8~3_combout ),
	.cout());
// synopsys translate_off
defparam \Mux8~3 .lut_mask = 16'hDAD0;
defparam \Mux8~3 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X70_Y38_N6
cycloneive_lcell_comb \register[16][23]~feeder (
// Equation(s):
// \register[16][23]~feeder_combout  = \register~72_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(\register~72_combout ),
	.datad(gnd),
	.cin(gnd),
	.combout(\register[16][23]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \register[16][23]~feeder .lut_mask = 16'hF0F0;
defparam \register[16][23]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X70_Y38_N7
dffeas \register[16][23] (
	.clk(!CLK),
	.d(\register[16][23]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~36_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\register[16][23]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \register[16][23] .is_wysiwyg = "true";
defparam \register[16][23] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X70_Y38_N28
cycloneive_lcell_comb \Mux8~4 (
// Equation(s):
// \Mux8~4_combout  = (Selector2 & ((Selector3) # ((\register[24][23]~q )))) # (!Selector2 & (!Selector3 & ((\register[16][23]~q ))))

	.dataa(Selector2),
	.datab(Selector3),
	.datac(\register[24][23]~q ),
	.datad(\register[16][23]~q ),
	.cin(gnd),
	.combout(\Mux8~4_combout ),
	.cout());
// synopsys translate_off
defparam \Mux8~4 .lut_mask = 16'hB9A8;
defparam \Mux8~4 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X70_Y38_N30
cycloneive_lcell_comb \Mux8~5 (
// Equation(s):
// \Mux8~5_combout  = (Selector3 & ((\Mux8~4_combout  & ((\register[28][23]~q ))) # (!\Mux8~4_combout  & (\register[20][23]~q )))) # (!Selector3 & (((\Mux8~4_combout ))))

	.dataa(Selector3),
	.datab(\register[20][23]~q ),
	.datac(\register[28][23]~q ),
	.datad(\Mux8~4_combout ),
	.cin(gnd),
	.combout(\Mux8~5_combout ),
	.cout());
// synopsys translate_off
defparam \Mux8~5 .lut_mask = 16'hF588;
defparam \Mux8~5 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X70_Y37_N20
cycloneive_lcell_comb \Mux8~6 (
// Equation(s):
// \Mux8~6_combout  = (Selector5 & (((Selector41)))) # (!Selector5 & ((Selector41 & (\Mux8~3_combout )) # (!Selector41 & ((\Mux8~5_combout )))))

	.dataa(Selector5),
	.datab(\Mux8~3_combout ),
	.datac(Selector41),
	.datad(\Mux8~5_combout ),
	.cin(gnd),
	.combout(\Mux8~6_combout ),
	.cout());
// synopsys translate_off
defparam \Mux8~6 .lut_mask = 16'hE5E0;
defparam \Mux8~6 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X63_Y30_N4
cycloneive_lcell_comb \Mux8~17 (
// Equation(s):
// \Mux8~17_combout  = (Selector41 & (((Selector5)))) # (!Selector41 & ((Selector5 & ((\register[13][23]~q ))) # (!Selector5 & (\register[12][23]~q ))))

	.dataa(\register[12][23]~q ),
	.datab(Selector41),
	.datac(\register[13][23]~q ),
	.datad(Selector5),
	.cin(gnd),
	.combout(\Mux8~17_combout ),
	.cout());
// synopsys translate_off
defparam \Mux8~17 .lut_mask = 16'hFC22;
defparam \Mux8~17 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X70_Y33_N20
cycloneive_lcell_comb \Mux8~18 (
// Equation(s):
// \Mux8~18_combout  = (Selector41 & ((\Mux8~17_combout  & ((\register[15][23]~q ))) # (!\Mux8~17_combout  & (\register[14][23]~q )))) # (!Selector41 & (((\Mux8~17_combout ))))

	.dataa(\register[14][23]~q ),
	.datab(Selector41),
	.datac(\register[15][23]~q ),
	.datad(\Mux8~17_combout ),
	.cin(gnd),
	.combout(\Mux8~18_combout ),
	.cout());
// synopsys translate_off
defparam \Mux8~18 .lut_mask = 16'hF388;
defparam \Mux8~18 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X66_Y40_N24
cycloneive_lcell_comb \Mux8~10 (
// Equation(s):
// \Mux8~10_combout  = (Selector41 & (((\register[10][23]~q ) # (Selector5)))) # (!Selector41 & (\register[8][23]~q  & ((!Selector5))))

	.dataa(\register[8][23]~q ),
	.datab(Selector41),
	.datac(\register[10][23]~q ),
	.datad(Selector5),
	.cin(gnd),
	.combout(\Mux8~10_combout ),
	.cout());
// synopsys translate_off
defparam \Mux8~10 .lut_mask = 16'hCCE2;
defparam \Mux8~10 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X66_Y40_N14
cycloneive_lcell_comb \Mux8~11 (
// Equation(s):
// \Mux8~11_combout  = (\Mux8~10_combout  & ((\register[11][23]~q ) # ((!Selector5)))) # (!\Mux8~10_combout  & (((\register[9][23]~q  & Selector5))))

	.dataa(\register[11][23]~q ),
	.datab(\register[9][23]~q ),
	.datac(\Mux8~10_combout ),
	.datad(Selector5),
	.cin(gnd),
	.combout(\Mux8~11_combout ),
	.cout());
// synopsys translate_off
defparam \Mux8~11 .lut_mask = 16'hACF0;
defparam \Mux8~11 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X69_Y33_N17
dffeas \register[3][23] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\register~72_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~48_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\register[3][23]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \register[3][23] .is_wysiwyg = "true";
defparam \register[3][23] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X69_Y33_N16
cycloneive_lcell_comb \Mux8~14 (
// Equation(s):
// \Mux8~14_combout  = (plif_ifidinstr_l_22 & ((Selector4 & ((\register[3][23]~q ))) # (!Selector4 & (\register[1][23]~q )))) # (!plif_ifidinstr_l_22 & (\register[1][23]~q ))

	.dataa(\register[1][23]~q ),
	.datab(plif_ifidinstr_l_22),
	.datac(\register[3][23]~q ),
	.datad(Selector4),
	.cin(gnd),
	.combout(\Mux8~14_combout ),
	.cout());
// synopsys translate_off
defparam \Mux8~14 .lut_mask = 16'hE2AA;
defparam \Mux8~14 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X70_Y37_N12
cycloneive_lcell_comb \Mux8~15 (
// Equation(s):
// \Mux8~15_combout  = (Selector5 & (((\Mux8~14_combout )))) # (!Selector5 & (\register[2][23]~q  & ((Selector41))))

	.dataa(Selector5),
	.datab(\register[2][23]~q ),
	.datac(\Mux8~14_combout ),
	.datad(Selector41),
	.cin(gnd),
	.combout(\Mux8~15_combout ),
	.cout());
// synopsys translate_off
defparam \Mux8~15 .lut_mask = 16'hE4A0;
defparam \Mux8~15 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X69_Y32_N20
cycloneive_lcell_comb \Mux8~12 (
// Equation(s):
// \Mux8~12_combout  = (Selector5 & (((\register[5][23]~q ) # (Selector41)))) # (!Selector5 & (\register[4][23]~q  & ((!Selector41))))

	.dataa(\register[4][23]~q ),
	.datab(Selector5),
	.datac(\register[5][23]~q ),
	.datad(Selector41),
	.cin(gnd),
	.combout(\Mux8~12_combout ),
	.cout());
// synopsys translate_off
defparam \Mux8~12 .lut_mask = 16'hCCE2;
defparam \Mux8~12 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X68_Y31_N30
cycloneive_lcell_comb \Mux8~13 (
// Equation(s):
// \Mux8~13_combout  = (Selector41 & ((\Mux8~12_combout  & (\register[7][23]~q )) # (!\Mux8~12_combout  & ((\register[6][23]~q ))))) # (!Selector41 & (\Mux8~12_combout ))

	.dataa(Selector41),
	.datab(\Mux8~12_combout ),
	.datac(\register[7][23]~q ),
	.datad(\register[6][23]~q ),
	.cin(gnd),
	.combout(\Mux8~13_combout ),
	.cout());
// synopsys translate_off
defparam \Mux8~13 .lut_mask = 16'hE6C4;
defparam \Mux8~13 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X70_Y37_N18
cycloneive_lcell_comb \Mux8~16 (
// Equation(s):
// \Mux8~16_combout  = (Selector2 & (((Selector3)))) # (!Selector2 & ((Selector3 & ((\Mux8~13_combout ))) # (!Selector3 & (\Mux8~15_combout ))))

	.dataa(\Mux8~15_combout ),
	.datab(Selector2),
	.datac(Selector3),
	.datad(\Mux8~13_combout ),
	.cin(gnd),
	.combout(\Mux8~16_combout ),
	.cout());
// synopsys translate_off
defparam \Mux8~16 .lut_mask = 16'hF2C2;
defparam \Mux8~16 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y37_N18
cycloneive_lcell_comb \Mux9~4 (
// Equation(s):
// \Mux9~4_combout  = (Selector2 & (Selector3)) # (!Selector2 & ((Selector3 & (\register[20][22]~q )) # (!Selector3 & ((\register[16][22]~q )))))

	.dataa(Selector2),
	.datab(Selector3),
	.datac(\register[20][22]~q ),
	.datad(\register[16][22]~q ),
	.cin(gnd),
	.combout(\Mux9~4_combout ),
	.cout());
// synopsys translate_off
defparam \Mux9~4 .lut_mask = 16'hD9C8;
defparam \Mux9~4 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y37_N20
cycloneive_lcell_comb \Mux9~5 (
// Equation(s):
// \Mux9~5_combout  = (Selector2 & ((\Mux9~4_combout  & ((\register[28][22]~q ))) # (!\Mux9~4_combout  & (\register[24][22]~q )))) # (!Selector2 & (((\Mux9~4_combout ))))

	.dataa(Selector2),
	.datab(\register[24][22]~q ),
	.datac(\register[28][22]~q ),
	.datad(\Mux9~4_combout ),
	.cin(gnd),
	.combout(\Mux9~5_combout ),
	.cout());
// synopsys translate_off
defparam \Mux9~5 .lut_mask = 16'hF588;
defparam \Mux9~5 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X69_Y35_N24
cycloneive_lcell_comb \Mux9~2 (
// Equation(s):
// \Mux9~2_combout  = (Selector3 & (((\register[22][22]~q ) # (Selector2)))) # (!Selector3 & (\register[18][22]~q  & ((!Selector2))))

	.dataa(\register[18][22]~q ),
	.datab(Selector3),
	.datac(\register[22][22]~q ),
	.datad(Selector2),
	.cin(gnd),
	.combout(\Mux9~2_combout ),
	.cout());
// synopsys translate_off
defparam \Mux9~2 .lut_mask = 16'hCCE2;
defparam \Mux9~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X68_Y37_N21
dffeas \register[26][22] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\register~73_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~54_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\register[26][22]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \register[26][22] .is_wysiwyg = "true";
defparam \register[26][22] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X68_Y37_N20
cycloneive_lcell_comb \Mux9~3 (
// Equation(s):
// \Mux9~3_combout  = (Selector2 & ((\Mux9~2_combout  & ((\register[30][22]~q ))) # (!\Mux9~2_combout  & (\register[26][22]~q )))) # (!Selector2 & (\Mux9~2_combout ))

	.dataa(Selector2),
	.datab(\Mux9~2_combout ),
	.datac(\register[26][22]~q ),
	.datad(\register[30][22]~q ),
	.cin(gnd),
	.combout(\Mux9~3_combout ),
	.cout());
// synopsys translate_off
defparam \Mux9~3 .lut_mask = 16'hEC64;
defparam \Mux9~3 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X68_Y36_N10
cycloneive_lcell_comb \Mux9~6 (
// Equation(s):
// \Mux9~6_combout  = (Selector41 & ((Selector5) # ((\Mux9~3_combout )))) # (!Selector41 & (!Selector5 & (\Mux9~5_combout )))

	.dataa(Selector41),
	.datab(Selector5),
	.datac(\Mux9~5_combout ),
	.datad(\Mux9~3_combout ),
	.cin(gnd),
	.combout(\Mux9~6_combout ),
	.cout());
// synopsys translate_off
defparam \Mux9~6 .lut_mask = 16'hBA98;
defparam \Mux9~6 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y39_N22
cycloneive_lcell_comb \Mux9~7 (
// Equation(s):
// \Mux9~7_combout  = (Selector3 & (((Selector2)))) # (!Selector3 & ((Selector2 & ((\register[27][22]~q ))) # (!Selector2 & (\register[19][22]~q ))))

	.dataa(Selector3),
	.datab(\register[19][22]~q ),
	.datac(\register[27][22]~q ),
	.datad(Selector2),
	.cin(gnd),
	.combout(\Mux9~7_combout ),
	.cout());
// synopsys translate_off
defparam \Mux9~7 .lut_mask = 16'hFA44;
defparam \Mux9~7 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X62_Y38_N7
dffeas \register[23][22] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\register~73_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~37_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\register[23][22]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \register[23][22] .is_wysiwyg = "true";
defparam \register[23][22] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X62_Y38_N6
cycloneive_lcell_comb \Mux9~8 (
// Equation(s):
// \Mux9~8_combout  = (\Mux9~7_combout  & (((\register[31][22]~q )) # (!Selector3))) # (!\Mux9~7_combout  & (Selector3 & (\register[23][22]~q )))

	.dataa(\Mux9~7_combout ),
	.datab(Selector3),
	.datac(\register[23][22]~q ),
	.datad(\register[31][22]~q ),
	.cin(gnd),
	.combout(\Mux9~8_combout ),
	.cout());
// synopsys translate_off
defparam \Mux9~8 .lut_mask = 16'hEA62;
defparam \Mux9~8 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y36_N22
cycloneive_lcell_comb \Mux9~0 (
// Equation(s):
// \Mux9~0_combout  = (Selector2 & ((\register[25][22]~q ) # ((Selector3)))) # (!Selector2 & (((\register[17][22]~q  & !Selector3))))

	.dataa(Selector2),
	.datab(\register[25][22]~q ),
	.datac(\register[17][22]~q ),
	.datad(Selector3),
	.cin(gnd),
	.combout(\Mux9~0_combout ),
	.cout());
// synopsys translate_off
defparam \Mux9~0 .lut_mask = 16'hAAD8;
defparam \Mux9~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X68_Y36_N24
cycloneive_lcell_comb \Mux9~1 (
// Equation(s):
// \Mux9~1_combout  = (Selector3 & ((\Mux9~0_combout  & (\register[29][22]~q )) # (!\Mux9~0_combout  & ((\register[21][22]~q ))))) # (!Selector3 & (((\Mux9~0_combout ))))

	.dataa(\register[29][22]~q ),
	.datab(\register[21][22]~q ),
	.datac(Selector3),
	.datad(\Mux9~0_combout ),
	.cin(gnd),
	.combout(\Mux9~1_combout ),
	.cout());
// synopsys translate_off
defparam \Mux9~1 .lut_mask = 16'hAFC0;
defparam \Mux9~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X69_Y31_N0
cycloneive_lcell_comb \Mux9~10 (
// Equation(s):
// \Mux9~10_combout  = (Selector5 & ((Selector41) # ((\register[5][22]~q )))) # (!Selector5 & (!Selector41 & ((\register[4][22]~q ))))

	.dataa(Selector5),
	.datab(Selector41),
	.datac(\register[5][22]~q ),
	.datad(\register[4][22]~q ),
	.cin(gnd),
	.combout(\Mux9~10_combout ),
	.cout());
// synopsys translate_off
defparam \Mux9~10 .lut_mask = 16'hB9A8;
defparam \Mux9~10 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y32_N16
cycloneive_lcell_comb \register[6][22]~feeder (
// Equation(s):
// \register[6][22]~feeder_combout  = \register~73_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(\register~73_combout ),
	.datad(gnd),
	.cin(gnd),
	.combout(\register[6][22]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \register[6][22]~feeder .lut_mask = 16'hF0F0;
defparam \register[6][22]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X62_Y32_N17
dffeas \register[6][22] (
	.clk(!CLK),
	.d(\register[6][22]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~58_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\register[6][22]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \register[6][22] .is_wysiwyg = "true";
defparam \register[6][22] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X62_Y32_N18
cycloneive_lcell_comb \Mux9~11 (
// Equation(s):
// \Mux9~11_combout  = (Selector41 & ((\Mux9~10_combout  & (\register[7][22]~q )) # (!\Mux9~10_combout  & ((\register[6][22]~q ))))) # (!Selector41 & (((\Mux9~10_combout ))))

	.dataa(\register[7][22]~q ),
	.datab(Selector41),
	.datac(\Mux9~10_combout ),
	.datad(\register[6][22]~q ),
	.cin(gnd),
	.combout(\Mux9~11_combout ),
	.cout());
// synopsys translate_off
defparam \Mux9~11 .lut_mask = 16'hBCB0;
defparam \Mux9~11 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y30_N4
cycloneive_lcell_comb \Mux9~17 (
// Equation(s):
// \Mux9~17_combout  = (Selector41 & (((Selector5)))) # (!Selector41 & ((Selector5 & ((\register[13][22]~q ))) # (!Selector5 & (\register[12][22]~q ))))

	.dataa(\register[12][22]~q ),
	.datab(Selector41),
	.datac(\register[13][22]~q ),
	.datad(Selector5),
	.cin(gnd),
	.combout(\Mux9~17_combout ),
	.cout());
// synopsys translate_off
defparam \Mux9~17 .lut_mask = 16'hFC22;
defparam \Mux9~17 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y32_N30
cycloneive_lcell_comb \Mux9~18 (
// Equation(s):
// \Mux9~18_combout  = (Selector41 & ((\Mux9~17_combout  & (\register[15][22]~q )) # (!\Mux9~17_combout  & ((\register[14][22]~q ))))) # (!Selector41 & (((\Mux9~17_combout ))))

	.dataa(\register[15][22]~q ),
	.datab(Selector41),
	.datac(\register[14][22]~q ),
	.datad(\Mux9~17_combout ),
	.cin(gnd),
	.combout(\Mux9~18_combout ),
	.cout());
// synopsys translate_off
defparam \Mux9~18 .lut_mask = 16'hBBC0;
defparam \Mux9~18 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X68_Y36_N26
cycloneive_lcell_comb \Mux9~15 (
// Equation(s):
// \Mux9~15_combout  = (Selector5 & (\Mux9~14_combout )) # (!Selector5 & (((\register[2][22]~q  & Selector41))))

	.dataa(\Mux9~14_combout ),
	.datab(\register[2][22]~q ),
	.datac(Selector41),
	.datad(Selector5),
	.cin(gnd),
	.combout(\Mux9~15_combout ),
	.cout());
// synopsys translate_off
defparam \Mux9~15 .lut_mask = 16'hAAC0;
defparam \Mux9~15 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X65_Y40_N14
cycloneive_lcell_comb \Mux9~13 (
// Equation(s):
// \Mux9~13_combout  = (\Mux9~12_combout  & (((\register[11][22]~q ) # (!Selector5)))) # (!\Mux9~12_combout  & (\register[9][22]~q  & ((Selector5))))

	.dataa(\Mux9~12_combout ),
	.datab(\register[9][22]~q ),
	.datac(\register[11][22]~q ),
	.datad(Selector5),
	.cin(gnd),
	.combout(\Mux9~13_combout ),
	.cout());
// synopsys translate_off
defparam \Mux9~13 .lut_mask = 16'hE4AA;
defparam \Mux9~13 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X68_Y36_N28
cycloneive_lcell_comb \Mux9~16 (
// Equation(s):
// \Mux9~16_combout  = (Selector2 & ((Selector3) # ((\Mux9~13_combout )))) # (!Selector2 & (!Selector3 & (\Mux9~15_combout )))

	.dataa(Selector2),
	.datab(Selector3),
	.datac(\Mux9~15_combout ),
	.datad(\Mux9~13_combout ),
	.cin(gnd),
	.combout(\Mux9~16_combout ),
	.cout());
// synopsys translate_off
defparam \Mux9~16 .lut_mask = 16'hBA98;
defparam \Mux9~16 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y35_N22
cycloneive_lcell_comb \Mux10~7 (
// Equation(s):
// \Mux10~7_combout  = (Selector2 & (Selector3)) # (!Selector2 & ((Selector3 & (\register[23][21]~q )) # (!Selector3 & ((\register[19][21]~q )))))

	.dataa(Selector2),
	.datab(Selector3),
	.datac(\register[23][21]~q ),
	.datad(\register[19][21]~q ),
	.cin(gnd),
	.combout(\Mux10~7_combout ),
	.cout());
// synopsys translate_off
defparam \Mux10~7 .lut_mask = 16'hD9C8;
defparam \Mux10~7 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y38_N30
cycloneive_lcell_comb \Mux10~8 (
// Equation(s):
// \Mux10~8_combout  = (Selector2 & ((\Mux10~7_combout  & (\register[31][21]~q )) # (!\Mux10~7_combout  & ((\register[27][21]~q ))))) # (!Selector2 & (\Mux10~7_combout ))

	.dataa(Selector2),
	.datab(\Mux10~7_combout ),
	.datac(\register[31][21]~q ),
	.datad(\register[27][21]~q ),
	.cin(gnd),
	.combout(\Mux10~8_combout ),
	.cout());
// synopsys translate_off
defparam \Mux10~8 .lut_mask = 16'hE6C4;
defparam \Mux10~8 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X63_Y34_N8
cycloneive_lcell_comb \Mux10~0 (
// Equation(s):
// \Mux10~0_combout  = (Selector2 & (((Selector3)))) # (!Selector2 & ((Selector3 & ((\register[21][21]~q ))) # (!Selector3 & (\register[17][21]~q ))))

	.dataa(Selector2),
	.datab(\register[17][21]~q ),
	.datac(\register[21][21]~q ),
	.datad(Selector3),
	.cin(gnd),
	.combout(\Mux10~0_combout ),
	.cout());
// synopsys translate_off
defparam \Mux10~0 .lut_mask = 16'hFA44;
defparam \Mux10~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y34_N0
cycloneive_lcell_comb \Mux10~1 (
// Equation(s):
// \Mux10~1_combout  = (\Mux10~0_combout  & (((\register[29][21]~q ) # (!Selector2)))) # (!\Mux10~0_combout  & (\register[25][21]~q  & ((Selector2))))

	.dataa(\register[25][21]~q ),
	.datab(\register[29][21]~q ),
	.datac(\Mux10~0_combout ),
	.datad(Selector2),
	.cin(gnd),
	.combout(\Mux10~1_combout ),
	.cout());
// synopsys translate_off
defparam \Mux10~1 .lut_mask = 16'hCAF0;
defparam \Mux10~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X69_Y34_N2
cycloneive_lcell_comb \register[16][21]~feeder (
// Equation(s):
// \register[16][21]~feeder_combout  = \register~74_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(\register~74_combout ),
	.datad(gnd),
	.cin(gnd),
	.combout(\register[16][21]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \register[16][21]~feeder .lut_mask = 16'hF0F0;
defparam \register[16][21]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X69_Y34_N3
dffeas \register[16][21] (
	.clk(!CLK),
	.d(\register[16][21]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~36_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\register[16][21]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \register[16][21] .is_wysiwyg = "true";
defparam \register[16][21] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X69_Y34_N20
cycloneive_lcell_comb \Mux10~4 (
// Equation(s):
// \Mux10~4_combout  = (Selector3 & (((Selector2)))) # (!Selector3 & ((Selector2 & ((\register[24][21]~q ))) # (!Selector2 & (\register[16][21]~q ))))

	.dataa(Selector3),
	.datab(\register[16][21]~q ),
	.datac(\register[24][21]~q ),
	.datad(Selector2),
	.cin(gnd),
	.combout(\Mux10~4_combout ),
	.cout());
// synopsys translate_off
defparam \Mux10~4 .lut_mask = 16'hFA44;
defparam \Mux10~4 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y38_N22
cycloneive_lcell_comb \Mux10~5 (
// Equation(s):
// \Mux10~5_combout  = (Selector3 & ((\Mux10~4_combout  & (\register[28][21]~q )) # (!\Mux10~4_combout  & ((\register[20][21]~q ))))) # (!Selector3 & (((\Mux10~4_combout ))))

	.dataa(\register[28][21]~q ),
	.datab(\register[20][21]~q ),
	.datac(Selector3),
	.datad(\Mux10~4_combout ),
	.cin(gnd),
	.combout(\Mux10~5_combout ),
	.cout());
// synopsys translate_off
defparam \Mux10~5 .lut_mask = 16'hAFC0;
defparam \Mux10~5 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X69_Y39_N14
cycloneive_lcell_comb \Mux10~2 (
// Equation(s):
// \Mux10~2_combout  = (Selector3 & (((Selector2)))) # (!Selector3 & ((Selector2 & ((\register[26][21]~q ))) # (!Selector2 & (\register[18][21]~q ))))

	.dataa(Selector3),
	.datab(\register[18][21]~q ),
	.datac(\register[26][21]~q ),
	.datad(Selector2),
	.cin(gnd),
	.combout(\Mux10~2_combout ),
	.cout());
// synopsys translate_off
defparam \Mux10~2 .lut_mask = 16'hFA44;
defparam \Mux10~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X67_Y37_N18
cycloneive_lcell_comb \Mux10~3 (
// Equation(s):
// \Mux10~3_combout  = (Selector3 & ((\Mux10~2_combout  & (\register[30][21]~q )) # (!\Mux10~2_combout  & ((\register[22][21]~q ))))) # (!Selector3 & (((\Mux10~2_combout ))))

	.dataa(\register[30][21]~q ),
	.datab(Selector3),
	.datac(\register[22][21]~q ),
	.datad(\Mux10~2_combout ),
	.cin(gnd),
	.combout(\Mux10~3_combout ),
	.cout());
// synopsys translate_off
defparam \Mux10~3 .lut_mask = 16'hBBC0;
defparam \Mux10~3 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y38_N16
cycloneive_lcell_comb \Mux10~6 (
// Equation(s):
// \Mux10~6_combout  = (Selector5 & (((Selector41)))) # (!Selector5 & ((Selector41 & ((\Mux10~3_combout ))) # (!Selector41 & (\Mux10~5_combout ))))

	.dataa(\Mux10~5_combout ),
	.datab(Selector5),
	.datac(Selector41),
	.datad(\Mux10~3_combout ),
	.cin(gnd),
	.combout(\Mux10~6_combout ),
	.cout());
// synopsys translate_off
defparam \Mux10~6 .lut_mask = 16'hF2C2;
defparam \Mux10~6 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y30_N2
cycloneive_lcell_comb \Mux10~17 (
// Equation(s):
// \Mux10~17_combout  = (Selector5 & ((\register[13][21]~q ) # ((Selector41)))) # (!Selector5 & (((\register[12][21]~q  & !Selector41))))

	.dataa(Selector5),
	.datab(\register[13][21]~q ),
	.datac(\register[12][21]~q ),
	.datad(Selector41),
	.cin(gnd),
	.combout(\Mux10~17_combout ),
	.cout());
// synopsys translate_off
defparam \Mux10~17 .lut_mask = 16'hAAD8;
defparam \Mux10~17 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y38_N20
cycloneive_lcell_comb \Mux10~18 (
// Equation(s):
// \Mux10~18_combout  = (Selector41 & ((\Mux10~17_combout  & (\register[15][21]~q )) # (!\Mux10~17_combout  & ((\register[14][21]~q ))))) # (!Selector41 & (((\Mux10~17_combout ))))

	.dataa(\register[15][21]~q ),
	.datab(\register[14][21]~q ),
	.datac(Selector41),
	.datad(\Mux10~17_combout ),
	.cin(gnd),
	.combout(\Mux10~18_combout ),
	.cout());
// synopsys translate_off
defparam \Mux10~18 .lut_mask = 16'hAFC0;
defparam \Mux10~18 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X66_Y40_N17
dffeas \register[10][21] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\register~74_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~45_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\register[10][21]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \register[10][21] .is_wysiwyg = "true";
defparam \register[10][21] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X66_Y40_N16
cycloneive_lcell_comb \Mux10~10 (
// Equation(s):
// \Mux10~10_combout  = (Selector5 & (((Selector41)))) # (!Selector5 & ((Selector41 & ((\register[10][21]~q ))) # (!Selector41 & (\register[8][21]~q ))))

	.dataa(\register[8][21]~q ),
	.datab(Selector5),
	.datac(\register[10][21]~q ),
	.datad(Selector41),
	.cin(gnd),
	.combout(\Mux10~10_combout ),
	.cout());
// synopsys translate_off
defparam \Mux10~10 .lut_mask = 16'hFC22;
defparam \Mux10~10 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X63_Y34_N18
cycloneive_lcell_comb \Mux10~11 (
// Equation(s):
// \Mux10~11_combout  = (\Mux10~10_combout  & (((\register[11][21]~q ) # (!Selector5)))) # (!\Mux10~10_combout  & (\register[9][21]~q  & ((Selector5))))

	.dataa(\register[9][21]~q ),
	.datab(\register[11][21]~q ),
	.datac(\Mux10~10_combout ),
	.datad(Selector5),
	.cin(gnd),
	.combout(\Mux10~11_combout ),
	.cout());
// synopsys translate_off
defparam \Mux10~11 .lut_mask = 16'hCAF0;
defparam \Mux10~11 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X68_Y31_N10
cycloneive_lcell_comb \Mux10~13 (
// Equation(s):
// \Mux10~13_combout  = (\Mux10~12_combout  & (((\register[7][21]~q ) # (!Selector41)))) # (!\Mux10~12_combout  & (\register[6][21]~q  & ((Selector41))))

	.dataa(\Mux10~12_combout ),
	.datab(\register[6][21]~q ),
	.datac(\register[7][21]~q ),
	.datad(Selector41),
	.cin(gnd),
	.combout(\Mux10~13_combout ),
	.cout());
// synopsys translate_off
defparam \Mux10~13 .lut_mask = 16'hE4AA;
defparam \Mux10~13 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X65_Y33_N4
cycloneive_lcell_comb \Mux10~14 (
// Equation(s):
// \Mux10~14_combout  = (Selector4 & ((plif_ifidinstr_l_22 & ((\register[3][21]~q ))) # (!plif_ifidinstr_l_22 & (\register[1][21]~q )))) # (!Selector4 & (\register[1][21]~q ))

	.dataa(Selector4),
	.datab(\register[1][21]~q ),
	.datac(\register[3][21]~q ),
	.datad(plif_ifidinstr_l_22),
	.cin(gnd),
	.combout(\Mux10~14_combout ),
	.cout());
// synopsys translate_off
defparam \Mux10~14 .lut_mask = 16'hE4CC;
defparam \Mux10~14 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X67_Y34_N20
cycloneive_lcell_comb \Mux10~15 (
// Equation(s):
// \Mux10~15_combout  = (Selector5 & (((\Mux10~14_combout )))) # (!Selector5 & (Selector41 & (\register[2][21]~q )))

	.dataa(Selector41),
	.datab(Selector5),
	.datac(\register[2][21]~q ),
	.datad(\Mux10~14_combout ),
	.cin(gnd),
	.combout(\Mux10~15_combout ),
	.cout());
// synopsys translate_off
defparam \Mux10~15 .lut_mask = 16'hEC20;
defparam \Mux10~15 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y38_N2
cycloneive_lcell_comb \Mux10~16 (
// Equation(s):
// \Mux10~16_combout  = (Selector2 & (Selector3)) # (!Selector2 & ((Selector3 & (\Mux10~13_combout )) # (!Selector3 & ((\Mux10~15_combout )))))

	.dataa(Selector2),
	.datab(Selector3),
	.datac(\Mux10~13_combout ),
	.datad(\Mux10~15_combout ),
	.cin(gnd),
	.combout(\Mux10~16_combout ),
	.cout());
// synopsys translate_off
defparam \Mux10~16 .lut_mask = 16'hD9C8;
defparam \Mux10~16 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y39_N10
cycloneive_lcell_comb \Mux11~7 (
// Equation(s):
// \Mux11~7_combout  = (Selector3 & (Selector2)) # (!Selector3 & ((Selector2 & (\register[27][20]~q )) # (!Selector2 & ((\register[19][20]~q )))))

	.dataa(Selector3),
	.datab(Selector2),
	.datac(\register[27][20]~q ),
	.datad(\register[19][20]~q ),
	.cin(gnd),
	.combout(\Mux11~7_combout ),
	.cout());
// synopsys translate_off
defparam \Mux11~7 .lut_mask = 16'hD9C8;
defparam \Mux11~7 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y40_N4
cycloneive_lcell_comb \Mux11~8 (
// Equation(s):
// \Mux11~8_combout  = (Selector3 & ((\Mux11~7_combout  & ((\register[31][20]~q ))) # (!\Mux11~7_combout  & (\register[23][20]~q )))) # (!Selector3 & (((\Mux11~7_combout ))))

	.dataa(Selector3),
	.datab(\register[23][20]~q ),
	.datac(\register[31][20]~q ),
	.datad(\Mux11~7_combout ),
	.cin(gnd),
	.combout(\Mux11~8_combout ),
	.cout());
// synopsys translate_off
defparam \Mux11~8 .lut_mask = 16'hF588;
defparam \Mux11~8 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y34_N4
cycloneive_lcell_comb \Mux11~0 (
// Equation(s):
// \Mux11~0_combout  = (Selector3 & (((Selector2)))) # (!Selector3 & ((Selector2 & ((\register[25][20]~q ))) # (!Selector2 & (\register[17][20]~q ))))

	.dataa(\register[17][20]~q ),
	.datab(Selector3),
	.datac(\register[25][20]~q ),
	.datad(Selector2),
	.cin(gnd),
	.combout(\Mux11~0_combout ),
	.cout());
// synopsys translate_off
defparam \Mux11~0 .lut_mask = 16'hFC22;
defparam \Mux11~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y34_N14
cycloneive_lcell_comb \Mux11~1 (
// Equation(s):
// \Mux11~1_combout  = (\Mux11~0_combout  & (((\register[29][20]~q ) # (!Selector3)))) # (!\Mux11~0_combout  & (\register[21][20]~q  & (Selector3)))

	.dataa(\register[21][20]~q ),
	.datab(\Mux11~0_combout ),
	.datac(Selector3),
	.datad(\register[29][20]~q ),
	.cin(gnd),
	.combout(\Mux11~1_combout ),
	.cout());
// synopsys translate_off
defparam \Mux11~1 .lut_mask = 16'hEC2C;
defparam \Mux11~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X65_Y39_N1
dffeas \register[16][20] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\register~75_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~36_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\register[16][20]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \register[16][20] .is_wysiwyg = "true";
defparam \register[16][20] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X65_Y39_N14
cycloneive_lcell_comb \Mux11~4 (
// Equation(s):
// \Mux11~4_combout  = (Selector2 & (((Selector3)))) # (!Selector2 & ((Selector3 & ((\register[20][20]~q ))) # (!Selector3 & (\register[16][20]~q ))))

	.dataa(Selector2),
	.datab(\register[16][20]~q ),
	.datac(\register[20][20]~q ),
	.datad(Selector3),
	.cin(gnd),
	.combout(\Mux11~4_combout ),
	.cout());
// synopsys translate_off
defparam \Mux11~4 .lut_mask = 16'hFA44;
defparam \Mux11~4 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X66_Y39_N4
cycloneive_lcell_comb \Mux11~5 (
// Equation(s):
// \Mux11~5_combout  = (Selector2 & ((\Mux11~4_combout  & ((\register[28][20]~q ))) # (!\Mux11~4_combout  & (\register[24][20]~q )))) # (!Selector2 & (((\Mux11~4_combout ))))

	.dataa(\register[24][20]~q ),
	.datab(Selector2),
	.datac(\register[28][20]~q ),
	.datad(\Mux11~4_combout ),
	.cin(gnd),
	.combout(\Mux11~5_combout ),
	.cout());
// synopsys translate_off
defparam \Mux11~5 .lut_mask = 16'hF388;
defparam \Mux11~5 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X69_Y39_N1
dffeas \register[18][20] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\register~75_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~33_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\register[18][20]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \register[18][20] .is_wysiwyg = "true";
defparam \register[18][20] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X69_Y39_N0
cycloneive_lcell_comb \Mux11~2 (
// Equation(s):
// \Mux11~2_combout  = (Selector3 & ((Selector2) # ((\register[22][20]~q )))) # (!Selector3 & (!Selector2 & (\register[18][20]~q )))

	.dataa(Selector3),
	.datab(Selector2),
	.datac(\register[18][20]~q ),
	.datad(\register[22][20]~q ),
	.cin(gnd),
	.combout(\Mux11~2_combout ),
	.cout());
// synopsys translate_off
defparam \Mux11~2 .lut_mask = 16'hBA98;
defparam \Mux11~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y40_N12
cycloneive_lcell_comb \Mux11~3 (
// Equation(s):
// \Mux11~3_combout  = (Selector2 & ((\Mux11~2_combout  & ((\register[30][20]~q ))) # (!\Mux11~2_combout  & (\register[26][20]~q )))) # (!Selector2 & (((\Mux11~2_combout ))))

	.dataa(\register[26][20]~q ),
	.datab(Selector2),
	.datac(\Mux11~2_combout ),
	.datad(\register[30][20]~q ),
	.cin(gnd),
	.combout(\Mux11~3_combout ),
	.cout());
// synopsys translate_off
defparam \Mux11~3 .lut_mask = 16'hF838;
defparam \Mux11~3 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y40_N10
cycloneive_lcell_comb \Mux11~6 (
// Equation(s):
// \Mux11~6_combout  = (Selector5 & (Selector41)) # (!Selector5 & ((Selector41 & ((\Mux11~3_combout ))) # (!Selector41 & (\Mux11~5_combout ))))

	.dataa(Selector5),
	.datab(Selector41),
	.datac(\Mux11~5_combout ),
	.datad(\Mux11~3_combout ),
	.cin(gnd),
	.combout(\Mux11~6_combout ),
	.cout());
// synopsys translate_off
defparam \Mux11~6 .lut_mask = 16'hDC98;
defparam \Mux11~6 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X62_Y41_N23
dffeas \register[8][20] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\register~75_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~46_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\register[8][20]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \register[8][20] .is_wysiwyg = "true";
defparam \register[8][20] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X62_Y41_N22
cycloneive_lcell_comb \Mux11~12 (
// Equation(s):
// \Mux11~12_combout  = (Selector41 & ((Selector5) # ((\register[10][20]~q )))) # (!Selector41 & (!Selector5 & (\register[8][20]~q )))

	.dataa(Selector41),
	.datab(Selector5),
	.datac(\register[8][20]~q ),
	.datad(\register[10][20]~q ),
	.cin(gnd),
	.combout(\Mux11~12_combout ),
	.cout());
// synopsys translate_off
defparam \Mux11~12 .lut_mask = 16'hBA98;
defparam \Mux11~12 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X65_Y40_N2
cycloneive_lcell_comb \Mux11~13 (
// Equation(s):
// \Mux11~13_combout  = (Selector5 & ((\Mux11~12_combout  & ((\register[11][20]~q ))) # (!\Mux11~12_combout  & (\register[9][20]~q )))) # (!Selector5 & (((\Mux11~12_combout ))))

	.dataa(\register[9][20]~q ),
	.datab(Selector5),
	.datac(\register[11][20]~q ),
	.datad(\Mux11~12_combout ),
	.cin(gnd),
	.combout(\Mux11~13_combout ),
	.cout());
// synopsys translate_off
defparam \Mux11~13 .lut_mask = 16'hF388;
defparam \Mux11~13 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X65_Y36_N24
cycloneive_lcell_comb \Mux11~14 (
// Equation(s):
// \Mux11~14_combout  = (Selector4 & ((plif_ifidinstr_l_22 & (\register[3][20]~q )) # (!plif_ifidinstr_l_22 & ((\register[1][20]~q ))))) # (!Selector4 & (((\register[1][20]~q ))))

	.dataa(Selector4),
	.datab(plif_ifidinstr_l_22),
	.datac(\register[3][20]~q ),
	.datad(\register[1][20]~q ),
	.cin(gnd),
	.combout(\Mux11~14_combout ),
	.cout());
// synopsys translate_off
defparam \Mux11~14 .lut_mask = 16'hF780;
defparam \Mux11~14 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X66_Y34_N26
cycloneive_lcell_comb \Mux11~15 (
// Equation(s):
// \Mux11~15_combout  = (Selector5 & (((\Mux11~14_combout )))) # (!Selector5 & (Selector41 & (\register[2][20]~q )))

	.dataa(Selector41),
	.datab(Selector5),
	.datac(\register[2][20]~q ),
	.datad(\Mux11~14_combout ),
	.cin(gnd),
	.combout(\Mux11~15_combout ),
	.cout());
// synopsys translate_off
defparam \Mux11~15 .lut_mask = 16'hEC20;
defparam \Mux11~15 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y40_N24
cycloneive_lcell_comb \Mux11~16 (
// Equation(s):
// \Mux11~16_combout  = (Selector3 & (Selector2)) # (!Selector3 & ((Selector2 & (\Mux11~13_combout )) # (!Selector2 & ((\Mux11~15_combout )))))

	.dataa(Selector3),
	.datab(Selector2),
	.datac(\Mux11~13_combout ),
	.datad(\Mux11~15_combout ),
	.cin(gnd),
	.combout(\Mux11~16_combout ),
	.cout());
// synopsys translate_off
defparam \Mux11~16 .lut_mask = 16'hD9C8;
defparam \Mux11~16 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y30_N14
cycloneive_lcell_comb \Mux11~17 (
// Equation(s):
// \Mux11~17_combout  = (Selector5 & ((Selector41) # ((\register[13][20]~q )))) # (!Selector5 & (!Selector41 & (\register[12][20]~q )))

	.dataa(Selector5),
	.datab(Selector41),
	.datac(\register[12][20]~q ),
	.datad(\register[13][20]~q ),
	.cin(gnd),
	.combout(\Mux11~17_combout ),
	.cout());
// synopsys translate_off
defparam \Mux11~17 .lut_mask = 16'hBA98;
defparam \Mux11~17 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y34_N6
cycloneive_lcell_comb \Mux11~18 (
// Equation(s):
// \Mux11~18_combout  = (\Mux11~17_combout  & (((\register[15][20]~q )) # (!Selector41))) # (!\Mux11~17_combout  & (Selector41 & (\register[14][20]~q )))

	.dataa(\Mux11~17_combout ),
	.datab(Selector41),
	.datac(\register[14][20]~q ),
	.datad(\register[15][20]~q ),
	.cin(gnd),
	.combout(\Mux11~18_combout ),
	.cout());
// synopsys translate_off
defparam \Mux11~18 .lut_mask = 16'hEA62;
defparam \Mux11~18 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X67_Y32_N23
dffeas \register[4][20] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\register~75_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~60_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\register[4][20]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \register[4][20] .is_wysiwyg = "true";
defparam \register[4][20] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X67_Y32_N22
cycloneive_lcell_comb \Mux11~10 (
// Equation(s):
// \Mux11~10_combout  = (Selector41 & (((Selector5)))) # (!Selector41 & ((Selector5 & (\register[5][20]~q )) # (!Selector5 & ((\register[4][20]~q )))))

	.dataa(Selector41),
	.datab(\register[5][20]~q ),
	.datac(\register[4][20]~q ),
	.datad(Selector5),
	.cin(gnd),
	.combout(\Mux11~10_combout ),
	.cout());
// synopsys translate_off
defparam \Mux11~10 .lut_mask = 16'hEE50;
defparam \Mux11~10 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X68_Y31_N4
cycloneive_lcell_comb \Mux11~11 (
// Equation(s):
// \Mux11~11_combout  = (Selector41 & ((\Mux11~10_combout  & (\register[7][20]~q )) # (!\Mux11~10_combout  & ((\register[6][20]~q ))))) # (!Selector41 & (((\Mux11~10_combout ))))

	.dataa(Selector41),
	.datab(\register[7][20]~q ),
	.datac(\register[6][20]~q ),
	.datad(\Mux11~10_combout ),
	.cin(gnd),
	.combout(\Mux11~11_combout ),
	.cout());
// synopsys translate_off
defparam \Mux11~11 .lut_mask = 16'hDDA0;
defparam \Mux11~11 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X63_Y34_N24
cycloneive_lcell_comb \Mux12~0 (
// Equation(s):
// \Mux12~0_combout  = (Selector2 & (((Selector3)))) # (!Selector2 & ((Selector3 & ((\register[21][19]~q ))) # (!Selector3 & (\register[17][19]~q ))))

	.dataa(Selector2),
	.datab(\register[17][19]~q ),
	.datac(\register[21][19]~q ),
	.datad(Selector3),
	.cin(gnd),
	.combout(\Mux12~0_combout ),
	.cout());
// synopsys translate_off
defparam \Mux12~0 .lut_mask = 16'hFA44;
defparam \Mux12~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y36_N4
cycloneive_lcell_comb \Mux12~1 (
// Equation(s):
// \Mux12~1_combout  = (\Mux12~0_combout  & (((\register[29][19]~q ) # (!Selector2)))) # (!\Mux12~0_combout  & (\register[25][19]~q  & (Selector2)))

	.dataa(\register[25][19]~q ),
	.datab(\Mux12~0_combout ),
	.datac(Selector2),
	.datad(\register[29][19]~q ),
	.cin(gnd),
	.combout(\Mux12~1_combout ),
	.cout());
// synopsys translate_off
defparam \Mux12~1 .lut_mask = 16'hEC2C;
defparam \Mux12~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y35_N0
cycloneive_lcell_comb \Mux12~7 (
// Equation(s):
// \Mux12~7_combout  = (Selector2 & (Selector3)) # (!Selector2 & ((Selector3 & (\register[23][19]~q )) # (!Selector3 & ((\register[19][19]~q )))))

	.dataa(Selector2),
	.datab(Selector3),
	.datac(\register[23][19]~q ),
	.datad(\register[19][19]~q ),
	.cin(gnd),
	.combout(\Mux12~7_combout ),
	.cout());
// synopsys translate_off
defparam \Mux12~7 .lut_mask = 16'hD9C8;
defparam \Mux12~7 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X67_Y36_N30
cycloneive_lcell_comb \register[27][19]~feeder (
// Equation(s):
// \register[27][19]~feeder_combout  = \register~76_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(\register~76_combout ),
	.cin(gnd),
	.combout(\register[27][19]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \register[27][19]~feeder .lut_mask = 16'hFF00;
defparam \register[27][19]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X67_Y36_N31
dffeas \register[27][19] (
	.clk(!CLK),
	.d(\register[27][19]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~38_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\register[27][19]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \register[27][19] .is_wysiwyg = "true";
defparam \register[27][19] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X67_Y36_N20
cycloneive_lcell_comb \Mux12~8 (
// Equation(s):
// \Mux12~8_combout  = (\Mux12~7_combout  & ((\register[31][19]~q ) # ((!Selector2)))) # (!\Mux12~7_combout  & (((\register[27][19]~q  & Selector2))))

	.dataa(\register[31][19]~q ),
	.datab(\Mux12~7_combout ),
	.datac(\register[27][19]~q ),
	.datad(Selector2),
	.cin(gnd),
	.combout(\Mux12~8_combout ),
	.cout());
// synopsys translate_off
defparam \Mux12~8 .lut_mask = 16'hB8CC;
defparam \Mux12~8 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X69_Y39_N17
dffeas \register[18][19] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\register~76_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~33_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\register[18][19]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \register[18][19] .is_wysiwyg = "true";
defparam \register[18][19] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X69_Y39_N16
cycloneive_lcell_comb \Mux12~2 (
// Equation(s):
// \Mux12~2_combout  = (Selector2 & ((\register[26][19]~q ) # ((Selector3)))) # (!Selector2 & (((\register[18][19]~q  & !Selector3))))

	.dataa(\register[26][19]~q ),
	.datab(Selector2),
	.datac(\register[18][19]~q ),
	.datad(Selector3),
	.cin(gnd),
	.combout(\Mux12~2_combout ),
	.cout());
// synopsys translate_off
defparam \Mux12~2 .lut_mask = 16'hCCB8;
defparam \Mux12~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X68_Y39_N18
cycloneive_lcell_comb \Mux12~3 (
// Equation(s):
// \Mux12~3_combout  = (Selector3 & ((\Mux12~2_combout  & ((\register[30][19]~q ))) # (!\Mux12~2_combout  & (\register[22][19]~q )))) # (!Selector3 & (((\Mux12~2_combout ))))

	.dataa(Selector3),
	.datab(\register[22][19]~q ),
	.datac(\register[30][19]~q ),
	.datad(\Mux12~2_combout ),
	.cin(gnd),
	.combout(\Mux12~3_combout ),
	.cout());
// synopsys translate_off
defparam \Mux12~3 .lut_mask = 16'hF588;
defparam \Mux12~3 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X66_Y39_N20
cycloneive_lcell_comb \Mux12~4 (
// Equation(s):
// \Mux12~4_combout  = (Selector3 & (Selector2)) # (!Selector3 & ((Selector2 & (\register[24][19]~q )) # (!Selector2 & ((\register[16][19]~q )))))

	.dataa(Selector3),
	.datab(Selector2),
	.datac(\register[24][19]~q ),
	.datad(\register[16][19]~q ),
	.cin(gnd),
	.combout(\Mux12~4_combout ),
	.cout());
// synopsys translate_off
defparam \Mux12~4 .lut_mask = 16'hD9C8;
defparam \Mux12~4 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X67_Y39_N10
cycloneive_lcell_comb \Mux12~5 (
// Equation(s):
// \Mux12~5_combout  = (Selector3 & ((\Mux12~4_combout  & (\register[28][19]~q )) # (!\Mux12~4_combout  & ((\register[20][19]~q ))))) # (!Selector3 & (((\Mux12~4_combout ))))

	.dataa(\register[28][19]~q ),
	.datab(Selector3),
	.datac(\register[20][19]~q ),
	.datad(\Mux12~4_combout ),
	.cin(gnd),
	.combout(\Mux12~5_combout ),
	.cout());
// synopsys translate_off
defparam \Mux12~5 .lut_mask = 16'hBBC0;
defparam \Mux12~5 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X67_Y36_N18
cycloneive_lcell_comb \Mux12~6 (
// Equation(s):
// \Mux12~6_combout  = (Selector5 & (((Selector41)))) # (!Selector5 & ((Selector41 & (\Mux12~3_combout )) # (!Selector41 & ((\Mux12~5_combout )))))

	.dataa(\Mux12~3_combout ),
	.datab(Selector5),
	.datac(\Mux12~5_combout ),
	.datad(Selector41),
	.cin(gnd),
	.combout(\Mux12~6_combout ),
	.cout());
// synopsys translate_off
defparam \Mux12~6 .lut_mask = 16'hEE30;
defparam \Mux12~6 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y36_N24
cycloneive_lcell_comb \Mux12~17 (
// Equation(s):
// \Mux12~17_combout  = (Selector41 & (((Selector5)))) # (!Selector41 & ((Selector5 & (\register[13][19]~q )) # (!Selector5 & ((\register[12][19]~q )))))

	.dataa(\register[13][19]~q ),
	.datab(\register[12][19]~q ),
	.datac(Selector41),
	.datad(Selector5),
	.cin(gnd),
	.combout(\Mux12~17_combout ),
	.cout());
// synopsys translate_off
defparam \Mux12~17 .lut_mask = 16'hFA0C;
defparam \Mux12~17 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y36_N6
cycloneive_lcell_comb \Mux12~18 (
// Equation(s):
// \Mux12~18_combout  = (Selector41 & ((\Mux12~17_combout  & (\register[15][19]~q )) # (!\Mux12~17_combout  & ((\register[14][19]~q ))))) # (!Selector41 & (((\Mux12~17_combout ))))

	.dataa(Selector41),
	.datab(\register[15][19]~q ),
	.datac(\register[14][19]~q ),
	.datad(\Mux12~17_combout ),
	.cin(gnd),
	.combout(\Mux12~18_combout ),
	.cout());
// synopsys translate_off
defparam \Mux12~18 .lut_mask = 16'hDDA0;
defparam \Mux12~18 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X68_Y32_N2
cycloneive_lcell_comb \Mux12~13 (
// Equation(s):
// \Mux12~13_combout  = (\Mux12~12_combout  & (((\register[7][19]~q )) # (!Selector41))) # (!\Mux12~12_combout  & (Selector41 & ((\register[6][19]~q ))))

	.dataa(\Mux12~12_combout ),
	.datab(Selector41),
	.datac(\register[7][19]~q ),
	.datad(\register[6][19]~q ),
	.cin(gnd),
	.combout(\Mux12~13_combout ),
	.cout());
// synopsys translate_off
defparam \Mux12~13 .lut_mask = 16'hE6A2;
defparam \Mux12~13 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y36_N30
cycloneive_lcell_comb \register[2][19]~feeder (
// Equation(s):
// \register[2][19]~feeder_combout  = \register~76_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(\register~76_combout ),
	.cin(gnd),
	.combout(\register[2][19]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \register[2][19]~feeder .lut_mask = 16'hFF00;
defparam \register[2][19]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X59_Y36_N31
dffeas \register[2][19] (
	.clk(!CLK),
	.d(\register[2][19]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~50_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\register[2][19]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \register[2][19] .is_wysiwyg = "true";
defparam \register[2][19] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X65_Y36_N16
cycloneive_lcell_comb \Mux12~14 (
// Equation(s):
// \Mux12~14_combout  = (Selector4 & ((plif_ifidinstr_l_22 & (\register[3][19]~q )) # (!plif_ifidinstr_l_22 & ((\register[1][19]~q ))))) # (!Selector4 & (((\register[1][19]~q ))))

	.dataa(Selector4),
	.datab(plif_ifidinstr_l_22),
	.datac(\register[3][19]~q ),
	.datad(\register[1][19]~q ),
	.cin(gnd),
	.combout(\Mux12~14_combout ),
	.cout());
// synopsys translate_off
defparam \Mux12~14 .lut_mask = 16'hF780;
defparam \Mux12~14 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y36_N22
cycloneive_lcell_comb \Mux12~15 (
// Equation(s):
// \Mux12~15_combout  = (Selector5 & (((\Mux12~14_combout )))) # (!Selector5 & (Selector41 & (\register[2][19]~q )))

	.dataa(Selector41),
	.datab(Selector5),
	.datac(\register[2][19]~q ),
	.datad(\Mux12~14_combout ),
	.cin(gnd),
	.combout(\Mux12~15_combout ),
	.cout());
// synopsys translate_off
defparam \Mux12~15 .lut_mask = 16'hEC20;
defparam \Mux12~15 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X67_Y36_N4
cycloneive_lcell_comb \Mux12~16 (
// Equation(s):
// \Mux12~16_combout  = (Selector3 & ((\Mux12~13_combout ) # ((Selector2)))) # (!Selector3 & (((\Mux12~15_combout  & !Selector2))))

	.dataa(\Mux12~13_combout ),
	.datab(\Mux12~15_combout ),
	.datac(Selector3),
	.datad(Selector2),
	.cin(gnd),
	.combout(\Mux12~16_combout ),
	.cout());
// synopsys translate_off
defparam \Mux12~16 .lut_mask = 16'hF0AC;
defparam \Mux12~16 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X66_Y40_N8
cycloneive_lcell_comb \Mux12~10 (
// Equation(s):
// \Mux12~10_combout  = (Selector5 & (((Selector41)))) # (!Selector5 & ((Selector41 & ((\register[10][19]~q ))) # (!Selector41 & (\register[8][19]~q ))))

	.dataa(\register[8][19]~q ),
	.datab(Selector5),
	.datac(\register[10][19]~q ),
	.datad(Selector41),
	.cin(gnd),
	.combout(\Mux12~10_combout ),
	.cout());
// synopsys translate_off
defparam \Mux12~10 .lut_mask = 16'hFC22;
defparam \Mux12~10 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X65_Y40_N16
cycloneive_lcell_comb \Mux12~11 (
// Equation(s):
// \Mux12~11_combout  = (\Mux12~10_combout  & ((\register[11][19]~q ) # ((!Selector5)))) # (!\Mux12~10_combout  & (((\register[9][19]~q  & Selector5))))

	.dataa(\register[11][19]~q ),
	.datab(\Mux12~10_combout ),
	.datac(\register[9][19]~q ),
	.datad(Selector5),
	.cin(gnd),
	.combout(\Mux12~11_combout ),
	.cout());
// synopsys translate_off
defparam \Mux12~11 .lut_mask = 16'hB8CC;
defparam \Mux12~11 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y38_N4
cycloneive_lcell_comb \Mux13~7 (
// Equation(s):
// \Mux13~7_combout  = (Selector3 & (Selector2)) # (!Selector3 & ((Selector2 & ((\register[27][18]~q ))) # (!Selector2 & (\register[19][18]~q ))))

	.dataa(Selector3),
	.datab(Selector2),
	.datac(\register[19][18]~q ),
	.datad(\register[27][18]~q ),
	.cin(gnd),
	.combout(\Mux13~7_combout ),
	.cout());
// synopsys translate_off
defparam \Mux13~7 .lut_mask = 16'hDC98;
defparam \Mux13~7 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X63_Y36_N26
cycloneive_lcell_comb \Mux13~8 (
// Equation(s):
// \Mux13~8_combout  = (Selector3 & ((\Mux13~7_combout  & (\register[31][18]~q )) # (!\Mux13~7_combout  & ((\register[23][18]~q ))))) # (!Selector3 & (((\Mux13~7_combout ))))

	.dataa(\register[31][18]~q ),
	.datab(\register[23][18]~q ),
	.datac(Selector3),
	.datad(\Mux13~7_combout ),
	.cin(gnd),
	.combout(\Mux13~8_combout ),
	.cout());
// synopsys translate_off
defparam \Mux13~8 .lut_mask = 16'hAFC0;
defparam \Mux13~8 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y36_N8
cycloneive_lcell_comb \Mux13~0 (
// Equation(s):
// \Mux13~0_combout  = (Selector3 & (Selector2)) # (!Selector3 & ((Selector2 & ((\register[25][18]~q ))) # (!Selector2 & (\register[17][18]~q ))))

	.dataa(Selector3),
	.datab(Selector2),
	.datac(\register[17][18]~q ),
	.datad(\register[25][18]~q ),
	.cin(gnd),
	.combout(\Mux13~0_combout ),
	.cout());
// synopsys translate_off
defparam \Mux13~0 .lut_mask = 16'hDC98;
defparam \Mux13~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X63_Y36_N8
cycloneive_lcell_comb \Mux13~1 (
// Equation(s):
// \Mux13~1_combout  = (Selector3 & ((\Mux13~0_combout  & ((\register[29][18]~q ))) # (!\Mux13~0_combout  & (\register[21][18]~q )))) # (!Selector3 & (((\Mux13~0_combout ))))

	.dataa(\register[21][18]~q ),
	.datab(\register[29][18]~q ),
	.datac(Selector3),
	.datad(\Mux13~0_combout ),
	.cin(gnd),
	.combout(\Mux13~1_combout ),
	.cout());
// synopsys translate_off
defparam \Mux13~1 .lut_mask = 16'hCFA0;
defparam \Mux13~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X69_Y39_N20
cycloneive_lcell_comb \Mux13~2 (
// Equation(s):
// \Mux13~2_combout  = (Selector3 & ((Selector2) # ((\register[22][18]~q )))) # (!Selector3 & (!Selector2 & (\register[18][18]~q )))

	.dataa(Selector3),
	.datab(Selector2),
	.datac(\register[18][18]~q ),
	.datad(\register[22][18]~q ),
	.cin(gnd),
	.combout(\Mux13~2_combout ),
	.cout());
// synopsys translate_off
defparam \Mux13~2 .lut_mask = 16'hBA98;
defparam \Mux13~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X63_Y36_N22
cycloneive_lcell_comb \Mux13~3 (
// Equation(s):
// \Mux13~3_combout  = (Selector2 & ((\Mux13~2_combout  & (\register[30][18]~q )) # (!\Mux13~2_combout  & ((\register[26][18]~q ))))) # (!Selector2 & (((\Mux13~2_combout ))))

	.dataa(Selector2),
	.datab(\register[30][18]~q ),
	.datac(\Mux13~2_combout ),
	.datad(\register[26][18]~q ),
	.cin(gnd),
	.combout(\Mux13~3_combout ),
	.cout());
// synopsys translate_off
defparam \Mux13~3 .lut_mask = 16'hDAD0;
defparam \Mux13~3 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X66_Y39_N31
dffeas \register[28][18] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\register~77_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~57_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\register[28][18]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \register[28][18] .is_wysiwyg = "true";
defparam \register[28][18] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X66_Y39_N30
cycloneive_lcell_comb \Mux13~5 (
// Equation(s):
// \Mux13~5_combout  = (\Mux13~4_combout  & (((\register[28][18]~q )) # (!Selector2))) # (!\Mux13~4_combout  & (Selector2 & ((\register[24][18]~q ))))

	.dataa(\Mux13~4_combout ),
	.datab(Selector2),
	.datac(\register[28][18]~q ),
	.datad(\register[24][18]~q ),
	.cin(gnd),
	.combout(\Mux13~5_combout ),
	.cout());
// synopsys translate_off
defparam \Mux13~5 .lut_mask = 16'hE6A2;
defparam \Mux13~5 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X63_Y36_N20
cycloneive_lcell_comb \Mux13~6 (
// Equation(s):
// \Mux13~6_combout  = (Selector41 & ((Selector5) # ((\Mux13~3_combout )))) # (!Selector41 & (!Selector5 & ((\Mux13~5_combout ))))

	.dataa(Selector41),
	.datab(Selector5),
	.datac(\Mux13~3_combout ),
	.datad(\Mux13~5_combout ),
	.cin(gnd),
	.combout(\Mux13~6_combout ),
	.cout());
// synopsys translate_off
defparam \Mux13~6 .lut_mask = 16'hB9A8;
defparam \Mux13~6 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X65_Y40_N22
cycloneive_lcell_comb \Mux13~13 (
// Equation(s):
// \Mux13~13_combout  = (\Mux13~12_combout  & (((\register[11][18]~q ) # (!Selector5)))) # (!\Mux13~12_combout  & (\register[9][18]~q  & ((Selector5))))

	.dataa(\Mux13~12_combout ),
	.datab(\register[9][18]~q ),
	.datac(\register[11][18]~q ),
	.datad(Selector5),
	.cin(gnd),
	.combout(\Mux13~13_combout ),
	.cout());
// synopsys translate_off
defparam \Mux13~13 .lut_mask = 16'hE4AA;
defparam \Mux13~13 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X65_Y33_N11
dffeas \register[1][18] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\register~77_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~49_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\register[1][18]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \register[1][18] .is_wysiwyg = "true";
defparam \register[1][18] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X65_Y33_N10
cycloneive_lcell_comb \Mux13~14 (
// Equation(s):
// \Mux13~14_combout  = (Selector4 & ((plif_ifidinstr_l_22 & (\register[3][18]~q )) # (!plif_ifidinstr_l_22 & ((\register[1][18]~q ))))) # (!Selector4 & (((\register[1][18]~q ))))

	.dataa(\register[3][18]~q ),
	.datab(Selector4),
	.datac(\register[1][18]~q ),
	.datad(plif_ifidinstr_l_22),
	.cin(gnd),
	.combout(\Mux13~14_combout ),
	.cout());
// synopsys translate_off
defparam \Mux13~14 .lut_mask = 16'hB8F0;
defparam \Mux13~14 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X63_Y36_N18
cycloneive_lcell_comb \Mux13~15 (
// Equation(s):
// \Mux13~15_combout  = (Selector5 & (((\Mux13~14_combout )))) # (!Selector5 & (Selector41 & ((\register[2][18]~q ))))

	.dataa(Selector41),
	.datab(Selector5),
	.datac(\Mux13~14_combout ),
	.datad(\register[2][18]~q ),
	.cin(gnd),
	.combout(\Mux13~15_combout ),
	.cout());
// synopsys translate_off
defparam \Mux13~15 .lut_mask = 16'hE2C0;
defparam \Mux13~15 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X63_Y36_N28
cycloneive_lcell_comb \Mux13~16 (
// Equation(s):
// \Mux13~16_combout  = (Selector2 & ((Selector3) # ((\Mux13~13_combout )))) # (!Selector2 & (!Selector3 & ((\Mux13~15_combout ))))

	.dataa(Selector2),
	.datab(Selector3),
	.datac(\Mux13~13_combout ),
	.datad(\Mux13~15_combout ),
	.cin(gnd),
	.combout(\Mux13~16_combout ),
	.cout());
// synopsys translate_off
defparam \Mux13~16 .lut_mask = 16'hB9A8;
defparam \Mux13~16 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X67_Y32_N31
dffeas \register[4][18] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\register~77_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~60_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\register[4][18]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \register[4][18] .is_wysiwyg = "true";
defparam \register[4][18] .power_up = "low";
// synopsys translate_on

// Location: FF_X67_Y32_N5
dffeas \register[5][18] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\register~77_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~59_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\register[5][18]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \register[5][18] .is_wysiwyg = "true";
defparam \register[5][18] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X67_Y32_N30
cycloneive_lcell_comb \Mux13~10 (
// Equation(s):
// \Mux13~10_combout  = (Selector41 & (Selector5)) # (!Selector41 & ((Selector5 & ((\register[5][18]~q ))) # (!Selector5 & (\register[4][18]~q ))))

	.dataa(Selector41),
	.datab(Selector5),
	.datac(\register[4][18]~q ),
	.datad(\register[5][18]~q ),
	.cin(gnd),
	.combout(\Mux13~10_combout ),
	.cout());
// synopsys translate_off
defparam \Mux13~10 .lut_mask = 16'hDC98;
defparam \Mux13~10 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X67_Y33_N10
cycloneive_lcell_comb \Mux13~11 (
// Equation(s):
// \Mux13~11_combout  = (Selector41 & ((\Mux13~10_combout  & (\register[7][18]~q )) # (!\Mux13~10_combout  & ((\register[6][18]~q ))))) # (!Selector41 & (((\Mux13~10_combout ))))

	.dataa(Selector41),
	.datab(\register[7][18]~q ),
	.datac(\register[6][18]~q ),
	.datad(\Mux13~10_combout ),
	.cin(gnd),
	.combout(\Mux13~11_combout ),
	.cout());
// synopsys translate_off
defparam \Mux13~11 .lut_mask = 16'hDDA0;
defparam \Mux13~11 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y36_N4
cycloneive_lcell_comb \Mux13~17 (
// Equation(s):
// \Mux13~17_combout  = (Selector5 & ((\register[13][18]~q ) # ((Selector41)))) # (!Selector5 & (((!Selector41 & \register[12][18]~q ))))

	.dataa(\register[13][18]~q ),
	.datab(Selector5),
	.datac(Selector41),
	.datad(\register[12][18]~q ),
	.cin(gnd),
	.combout(\Mux13~17_combout ),
	.cout());
// synopsys translate_off
defparam \Mux13~17 .lut_mask = 16'hCBC8;
defparam \Mux13~17 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X63_Y36_N2
cycloneive_lcell_comb \Mux13~18 (
// Equation(s):
// \Mux13~18_combout  = (Selector41 & ((\Mux13~17_combout  & ((\register[15][18]~q ))) # (!\Mux13~17_combout  & (\register[14][18]~q )))) # (!Selector41 & (((\Mux13~17_combout ))))

	.dataa(Selector41),
	.datab(\register[14][18]~q ),
	.datac(\register[15][18]~q ),
	.datad(\Mux13~17_combout ),
	.cin(gnd),
	.combout(\Mux13~18_combout ),
	.cout());
// synopsys translate_off
defparam \Mux13~18 .lut_mask = 16'hF588;
defparam \Mux13~18 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X60_Y38_N3
dffeas \register[19][17] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\register~78_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~39_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\register[19][17]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \register[19][17] .is_wysiwyg = "true";
defparam \register[19][17] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X60_Y38_N2
cycloneive_lcell_comb \Mux14~7 (
// Equation(s):
// \Mux14~7_combout  = (Selector3 & ((Selector2) # ((\register[23][17]~q )))) # (!Selector3 & (!Selector2 & (\register[19][17]~q )))

	.dataa(Selector3),
	.datab(Selector2),
	.datac(\register[19][17]~q ),
	.datad(\register[23][17]~q ),
	.cin(gnd),
	.combout(\Mux14~7_combout ),
	.cout());
// synopsys translate_off
defparam \Mux14~7 .lut_mask = 16'hBA98;
defparam \Mux14~7 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y40_N14
cycloneive_lcell_comb \Mux14~8 (
// Equation(s):
// \Mux14~8_combout  = (Selector2 & ((\Mux14~7_combout  & (\register[31][17]~q )) # (!\Mux14~7_combout  & ((\register[27][17]~q ))))) # (!Selector2 & (\Mux14~7_combout ))

	.dataa(Selector2),
	.datab(\Mux14~7_combout ),
	.datac(\register[31][17]~q ),
	.datad(\register[27][17]~q ),
	.cin(gnd),
	.combout(\Mux14~8_combout ),
	.cout());
// synopsys translate_off
defparam \Mux14~8 .lut_mask = 16'hE6C4;
defparam \Mux14~8 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X63_Y34_N6
cycloneive_lcell_comb \Mux14~0 (
// Equation(s):
// \Mux14~0_combout  = (Selector2 & (((Selector3)))) # (!Selector2 & ((Selector3 & ((\register[21][17]~q ))) # (!Selector3 & (\register[17][17]~q ))))

	.dataa(Selector2),
	.datab(\register[17][17]~q ),
	.datac(\register[21][17]~q ),
	.datad(Selector3),
	.cin(gnd),
	.combout(\Mux14~0_combout ),
	.cout());
// synopsys translate_off
defparam \Mux14~0 .lut_mask = 16'hFA44;
defparam \Mux14~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y40_N22
cycloneive_lcell_comb \Mux14~1 (
// Equation(s):
// \Mux14~1_combout  = (Selector2 & ((\Mux14~0_combout  & (\register[29][17]~q )) # (!\Mux14~0_combout  & ((\register[25][17]~q ))))) # (!Selector2 & (((\Mux14~0_combout ))))

	.dataa(Selector2),
	.datab(\register[29][17]~q ),
	.datac(\register[25][17]~q ),
	.datad(\Mux14~0_combout ),
	.cin(gnd),
	.combout(\Mux14~1_combout ),
	.cout());
// synopsys translate_off
defparam \Mux14~1 .lut_mask = 16'hDDA0;
defparam \Mux14~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X68_Y39_N9
dffeas \register[22][17] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\register~78_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~55_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\register[22][17]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \register[22][17] .is_wysiwyg = "true";
defparam \register[22][17] .power_up = "low";
// synopsys translate_on

// Location: FF_X69_Y39_N23
dffeas \register[26][17] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\register~78_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~54_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\register[26][17]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \register[26][17] .is_wysiwyg = "true";
defparam \register[26][17] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X69_Y39_N22
cycloneive_lcell_comb \Mux14~2 (
// Equation(s):
// \Mux14~2_combout  = (Selector3 & (Selector2)) # (!Selector3 & ((Selector2 & (\register[26][17]~q )) # (!Selector2 & ((\register[18][17]~q )))))

	.dataa(Selector3),
	.datab(Selector2),
	.datac(\register[26][17]~q ),
	.datad(\register[18][17]~q ),
	.cin(gnd),
	.combout(\Mux14~2_combout ),
	.cout());
// synopsys translate_off
defparam \Mux14~2 .lut_mask = 16'hD9C8;
defparam \Mux14~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X68_Y39_N8
cycloneive_lcell_comb \Mux14~3 (
// Equation(s):
// \Mux14~3_combout  = (Selector3 & ((\Mux14~2_combout  & (\register[30][17]~q )) # (!\Mux14~2_combout  & ((\register[22][17]~q ))))) # (!Selector3 & (((\Mux14~2_combout ))))

	.dataa(Selector3),
	.datab(\register[30][17]~q ),
	.datac(\register[22][17]~q ),
	.datad(\Mux14~2_combout ),
	.cin(gnd),
	.combout(\Mux14~3_combout ),
	.cout());
// synopsys translate_off
defparam \Mux14~3 .lut_mask = 16'hDDA0;
defparam \Mux14~3 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y40_N16
cycloneive_lcell_comb \Mux14~4 (
// Equation(s):
// \Mux14~4_combout  = (Selector2 & (((\register[24][17]~q ) # (Selector3)))) # (!Selector2 & (\register[16][17]~q  & ((!Selector3))))

	.dataa(Selector2),
	.datab(\register[16][17]~q ),
	.datac(\register[24][17]~q ),
	.datad(Selector3),
	.cin(gnd),
	.combout(\Mux14~4_combout ),
	.cout());
// synopsys translate_off
defparam \Mux14~4 .lut_mask = 16'hAAE4;
defparam \Mux14~4 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y40_N24
cycloneive_lcell_comb \Mux14~5 (
// Equation(s):
// \Mux14~5_combout  = (\Mux14~4_combout  & ((\register[28][17]~q ) # ((!Selector3)))) # (!\Mux14~4_combout  & (((\register[20][17]~q  & Selector3))))

	.dataa(\register[28][17]~q ),
	.datab(\Mux14~4_combout ),
	.datac(\register[20][17]~q ),
	.datad(Selector3),
	.cin(gnd),
	.combout(\Mux14~5_combout ),
	.cout());
// synopsys translate_off
defparam \Mux14~5 .lut_mask = 16'hB8CC;
defparam \Mux14~5 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y40_N24
cycloneive_lcell_comb \Mux14~6 (
// Equation(s):
// \Mux14~6_combout  = (Selector5 & (Selector41)) # (!Selector5 & ((Selector41 & (\Mux14~3_combout )) # (!Selector41 & ((\Mux14~5_combout )))))

	.dataa(Selector5),
	.datab(Selector41),
	.datac(\Mux14~3_combout ),
	.datad(\Mux14~5_combout ),
	.cin(gnd),
	.combout(\Mux14~6_combout ),
	.cout());
// synopsys translate_off
defparam \Mux14~6 .lut_mask = 16'hD9C8;
defparam \Mux14~6 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y36_N18
cycloneive_lcell_comb \Mux14~17 (
// Equation(s):
// \Mux14~17_combout  = (Selector41 & (((Selector5)))) # (!Selector41 & ((Selector5 & ((\register[13][17]~q ))) # (!Selector5 & (\register[12][17]~q ))))

	.dataa(Selector41),
	.datab(\register[12][17]~q ),
	.datac(\register[13][17]~q ),
	.datad(Selector5),
	.cin(gnd),
	.combout(\Mux14~17_combout ),
	.cout());
// synopsys translate_off
defparam \Mux14~17 .lut_mask = 16'hFA44;
defparam \Mux14~17 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y40_N22
cycloneive_lcell_comb \Mux14~18 (
// Equation(s):
// \Mux14~18_combout  = (Selector41 & ((\Mux14~17_combout  & ((\register[15][17]~q ))) # (!\Mux14~17_combout  & (\register[14][17]~q )))) # (!Selector41 & (((\Mux14~17_combout ))))

	.dataa(\register[14][17]~q ),
	.datab(\register[15][17]~q ),
	.datac(Selector41),
	.datad(\Mux14~17_combout ),
	.cin(gnd),
	.combout(\Mux14~18_combout ),
	.cout());
// synopsys translate_off
defparam \Mux14~18 .lut_mask = 16'hCFA0;
defparam \Mux14~18 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X66_Y40_N11
dffeas \register[10][17] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\register~78_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~45_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\register[10][17]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \register[10][17] .is_wysiwyg = "true";
defparam \register[10][17] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X66_Y40_N10
cycloneive_lcell_comb \Mux14~10 (
// Equation(s):
// \Mux14~10_combout  = (Selector41 & (((\register[10][17]~q ) # (Selector5)))) # (!Selector41 & (\register[8][17]~q  & ((!Selector5))))

	.dataa(\register[8][17]~q ),
	.datab(Selector41),
	.datac(\register[10][17]~q ),
	.datad(Selector5),
	.cin(gnd),
	.combout(\Mux14~10_combout ),
	.cout());
// synopsys translate_off
defparam \Mux14~10 .lut_mask = 16'hCCE2;
defparam \Mux14~10 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X63_Y40_N0
cycloneive_lcell_comb \Mux14~11 (
// Equation(s):
// \Mux14~11_combout  = (\Mux14~10_combout  & ((\register[11][17]~q ) # ((!Selector5)))) # (!\Mux14~10_combout  & (((\register[9][17]~q  & Selector5))))

	.dataa(\register[11][17]~q ),
	.datab(\Mux14~10_combout ),
	.datac(\register[9][17]~q ),
	.datad(Selector5),
	.cin(gnd),
	.combout(\Mux14~11_combout ),
	.cout());
// synopsys translate_off
defparam \Mux14~11 .lut_mask = 16'hB8CC;
defparam \Mux14~11 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X69_Y33_N12
cycloneive_lcell_comb \Mux14~14 (
// Equation(s):
// \Mux14~14_combout  = (Selector5 & ((Selector41 & (\register[3][17]~q )) # (!Selector41 & ((\register[1][17]~q )))))

	.dataa(Selector41),
	.datab(Selector5),
	.datac(\register[3][17]~q ),
	.datad(\register[1][17]~q ),
	.cin(gnd),
	.combout(\Mux14~14_combout ),
	.cout());
// synopsys translate_off
defparam \Mux14~14 .lut_mask = 16'hC480;
defparam \Mux14~14 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y36_N2
cycloneive_lcell_comb \Mux14~15 (
// Equation(s):
// \Mux14~15_combout  = (\Mux14~14_combout ) # ((Selector41 & (!Selector5 & \register[2][17]~q )))

	.dataa(Selector41),
	.datab(Selector5),
	.datac(\register[2][17]~q ),
	.datad(\Mux14~14_combout ),
	.cin(gnd),
	.combout(\Mux14~15_combout ),
	.cout());
// synopsys translate_off
defparam \Mux14~15 .lut_mask = 16'hFF20;
defparam \Mux14~15 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X67_Y32_N20
cycloneive_lcell_comb \Mux14~12 (
// Equation(s):
// \Mux14~12_combout  = (Selector41 & (((Selector5)))) # (!Selector41 & ((Selector5 & ((\register[5][17]~q ))) # (!Selector5 & (\register[4][17]~q ))))

	.dataa(\register[4][17]~q ),
	.datab(Selector41),
	.datac(\register[5][17]~q ),
	.datad(Selector5),
	.cin(gnd),
	.combout(\Mux14~12_combout ),
	.cout());
// synopsys translate_off
defparam \Mux14~12 .lut_mask = 16'hFC22;
defparam \Mux14~12 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X68_Y32_N14
cycloneive_lcell_comb \Mux14~13 (
// Equation(s):
// \Mux14~13_combout  = (Selector41 & ((\Mux14~12_combout  & (\register[7][17]~q )) # (!\Mux14~12_combout  & ((\register[6][17]~q ))))) # (!Selector41 & (\Mux14~12_combout ))

	.dataa(Selector41),
	.datab(\Mux14~12_combout ),
	.datac(\register[7][17]~q ),
	.datad(\register[6][17]~q ),
	.cin(gnd),
	.combout(\Mux14~13_combout ),
	.cout());
// synopsys translate_off
defparam \Mux14~13 .lut_mask = 16'hE6C4;
defparam \Mux14~13 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y40_N18
cycloneive_lcell_comb \Mux14~16 (
// Equation(s):
// \Mux14~16_combout  = (Selector3 & (((Selector2) # (\Mux14~13_combout )))) # (!Selector3 & (\Mux14~15_combout  & (!Selector2)))

	.dataa(\Mux14~15_combout ),
	.datab(Selector3),
	.datac(Selector2),
	.datad(\Mux14~13_combout ),
	.cin(gnd),
	.combout(\Mux14~16_combout ),
	.cout());
// synopsys translate_off
defparam \Mux14~16 .lut_mask = 16'hCEC2;
defparam \Mux14~16 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y38_N22
cycloneive_lcell_comb \Mux31~7 (
// Equation(s):
// \Mux31~7_combout  = (Selector3 & (Selector2)) # (!Selector3 & ((Selector2 & ((\register[27][0]~q ))) # (!Selector2 & (\register[19][0]~q ))))

	.dataa(Selector3),
	.datab(Selector2),
	.datac(\register[19][0]~q ),
	.datad(\register[27][0]~q ),
	.cin(gnd),
	.combout(\Mux31~7_combout ),
	.cout());
// synopsys translate_off
defparam \Mux31~7 .lut_mask = 16'hDC98;
defparam \Mux31~7 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y40_N14
cycloneive_lcell_comb \Mux31~8 (
// Equation(s):
// \Mux31~8_combout  = (Selector3 & ((\Mux31~7_combout  & ((\register[31][0]~q ))) # (!\Mux31~7_combout  & (\register[23][0]~q )))) # (!Selector3 & (((\Mux31~7_combout ))))

	.dataa(Selector3),
	.datab(\register[23][0]~q ),
	.datac(\register[31][0]~q ),
	.datad(\Mux31~7_combout ),
	.cin(gnd),
	.combout(\Mux31~8_combout ),
	.cout());
// synopsys translate_off
defparam \Mux31~8 .lut_mask = 16'hF588;
defparam \Mux31~8 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y35_N28
cycloneive_lcell_comb \Mux31~0 (
// Equation(s):
// \Mux31~0_combout  = (Selector2 & ((Selector3) # ((\register[25][0]~q )))) # (!Selector2 & (!Selector3 & (\register[17][0]~q )))

	.dataa(Selector2),
	.datab(Selector3),
	.datac(\register[17][0]~q ),
	.datad(\register[25][0]~q ),
	.cin(gnd),
	.combout(\Mux31~0_combout ),
	.cout());
// synopsys translate_off
defparam \Mux31~0 .lut_mask = 16'hBA98;
defparam \Mux31~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y40_N26
cycloneive_lcell_comb \Mux31~1 (
// Equation(s):
// \Mux31~1_combout  = (\Mux31~0_combout  & ((\register[29][0]~q ) # ((!Selector3)))) # (!\Mux31~0_combout  & (((\register[21][0]~q  & Selector3))))

	.dataa(\register[29][0]~q ),
	.datab(\register[21][0]~q ),
	.datac(\Mux31~0_combout ),
	.datad(Selector3),
	.cin(gnd),
	.combout(\Mux31~1_combout ),
	.cout());
// synopsys translate_off
defparam \Mux31~1 .lut_mask = 16'hACF0;
defparam \Mux31~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X66_Y36_N4
cycloneive_lcell_comb \Mux31~4 (
// Equation(s):
// \Mux31~4_combout  = (Selector2 & (((Selector3)))) # (!Selector2 & ((Selector3 & (\register[20][0]~q )) # (!Selector3 & ((\register[16][0]~q )))))

	.dataa(\register[20][0]~q ),
	.datab(\register[16][0]~q ),
	.datac(Selector2),
	.datad(Selector3),
	.cin(gnd),
	.combout(\Mux31~4_combout ),
	.cout());
// synopsys translate_off
defparam \Mux31~4 .lut_mask = 16'hFA0C;
defparam \Mux31~4 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X66_Y36_N10
cycloneive_lcell_comb \Mux31~5 (
// Equation(s):
// \Mux31~5_combout  = (\Mux31~4_combout  & (((\register[28][0]~q ) # (!Selector2)))) # (!\Mux31~4_combout  & (\register[24][0]~q  & (Selector2)))

	.dataa(\register[24][0]~q ),
	.datab(\Mux31~4_combout ),
	.datac(Selector2),
	.datad(\register[28][0]~q ),
	.cin(gnd),
	.combout(\Mux31~5_combout ),
	.cout());
// synopsys translate_off
defparam \Mux31~5 .lut_mask = 16'hEC2C;
defparam \Mux31~5 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X70_Y39_N26
cycloneive_lcell_comb \register[22][0]~feeder (
// Equation(s):
// \register[22][0]~feeder_combout  = \register~93_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(\register~93_combout ),
	.cin(gnd),
	.combout(\register[22][0]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \register[22][0]~feeder .lut_mask = 16'hFF00;
defparam \register[22][0]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X70_Y39_N27
dffeas \register[22][0] (
	.clk(!CLK),
	.d(\register[22][0]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~55_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\register[22][0]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \register[22][0] .is_wysiwyg = "true";
defparam \register[22][0] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X69_Y39_N4
cycloneive_lcell_comb \Mux31~2 (
// Equation(s):
// \Mux31~2_combout  = (Selector3 & ((Selector2) # ((\register[22][0]~q )))) # (!Selector3 & (!Selector2 & (\register[18][0]~q )))

	.dataa(Selector3),
	.datab(Selector2),
	.datac(\register[18][0]~q ),
	.datad(\register[22][0]~q ),
	.cin(gnd),
	.combout(\Mux31~2_combout ),
	.cout());
// synopsys translate_off
defparam \Mux31~2 .lut_mask = 16'hBA98;
defparam \Mux31~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y36_N24
cycloneive_lcell_comb \Mux31~3 (
// Equation(s):
// \Mux31~3_combout  = (Selector2 & ((\Mux31~2_combout  & ((\register[30][0]~q ))) # (!\Mux31~2_combout  & (\register[26][0]~q )))) # (!Selector2 & (((\Mux31~2_combout ))))

	.dataa(Selector2),
	.datab(\register[26][0]~q ),
	.datac(\register[30][0]~q ),
	.datad(\Mux31~2_combout ),
	.cin(gnd),
	.combout(\Mux31~3_combout ),
	.cout());
// synopsys translate_off
defparam \Mux31~3 .lut_mask = 16'hF588;
defparam \Mux31~3 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y40_N20
cycloneive_lcell_comb \Mux31~6 (
// Equation(s):
// \Mux31~6_combout  = (Selector5 & (Selector41)) # (!Selector5 & ((Selector41 & ((\Mux31~3_combout ))) # (!Selector41 & (\Mux31~5_combout ))))

	.dataa(Selector5),
	.datab(Selector41),
	.datac(\Mux31~5_combout ),
	.datad(\Mux31~3_combout ),
	.cin(gnd),
	.combout(\Mux31~6_combout ),
	.cout());
// synopsys translate_off
defparam \Mux31~6 .lut_mask = 16'hDC98;
defparam \Mux31~6 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X63_Y40_N6
cycloneive_lcell_comb \Mux31~13 (
// Equation(s):
// \Mux31~13_combout  = (\Mux31~12_combout  & (((\register[11][0]~q ) # (!Selector5)))) # (!\Mux31~12_combout  & (\register[9][0]~q  & ((Selector5))))

	.dataa(\Mux31~12_combout ),
	.datab(\register[9][0]~q ),
	.datac(\register[11][0]~q ),
	.datad(Selector5),
	.cin(gnd),
	.combout(\Mux31~13_combout ),
	.cout());
// synopsys translate_off
defparam \Mux31~13 .lut_mask = 16'hE4AA;
defparam \Mux31~13 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X65_Y36_N23
dffeas \register[1][0] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\register~93_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~49_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\register[1][0]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \register[1][0] .is_wysiwyg = "true";
defparam \register[1][0] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X65_Y36_N22
cycloneive_lcell_comb \Mux31~14 (
// Equation(s):
// \Mux31~14_combout  = (Selector4 & ((plif_ifidinstr_l_22 & ((\register[3][0]~q ))) # (!plif_ifidinstr_l_22 & (\register[1][0]~q )))) # (!Selector4 & (((\register[1][0]~q ))))

	.dataa(Selector4),
	.datab(plif_ifidinstr_l_22),
	.datac(\register[1][0]~q ),
	.datad(\register[3][0]~q ),
	.cin(gnd),
	.combout(\Mux31~14_combout ),
	.cout());
// synopsys translate_off
defparam \Mux31~14 .lut_mask = 16'hF870;
defparam \Mux31~14 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y40_N2
cycloneive_lcell_comb \Mux31~15 (
// Equation(s):
// \Mux31~15_combout  = (Selector5 & (((\Mux31~14_combout )))) # (!Selector5 & (Selector41 & (\register[2][0]~q )))

	.dataa(Selector5),
	.datab(Selector41),
	.datac(\register[2][0]~q ),
	.datad(\Mux31~14_combout ),
	.cin(gnd),
	.combout(\Mux31~15_combout ),
	.cout());
// synopsys translate_off
defparam \Mux31~15 .lut_mask = 16'hEA40;
defparam \Mux31~15 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y40_N0
cycloneive_lcell_comb \Mux31~16 (
// Equation(s):
// \Mux31~16_combout  = (Selector3 & (((Selector2)))) # (!Selector3 & ((Selector2 & (\Mux31~13_combout )) # (!Selector2 & ((\Mux31~15_combout )))))

	.dataa(Selector3),
	.datab(\Mux31~13_combout ),
	.datac(Selector2),
	.datad(\Mux31~15_combout ),
	.cin(gnd),
	.combout(\Mux31~16_combout ),
	.cout());
// synopsys translate_off
defparam \Mux31~16 .lut_mask = 16'hE5E0;
defparam \Mux31~16 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X67_Y32_N16
cycloneive_lcell_comb \Mux31~10 (
// Equation(s):
// \Mux31~10_combout  = (Selector41 & (((Selector5)))) # (!Selector41 & ((Selector5 & ((\register[5][0]~q ))) # (!Selector5 & (\register[4][0]~q ))))

	.dataa(\register[4][0]~q ),
	.datab(Selector41),
	.datac(\register[5][0]~q ),
	.datad(Selector5),
	.cin(gnd),
	.combout(\Mux31~10_combout ),
	.cout());
// synopsys translate_off
defparam \Mux31~10 .lut_mask = 16'hFC22;
defparam \Mux31~10 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y32_N12
cycloneive_lcell_comb \Mux31~11 (
// Equation(s):
// \Mux31~11_combout  = (Selector41 & ((\Mux31~10_combout  & (\register[7][0]~q )) # (!\Mux31~10_combout  & ((\register[6][0]~q ))))) # (!Selector41 & (((\Mux31~10_combout ))))

	.dataa(\register[7][0]~q ),
	.datab(Selector41),
	.datac(\register[6][0]~q ),
	.datad(\Mux31~10_combout ),
	.cin(gnd),
	.combout(\Mux31~11_combout ),
	.cout());
// synopsys translate_off
defparam \Mux31~11 .lut_mask = 16'hBBC0;
defparam \Mux31~11 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y33_N20
cycloneive_lcell_comb \Mux31~17 (
// Equation(s):
// \Mux31~17_combout  = (Selector41 & (((Selector5)))) # (!Selector41 & ((Selector5 & ((\register[13][0]~q ))) # (!Selector5 & (\register[12][0]~q ))))

	.dataa(\register[12][0]~q ),
	.datab(Selector41),
	.datac(\register[13][0]~q ),
	.datad(Selector5),
	.cin(gnd),
	.combout(\Mux31~17_combout ),
	.cout());
// synopsys translate_off
defparam \Mux31~17 .lut_mask = 16'hFC22;
defparam \Mux31~17 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y32_N6
cycloneive_lcell_comb \Mux31~18 (
// Equation(s):
// \Mux31~18_combout  = (Selector41 & ((\Mux31~17_combout  & (\register[15][0]~q )) # (!\Mux31~17_combout  & ((\register[14][0]~q ))))) # (!Selector41 & (((\Mux31~17_combout ))))

	.dataa(\register[15][0]~q ),
	.datab(Selector41),
	.datac(\register[14][0]~q ),
	.datad(\Mux31~17_combout ),
	.cin(gnd),
	.combout(\Mux31~18_combout ),
	.cout());
// synopsys translate_off
defparam \Mux31~18 .lut_mask = 16'hBBC0;
defparam \Mux31~18 .sum_lutc_input = "datac";
// synopsys translate_on

endmodule

module memory_control (
	plif_exmemdmemWEN_l,
	plif_exmemdmemREN_l,
	dpifimemREN,
	always1,
	always0,
	ccifiwait_0,
	devpor,
	devclrn,
	devoe);
input 	plif_exmemdmemWEN_l;
input 	plif_exmemdmemREN_l;
input 	dpifimemREN;
input 	always1;
output 	always0;
output 	ccifiwait_0;

// Design Ports Information

input 	devpor;
input 	devclrn;
input 	devoe;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
assign unknown = 1'bx;



// Location: LCCOMB_X54_Y32_N22
cycloneive_lcell_comb \always0~0 (
// Equation(s):
// always0 = (plif_exmemdmemREN_l) # (plif_exmemdmemWEN_l)

	.dataa(plif_exmemdmemREN_l),
	.datab(gnd),
	.datac(gnd),
	.datad(plif_exmemdmemWEN_l),
	.cin(gnd),
	.combout(always0),
	.cout());
// synopsys translate_off
defparam \always0~0 .lut_mask = 16'hFFAA;
defparam \always0~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y33_N14
cycloneive_lcell_comb \ccif.iwait[0]~2 (
// Equation(s):
// ccifiwait_0 = ((plif_exmemdmemWEN_l) # ((plif_exmemdmemREN_l) # (dpifimemREN))) # (!always1)

	.dataa(always1),
	.datab(plif_exmemdmemWEN_l),
	.datac(plif_exmemdmemREN_l),
	.datad(dpifimemREN),
	.cin(gnd),
	.combout(ccifiwait_0),
	.cout());
// synopsys translate_off
defparam \ccif.iwait[0]~2 .lut_mask = 16'hFFFD;
defparam \ccif.iwait[0]~2 .sum_lutc_input = "datac";
// synopsys translate_on

endmodule

module ram (
	is_in_use_reg,
	ramaddr,
	ramaddr1,
	ramaddr2,
	ramaddr3,
	ramaddr4,
	ramaddr5,
	ramaddr6,
	ramaddr7,
	ramaddr8,
	ramaddr9,
	ramaddr10,
	ramaddr11,
	ramaddr12,
	ramaddr13,
	ramaddr14,
	ramaddr15,
	\ramif.ramaddr ,
	ramaddr16,
	ramaddr17,
	ramaddr18,
	ramaddr19,
	\ramif.ramWEN ,
	\ramif.ramREN ,
	always1,
	ramiframload_0,
	ramiframload_1,
	ramiframload_2,
	ramiframload_3,
	ramiframload_4,
	ramiframload_5,
	ramiframload_6,
	ramiframload_7,
	ramiframload_8,
	ramiframload_9,
	ramiframload_10,
	ramiframload_11,
	ramiframload_12,
	ramiframload_13,
	ramiframload_14,
	ramiframload_15,
	ramiframload_16,
	ramiframload_17,
	ramiframload_18,
	ramiframload_19,
	ramiframload_20,
	ramiframload_21,
	ramiframload_22,
	ramiframload_23,
	ramiframload_24,
	ramiframload_25,
	ramiframload_26,
	ramiframload_27,
	ramiframload_28,
	ramiframload_29,
	ramiframload_30,
	ramiframload_31,
	ir_loaded_address_reg_0,
	ir_loaded_address_reg_1,
	ir_loaded_address_reg_2,
	ir_loaded_address_reg_3,
	tdo,
	ramstore,
	ramstore1,
	ramstore2,
	ramstore3,
	ramstore4,
	ramstore5,
	ramstore6,
	ramstore7,
	ramstore8,
	ramstore9,
	ramstore10,
	ramstore11,
	ramstore12,
	ramstore13,
	ramstore14,
	ramstore15,
	ramstore16,
	ramstore17,
	ramstore18,
	ramstore19,
	ramstore20,
	ramstore21,
	ramstore22,
	ramstore23,
	ramstore24,
	ramstore25,
	ramstore26,
	ramstore27,
	ramstore28,
	ramstore29,
	ramstore30,
	ramstore31,
	ramaddr20,
	altera_internal_jtag,
	state_4,
	irf_reg_0_1,
	irf_reg_1_1,
	irf_reg_2_1,
	irf_reg_3_1,
	irf_reg_4_1,
	node_ena_1,
	clr_reg,
	virtual_ir_scan_reg,
	state_3,
	state_5,
	state_8,
	syiftbCTRL,
	syifaddr_1,
	syifaddr_0,
	nRST,
	altera_internal_jtag1,
	nRST1,
	CLK,
	devpor,
	devclrn,
	devoe);
output 	is_in_use_reg;
input 	ramaddr;
input 	ramaddr1;
input 	ramaddr2;
input 	ramaddr3;
input 	ramaddr4;
input 	ramaddr5;
input 	ramaddr6;
input 	ramaddr7;
input 	ramaddr8;
input 	ramaddr9;
input 	ramaddr10;
input 	ramaddr11;
input 	ramaddr12;
input 	ramaddr13;
input 	ramaddr14;
input 	ramaddr15;
input 	[31:0] \ramif.ramaddr ;
input 	ramaddr16;
input 	ramaddr17;
input 	ramaddr18;
input 	ramaddr19;
input 	\ramif.ramWEN ;
input 	\ramif.ramREN ;
output 	always1;
output 	ramiframload_0;
output 	ramiframload_1;
output 	ramiframload_2;
output 	ramiframload_3;
output 	ramiframload_4;
output 	ramiframload_5;
output 	ramiframload_6;
output 	ramiframload_7;
output 	ramiframload_8;
output 	ramiframload_9;
output 	ramiframload_10;
output 	ramiframload_11;
output 	ramiframload_12;
output 	ramiframload_13;
output 	ramiframload_14;
output 	ramiframload_15;
output 	ramiframload_16;
output 	ramiframload_17;
output 	ramiframload_18;
output 	ramiframload_19;
output 	ramiframload_20;
output 	ramiframload_21;
output 	ramiframload_22;
output 	ramiframload_23;
output 	ramiframload_24;
output 	ramiframload_25;
output 	ramiframload_26;
output 	ramiframload_27;
output 	ramiframload_28;
output 	ramiframload_29;
output 	ramiframload_30;
output 	ramiframload_31;
output 	ir_loaded_address_reg_0;
output 	ir_loaded_address_reg_1;
output 	ir_loaded_address_reg_2;
output 	ir_loaded_address_reg_3;
output 	tdo;
input 	ramstore;
input 	ramstore1;
input 	ramstore2;
input 	ramstore3;
input 	ramstore4;
input 	ramstore5;
input 	ramstore6;
input 	ramstore7;
input 	ramstore8;
input 	ramstore9;
input 	ramstore10;
input 	ramstore11;
input 	ramstore12;
input 	ramstore13;
input 	ramstore14;
input 	ramstore15;
input 	ramstore16;
input 	ramstore17;
input 	ramstore18;
input 	ramstore19;
input 	ramstore20;
input 	ramstore21;
input 	ramstore22;
input 	ramstore23;
input 	ramstore24;
input 	ramstore25;
input 	ramstore26;
input 	ramstore27;
input 	ramstore28;
input 	ramstore29;
input 	ramstore30;
input 	ramstore31;
input 	ramaddr20;
input 	altera_internal_jtag;
input 	state_4;
input 	irf_reg_0_1;
input 	irf_reg_1_1;
input 	irf_reg_2_1;
input 	irf_reg_3_1;
input 	irf_reg_4_1;
input 	node_ena_1;
input 	clr_reg;
input 	virtual_ir_scan_reg;
input 	state_3;
input 	state_5;
input 	state_8;
input 	syiftbCTRL;
input 	syifaddr_1;
input 	syifaddr_0;
input 	nRST;
input 	altera_internal_jtag1;
input 	nRST1;
input 	CLK;

// Design Ports Information

input 	devpor;
input 	devclrn;
input 	devoe;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
assign unknown = 1'bx;

wire \altsyncram_component|auto_generated|altsyncram1|ram_block3a32~portadataout ;
wire \altsyncram_component|auto_generated|altsyncram1|ram_block3a0~portadataout ;
wire \altsyncram_component|auto_generated|altsyncram1|ram_block3a33~portadataout ;
wire \altsyncram_component|auto_generated|altsyncram1|ram_block3a1~portadataout ;
wire \altsyncram_component|auto_generated|altsyncram1|ram_block3a34~portadataout ;
wire \altsyncram_component|auto_generated|altsyncram1|ram_block3a2~portadataout ;
wire \altsyncram_component|auto_generated|altsyncram1|ram_block3a35~portadataout ;
wire \altsyncram_component|auto_generated|altsyncram1|ram_block3a3~portadataout ;
wire \altsyncram_component|auto_generated|altsyncram1|ram_block3a36~portadataout ;
wire \altsyncram_component|auto_generated|altsyncram1|ram_block3a4~portadataout ;
wire \altsyncram_component|auto_generated|altsyncram1|ram_block3a37~portadataout ;
wire \altsyncram_component|auto_generated|altsyncram1|ram_block3a5~portadataout ;
wire \altsyncram_component|auto_generated|altsyncram1|ram_block3a38~portadataout ;
wire \altsyncram_component|auto_generated|altsyncram1|ram_block3a6~portadataout ;
wire \altsyncram_component|auto_generated|altsyncram1|ram_block3a39~portadataout ;
wire \altsyncram_component|auto_generated|altsyncram1|ram_block3a7~portadataout ;
wire \altsyncram_component|auto_generated|altsyncram1|ram_block3a40~portadataout ;
wire \altsyncram_component|auto_generated|altsyncram1|ram_block3a8~portadataout ;
wire \altsyncram_component|auto_generated|altsyncram1|ram_block3a41~portadataout ;
wire \altsyncram_component|auto_generated|altsyncram1|ram_block3a9~portadataout ;
wire \altsyncram_component|auto_generated|altsyncram1|ram_block3a42~portadataout ;
wire \altsyncram_component|auto_generated|altsyncram1|ram_block3a10~portadataout ;
wire \altsyncram_component|auto_generated|altsyncram1|ram_block3a43~portadataout ;
wire \altsyncram_component|auto_generated|altsyncram1|ram_block3a11~portadataout ;
wire \altsyncram_component|auto_generated|altsyncram1|ram_block3a44~portadataout ;
wire \altsyncram_component|auto_generated|altsyncram1|ram_block3a12~portadataout ;
wire \altsyncram_component|auto_generated|altsyncram1|ram_block3a45~portadataout ;
wire \altsyncram_component|auto_generated|altsyncram1|ram_block3a13~portadataout ;
wire \altsyncram_component|auto_generated|altsyncram1|ram_block3a46~portadataout ;
wire \altsyncram_component|auto_generated|altsyncram1|ram_block3a14~portadataout ;
wire \altsyncram_component|auto_generated|altsyncram1|ram_block3a47~portadataout ;
wire \altsyncram_component|auto_generated|altsyncram1|ram_block3a15~portadataout ;
wire \altsyncram_component|auto_generated|altsyncram1|ram_block3a48~portadataout ;
wire \altsyncram_component|auto_generated|altsyncram1|ram_block3a16~portadataout ;
wire \altsyncram_component|auto_generated|altsyncram1|ram_block3a49~portadataout ;
wire \altsyncram_component|auto_generated|altsyncram1|ram_block3a17~portadataout ;
wire \altsyncram_component|auto_generated|altsyncram1|ram_block3a50~portadataout ;
wire \altsyncram_component|auto_generated|altsyncram1|ram_block3a18~portadataout ;
wire \altsyncram_component|auto_generated|altsyncram1|ram_block3a51~portadataout ;
wire \altsyncram_component|auto_generated|altsyncram1|ram_block3a19~portadataout ;
wire \altsyncram_component|auto_generated|altsyncram1|ram_block3a52~portadataout ;
wire \altsyncram_component|auto_generated|altsyncram1|ram_block3a20~portadataout ;
wire \altsyncram_component|auto_generated|altsyncram1|ram_block3a53~portadataout ;
wire \altsyncram_component|auto_generated|altsyncram1|ram_block3a21~portadataout ;
wire \altsyncram_component|auto_generated|altsyncram1|ram_block3a54~portadataout ;
wire \altsyncram_component|auto_generated|altsyncram1|ram_block3a22~portadataout ;
wire \altsyncram_component|auto_generated|altsyncram1|ram_block3a55~portadataout ;
wire \altsyncram_component|auto_generated|altsyncram1|ram_block3a23~portadataout ;
wire \altsyncram_component|auto_generated|altsyncram1|ram_block3a56~portadataout ;
wire \altsyncram_component|auto_generated|altsyncram1|ram_block3a24~portadataout ;
wire \altsyncram_component|auto_generated|altsyncram1|ram_block3a57~portadataout ;
wire \altsyncram_component|auto_generated|altsyncram1|ram_block3a25~portadataout ;
wire \altsyncram_component|auto_generated|altsyncram1|ram_block3a58~portadataout ;
wire \altsyncram_component|auto_generated|altsyncram1|ram_block3a26~portadataout ;
wire \altsyncram_component|auto_generated|altsyncram1|ram_block3a59~portadataout ;
wire \altsyncram_component|auto_generated|altsyncram1|ram_block3a27~portadataout ;
wire \altsyncram_component|auto_generated|altsyncram1|ram_block3a60~portadataout ;
wire \altsyncram_component|auto_generated|altsyncram1|ram_block3a28~portadataout ;
wire \altsyncram_component|auto_generated|altsyncram1|ram_block3a61~portadataout ;
wire \altsyncram_component|auto_generated|altsyncram1|ram_block3a29~portadataout ;
wire \altsyncram_component|auto_generated|altsyncram1|ram_block3a62~portadataout ;
wire \altsyncram_component|auto_generated|altsyncram1|ram_block3a30~portadataout ;
wire \altsyncram_component|auto_generated|altsyncram1|ram_block3a63~portadataout ;
wire \altsyncram_component|auto_generated|altsyncram1|ram_block3a31~portadataout ;
wire \Equal2~0_combout ;
wire \Equal2~1_combout ;
wire \Equal2~2_combout ;
wire \Equal2~10_combout ;
wire \Equal2~13_combout ;
wire \Equal2~17_combout ;
wire \addr[3]~feeder_combout ;
wire \addr[18]~feeder_combout ;
wire \addr[24]~feeder_combout ;
wire \addr[28]~feeder_combout ;
wire \addr[7]~feeder_combout ;
wire \always0~0_combout ;
wire \always0~1_combout ;
wire \addr[6]~feeder_combout ;
wire \Equal2~5_combout ;
wire \addr[2]~feeder_combout ;
wire \Equal2~3_combout ;
wire \addr[5]~feeder_combout ;
wire \Equal2~4_combout ;
wire \Equal2~6_combout ;
wire \Equal2~8_combout ;
wire \Equal2~7_combout ;
wire \addr[12]~feeder_combout ;
wire \Equal2~9_combout ;
wire \Equal2~11_combout ;
wire \Equal2~18_combout ;
wire \Equal2~19_combout ;
wire \Equal2~20_combout ;
wire \Equal2~21_combout ;
wire \Equal2~15_combout ;
wire \Equal2~14_combout ;
wire \Equal2~12_combout ;
wire \Equal2~16_combout ;
wire \Equal2~22_combout ;
wire [1:0] en;
wire [31:0] addr;
wire [0:0] \altsyncram_component|auto_generated|altsyncram1|address_reg_a ;


altsyncram_1 altsyncram_component(
	.ram_block3a32(\altsyncram_component|auto_generated|altsyncram1|ram_block3a32~portadataout ),
	.ram_block3a0(\altsyncram_component|auto_generated|altsyncram1|ram_block3a0~portadataout ),
	.ram_block3a33(\altsyncram_component|auto_generated|altsyncram1|ram_block3a33~portadataout ),
	.ram_block3a1(\altsyncram_component|auto_generated|altsyncram1|ram_block3a1~portadataout ),
	.ram_block3a34(\altsyncram_component|auto_generated|altsyncram1|ram_block3a34~portadataout ),
	.ram_block3a2(\altsyncram_component|auto_generated|altsyncram1|ram_block3a2~portadataout ),
	.ram_block3a35(\altsyncram_component|auto_generated|altsyncram1|ram_block3a35~portadataout ),
	.ram_block3a3(\altsyncram_component|auto_generated|altsyncram1|ram_block3a3~portadataout ),
	.ram_block3a36(\altsyncram_component|auto_generated|altsyncram1|ram_block3a36~portadataout ),
	.ram_block3a4(\altsyncram_component|auto_generated|altsyncram1|ram_block3a4~portadataout ),
	.ram_block3a37(\altsyncram_component|auto_generated|altsyncram1|ram_block3a37~portadataout ),
	.ram_block3a5(\altsyncram_component|auto_generated|altsyncram1|ram_block3a5~portadataout ),
	.ram_block3a38(\altsyncram_component|auto_generated|altsyncram1|ram_block3a38~portadataout ),
	.ram_block3a6(\altsyncram_component|auto_generated|altsyncram1|ram_block3a6~portadataout ),
	.ram_block3a39(\altsyncram_component|auto_generated|altsyncram1|ram_block3a39~portadataout ),
	.ram_block3a7(\altsyncram_component|auto_generated|altsyncram1|ram_block3a7~portadataout ),
	.ram_block3a40(\altsyncram_component|auto_generated|altsyncram1|ram_block3a40~portadataout ),
	.ram_block3a8(\altsyncram_component|auto_generated|altsyncram1|ram_block3a8~portadataout ),
	.ram_block3a41(\altsyncram_component|auto_generated|altsyncram1|ram_block3a41~portadataout ),
	.ram_block3a9(\altsyncram_component|auto_generated|altsyncram1|ram_block3a9~portadataout ),
	.ram_block3a42(\altsyncram_component|auto_generated|altsyncram1|ram_block3a42~portadataout ),
	.ram_block3a10(\altsyncram_component|auto_generated|altsyncram1|ram_block3a10~portadataout ),
	.ram_block3a43(\altsyncram_component|auto_generated|altsyncram1|ram_block3a43~portadataout ),
	.ram_block3a11(\altsyncram_component|auto_generated|altsyncram1|ram_block3a11~portadataout ),
	.ram_block3a44(\altsyncram_component|auto_generated|altsyncram1|ram_block3a44~portadataout ),
	.ram_block3a12(\altsyncram_component|auto_generated|altsyncram1|ram_block3a12~portadataout ),
	.ram_block3a45(\altsyncram_component|auto_generated|altsyncram1|ram_block3a45~portadataout ),
	.ram_block3a13(\altsyncram_component|auto_generated|altsyncram1|ram_block3a13~portadataout ),
	.ram_block3a46(\altsyncram_component|auto_generated|altsyncram1|ram_block3a46~portadataout ),
	.ram_block3a14(\altsyncram_component|auto_generated|altsyncram1|ram_block3a14~portadataout ),
	.ram_block3a47(\altsyncram_component|auto_generated|altsyncram1|ram_block3a47~portadataout ),
	.ram_block3a15(\altsyncram_component|auto_generated|altsyncram1|ram_block3a15~portadataout ),
	.ram_block3a48(\altsyncram_component|auto_generated|altsyncram1|ram_block3a48~portadataout ),
	.ram_block3a16(\altsyncram_component|auto_generated|altsyncram1|ram_block3a16~portadataout ),
	.ram_block3a49(\altsyncram_component|auto_generated|altsyncram1|ram_block3a49~portadataout ),
	.ram_block3a17(\altsyncram_component|auto_generated|altsyncram1|ram_block3a17~portadataout ),
	.ram_block3a50(\altsyncram_component|auto_generated|altsyncram1|ram_block3a50~portadataout ),
	.ram_block3a18(\altsyncram_component|auto_generated|altsyncram1|ram_block3a18~portadataout ),
	.ram_block3a51(\altsyncram_component|auto_generated|altsyncram1|ram_block3a51~portadataout ),
	.ram_block3a19(\altsyncram_component|auto_generated|altsyncram1|ram_block3a19~portadataout ),
	.ram_block3a52(\altsyncram_component|auto_generated|altsyncram1|ram_block3a52~portadataout ),
	.ram_block3a20(\altsyncram_component|auto_generated|altsyncram1|ram_block3a20~portadataout ),
	.ram_block3a53(\altsyncram_component|auto_generated|altsyncram1|ram_block3a53~portadataout ),
	.ram_block3a21(\altsyncram_component|auto_generated|altsyncram1|ram_block3a21~portadataout ),
	.ram_block3a54(\altsyncram_component|auto_generated|altsyncram1|ram_block3a54~portadataout ),
	.ram_block3a22(\altsyncram_component|auto_generated|altsyncram1|ram_block3a22~portadataout ),
	.ram_block3a55(\altsyncram_component|auto_generated|altsyncram1|ram_block3a55~portadataout ),
	.ram_block3a23(\altsyncram_component|auto_generated|altsyncram1|ram_block3a23~portadataout ),
	.ram_block3a56(\altsyncram_component|auto_generated|altsyncram1|ram_block3a56~portadataout ),
	.ram_block3a24(\altsyncram_component|auto_generated|altsyncram1|ram_block3a24~portadataout ),
	.ram_block3a57(\altsyncram_component|auto_generated|altsyncram1|ram_block3a57~portadataout ),
	.ram_block3a25(\altsyncram_component|auto_generated|altsyncram1|ram_block3a25~portadataout ),
	.ram_block3a58(\altsyncram_component|auto_generated|altsyncram1|ram_block3a58~portadataout ),
	.ram_block3a26(\altsyncram_component|auto_generated|altsyncram1|ram_block3a26~portadataout ),
	.ram_block3a59(\altsyncram_component|auto_generated|altsyncram1|ram_block3a59~portadataout ),
	.ram_block3a27(\altsyncram_component|auto_generated|altsyncram1|ram_block3a27~portadataout ),
	.ram_block3a60(\altsyncram_component|auto_generated|altsyncram1|ram_block3a60~portadataout ),
	.ram_block3a28(\altsyncram_component|auto_generated|altsyncram1|ram_block3a28~portadataout ),
	.ram_block3a61(\altsyncram_component|auto_generated|altsyncram1|ram_block3a61~portadataout ),
	.ram_block3a29(\altsyncram_component|auto_generated|altsyncram1|ram_block3a29~portadataout ),
	.ram_block3a62(\altsyncram_component|auto_generated|altsyncram1|ram_block3a62~portadataout ),
	.ram_block3a30(\altsyncram_component|auto_generated|altsyncram1|ram_block3a30~portadataout ),
	.ram_block3a63(\altsyncram_component|auto_generated|altsyncram1|ram_block3a63~portadataout ),
	.ram_block3a31(\altsyncram_component|auto_generated|altsyncram1|ram_block3a31~portadataout ),
	.is_in_use_reg(is_in_use_reg),
	.address_reg_a_0(\altsyncram_component|auto_generated|altsyncram1|address_reg_a [0]),
	.address_a({ramaddr20,ramaddr15,ramaddr12,ramaddr13,ramaddr10,ramaddr11,ramaddr8,ramaddr9,ramaddr6,ramaddr7,ramaddr4,ramaddr5,ramaddr2,ramaddr3}),
	.ramaddr(ramaddr14),
	.ramWEN(\ramif.ramWEN ),
	.always1(always1),
	.ir_loaded_address_reg_0(ir_loaded_address_reg_0),
	.ir_loaded_address_reg_1(ir_loaded_address_reg_1),
	.ir_loaded_address_reg_2(ir_loaded_address_reg_2),
	.ir_loaded_address_reg_3(ir_loaded_address_reg_3),
	.tdo(tdo),
	.data_a({ramstore31,ramstore30,ramstore29,ramstore28,ramstore27,ramstore26,ramstore25,ramstore24,ramstore23,ramstore22,ramstore21,ramstore20,ramstore19,ramstore18,ramstore17,ramstore16,ramstore15,ramstore14,ramstore13,ramstore12,ramstore11,ramstore10,ramstore9,ramstore8,ramstore7,ramstore6,
ramstore5,ramstore4,ramstore3,ramstore2,ramstore1,ramstore}),
	.altera_internal_jtag(altera_internal_jtag),
	.state_4(state_4),
	.irf_reg_0_1(irf_reg_0_1),
	.irf_reg_1_1(irf_reg_1_1),
	.irf_reg_2_1(irf_reg_2_1),
	.irf_reg_3_1(irf_reg_3_1),
	.irf_reg_4_1(irf_reg_4_1),
	.node_ena_1(node_ena_1),
	.clr_reg(clr_reg),
	.virtual_ir_scan_reg(virtual_ir_scan_reg),
	.state_3(state_3),
	.state_5(state_5),
	.state_8(state_8),
	.altera_internal_jtag1(altera_internal_jtag1),
	.clock0(CLK),
	.devpor(devpor),
	.devclrn(devclrn),
	.devoe(devoe));

// Location: FF_X49_Y34_N3
dffeas \addr[1] (
	.clk(CLK),
	.d(\ramif.ramaddr [1]),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~1_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(addr[1]),
	.prn(vcc));
// synopsys translate_off
defparam \addr[1] .is_wysiwyg = "true";
defparam \addr[1] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X49_Y34_N12
cycloneive_lcell_comb \Equal2~0 (
// Equation(s):
// \Equal2~0_combout  = addr[1] $ (((\syif.addr[1]~input_o  & \syif.tbCTRL~input_o )))

	.dataa(syifaddr_1),
	.datab(syiftbCTRL),
	.datac(gnd),
	.datad(addr[1]),
	.cin(gnd),
	.combout(\Equal2~0_combout ),
	.cout());
// synopsys translate_off
defparam \Equal2~0 .lut_mask = 16'h7788;
defparam \Equal2~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X49_Y34_N15
dffeas \addr[0] (
	.clk(CLK),
	.d(\ramif.ramaddr [0]),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~1_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(addr[0]),
	.prn(vcc));
// synopsys translate_off
defparam \addr[0] .is_wysiwyg = "true";
defparam \addr[0] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X49_Y34_N22
cycloneive_lcell_comb \Equal2~1 (
// Equation(s):
// \Equal2~1_combout  = addr[0] $ (((\syif.tbCTRL~input_o  & (\syif.addr[0]~input_o )) # (!\syif.tbCTRL~input_o  & ((\ramaddr~1_combout )))))

	.dataa(syiftbCTRL),
	.datab(syifaddr_0),
	.datac(addr[0]),
	.datad(ramaddr1),
	.cin(gnd),
	.combout(\Equal2~1_combout ),
	.cout());
// synopsys translate_off
defparam \Equal2~1 .lut_mask = 16'h2D78;
defparam \Equal2~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X49_Y34_N4
cycloneive_lcell_comb \Equal2~2 (
// Equation(s):
// \Equal2~2_combout  = (!\Equal2~1_combout  & (\Equal2~0_combout  $ (((\syif.tbCTRL~input_o ) # (!\ramaddr~0_combout )))))

	.dataa(\Equal2~0_combout ),
	.datab(syiftbCTRL),
	.datac(\Equal2~1_combout ),
	.datad(ramaddr),
	.cin(gnd),
	.combout(\Equal2~2_combout ),
	.cout());
// synopsys translate_off
defparam \Equal2~2 .lut_mask = 16'h0605;
defparam \Equal2~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X54_Y35_N23
dffeas \addr[3] (
	.clk(CLK),
	.d(\addr[3]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~1_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(addr[3]),
	.prn(vcc));
// synopsys translate_off
defparam \addr[3] .is_wysiwyg = "true";
defparam \addr[3] .power_up = "low";
// synopsys translate_on

// Location: FF_X49_Y34_N27
dffeas \addr[4] (
	.clk(CLK),
	.d(gnd),
	.asdata(ramaddr5),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\always0~1_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(addr[4]),
	.prn(vcc));
// synopsys translate_off
defparam \addr[4] .is_wysiwyg = "true";
defparam \addr[4] .power_up = "low";
// synopsys translate_on

// Location: FF_X54_Y33_N9
dffeas \addr[8] (
	.clk(CLK),
	.d(ramaddr9),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~1_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(addr[8]),
	.prn(vcc));
// synopsys translate_off
defparam \addr[8] .is_wysiwyg = "true";
defparam \addr[8] .power_up = "low";
// synopsys translate_on

// Location: FF_X54_Y37_N23
dffeas \addr[11] (
	.clk(CLK),
	.d(ramaddr10),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~1_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(addr[11]),
	.prn(vcc));
// synopsys translate_off
defparam \addr[11] .is_wysiwyg = "true";
defparam \addr[11] .power_up = "low";
// synopsys translate_on

// Location: FF_X54_Y32_N23
dffeas \addr[13] (
	.clk(CLK),
	.d(gnd),
	.asdata(ramaddr12),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\always0~1_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(addr[13]),
	.prn(vcc));
// synopsys translate_off
defparam \addr[13] .is_wysiwyg = "true";
defparam \addr[13] .power_up = "low";
// synopsys translate_on

// Location: FF_X52_Y34_N29
dffeas \addr[14] (
	.clk(CLK),
	.d(gnd),
	.asdata(ramaddr15),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\always0~1_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(addr[14]),
	.prn(vcc));
// synopsys translate_off
defparam \addr[14] .is_wysiwyg = "true";
defparam \addr[14] .power_up = "low";
// synopsys translate_on

// Location: FF_X52_Y34_N19
dffeas \addr[15] (
	.clk(CLK),
	.d(gnd),
	.asdata(ramaddr20),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\always0~1_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(addr[15]),
	.prn(vcc));
// synopsys translate_off
defparam \addr[15] .is_wysiwyg = "true";
defparam \addr[15] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X52_Y34_N18
cycloneive_lcell_comb \Equal2~10 (
// Equation(s):
// \Equal2~10_combout  = (\ramaddr~27_combout  & (!addr[15] & (addr[14] $ (!\ramaddr~29_combout )))) # (!\ramaddr~27_combout  & (addr[15] & (addr[14] $ (!\ramaddr~29_combout ))))

	.dataa(ramaddr14),
	.datab(addr[14]),
	.datac(addr[15]),
	.datad(ramaddr15),
	.cin(gnd),
	.combout(\Equal2~10_combout ),
	.cout());
// synopsys translate_off
defparam \Equal2~10 .lut_mask = 16'h4812;
defparam \Equal2~10 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X50_Y34_N9
dffeas \addr[16] (
	.clk(CLK),
	.d(\ramif.ramaddr [16]),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~1_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(addr[16]),
	.prn(vcc));
// synopsys translate_off
defparam \addr[16] .is_wysiwyg = "true";
defparam \addr[16] .power_up = "low";
// synopsys translate_on

// Location: FF_X54_Y33_N13
dffeas \addr[18] (
	.clk(CLK),
	.d(\addr[18]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~1_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(addr[18]),
	.prn(vcc));
// synopsys translate_off
defparam \addr[18] .is_wysiwyg = "true";
defparam \addr[18] .power_up = "low";
// synopsys translate_on

// Location: FF_X54_Y33_N3
dffeas \addr[19] (
	.clk(CLK),
	.d(\ramif.ramaddr [19]),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~1_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(addr[19]),
	.prn(vcc));
// synopsys translate_off
defparam \addr[19] .is_wysiwyg = "true";
defparam \addr[19] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X54_Y33_N22
cycloneive_lcell_comb \Equal2~13 (
// Equation(s):
// \Equal2~13_combout  = (addr[18] & (\ramaddr~37_combout  & (\ramaddr~35_combout  $ (!addr[19])))) # (!addr[18] & (!\ramaddr~37_combout  & (\ramaddr~35_combout  $ (!addr[19]))))

	.dataa(addr[18]),
	.datab(\ramif.ramaddr [19]),
	.datac(addr[19]),
	.datad(ramaddr16),
	.cin(gnd),
	.combout(\Equal2~13_combout ),
	.cout());
// synopsys translate_off
defparam \Equal2~13 .lut_mask = 16'h8241;
defparam \Equal2~13 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X53_Y34_N9
dffeas \addr[22] (
	.clk(CLK),
	.d(\ramif.ramaddr [22]),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~1_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(addr[22]),
	.prn(vcc));
// synopsys translate_off
defparam \addr[22] .is_wysiwyg = "true";
defparam \addr[22] .power_up = "low";
// synopsys translate_on

// Location: FF_X54_Y35_N27
dffeas \addr[24] (
	.clk(CLK),
	.d(\addr[24]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~1_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(addr[24]),
	.prn(vcc));
// synopsys translate_off
defparam \addr[24] .is_wysiwyg = "true";
defparam \addr[24] .power_up = "low";
// synopsys translate_on

// Location: FF_X54_Y35_N13
dffeas \addr[25] (
	.clk(CLK),
	.d(gnd),
	.asdata(ramaddr17),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\always0~1_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(addr[25]),
	.prn(vcc));
// synopsys translate_off
defparam \addr[25] .is_wysiwyg = "true";
defparam \addr[25] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X54_Y35_N30
cycloneive_lcell_comb \Equal2~17 (
// Equation(s):
// \Equal2~17_combout  = (addr[25] & (\ramaddr~47_combout  & (\ramaddr~49_combout  $ (!addr[24])))) # (!addr[25] & (!\ramaddr~47_combout  & (\ramaddr~49_combout  $ (!addr[24]))))

	.dataa(addr[25]),
	.datab(ramaddr18),
	.datac(ramaddr17),
	.datad(addr[24]),
	.cin(gnd),
	.combout(\Equal2~17_combout ),
	.cout());
// synopsys translate_off
defparam \Equal2~17 .lut_mask = 16'h8421;
defparam \Equal2~17 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X54_Y34_N7
dffeas \addr[27] (
	.clk(CLK),
	.d(\ramif.ramaddr [27]),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~1_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(addr[27]),
	.prn(vcc));
// synopsys translate_off
defparam \addr[27] .is_wysiwyg = "true";
defparam \addr[27] .power_up = "low";
// synopsys translate_on

// Location: FF_X50_Y34_N23
dffeas \addr[28] (
	.clk(CLK),
	.d(\addr[28]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~1_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(addr[28]),
	.prn(vcc));
// synopsys translate_off
defparam \addr[28] .is_wysiwyg = "true";
defparam \addr[28] .power_up = "low";
// synopsys translate_on

// Location: FF_X53_Y34_N25
dffeas \addr[30] (
	.clk(CLK),
	.d(\ramif.ramaddr [30]),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~1_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(addr[30]),
	.prn(vcc));
// synopsys translate_off
defparam \addr[30] .is_wysiwyg = "true";
defparam \addr[30] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X54_Y35_N22
cycloneive_lcell_comb \addr[3]~feeder (
// Equation(s):
// \addr[3]~feeder_combout  = \ramaddr~3_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(ramaddr2),
	.datad(gnd),
	.cin(gnd),
	.combout(\addr[3]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \addr[3]~feeder .lut_mask = 16'hF0F0;
defparam \addr[3]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y33_N12
cycloneive_lcell_comb \addr[18]~feeder (
// Equation(s):
// \addr[18]~feeder_combout  = \ramaddr~37_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(ramaddr16),
	.cin(gnd),
	.combout(\addr[18]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \addr[18]~feeder .lut_mask = 16'hFF00;
defparam \addr[18]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y35_N26
cycloneive_lcell_comb \addr[24]~feeder (
// Equation(s):
// \addr[24]~feeder_combout  = \ramaddr~49_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(ramaddr18),
	.datad(gnd),
	.cin(gnd),
	.combout(\addr[24]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \addr[24]~feeder .lut_mask = 16'hF0F0;
defparam \addr[24]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X50_Y34_N22
cycloneive_lcell_comb \addr[28]~feeder (
// Equation(s):
// \addr[28]~feeder_combout  = \ramaddr~57_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(ramaddr19),
	.datad(gnd),
	.cin(gnd),
	.combout(\addr[28]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \addr[28]~feeder .lut_mask = 16'hF0F0;
defparam \addr[28]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y34_N2
cycloneive_lcell_comb \always1~0 (
// Equation(s):
// always1 = ((\Equal2~22_combout  & ((!\ramREN~1_combout ) # (!\ramWEN~0_combout )))) # (!\nRST~input_o )

	.dataa(\ramif.ramWEN ),
	.datab(\ramif.ramREN ),
	.datac(nRST),
	.datad(\Equal2~22_combout ),
	.cin(gnd),
	.combout(always1),
	.cout());
// synopsys translate_off
defparam \always1~0 .lut_mask = 16'h7F0F;
defparam \always1~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X50_Y33_N22
cycloneive_lcell_comb \ramif.ramload[0]~0 (
// Equation(s):
// ramiframload_0 = ((address_reg_a_0 & (ram_block3a321)) # (!address_reg_a_0 & ((ram_block3a01)))) # (!always1)

	.dataa(\altsyncram_component|auto_generated|altsyncram1|ram_block3a32~portadataout ),
	.datab(\altsyncram_component|auto_generated|altsyncram1|ram_block3a0~portadataout ),
	.datac(\altsyncram_component|auto_generated|altsyncram1|address_reg_a [0]),
	.datad(always1),
	.cin(gnd),
	.combout(ramiframload_0),
	.cout());
// synopsys translate_off
defparam \ramif.ramload[0]~0 .lut_mask = 16'hACFF;
defparam \ramif.ramload[0]~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y30_N24
cycloneive_lcell_comb \ramif.ramload[1]~1 (
// Equation(s):
// ramiframload_1 = (always1 & ((address_reg_a_0 & ((ram_block3a331))) # (!address_reg_a_0 & (ram_block3a110))))

	.dataa(\altsyncram_component|auto_generated|altsyncram1|address_reg_a [0]),
	.datab(always1),
	.datac(\altsyncram_component|auto_generated|altsyncram1|ram_block3a1~portadataout ),
	.datad(\altsyncram_component|auto_generated|altsyncram1|ram_block3a33~portadataout ),
	.cin(gnd),
	.combout(ramiframload_1),
	.cout());
// synopsys translate_off
defparam \ramif.ramload[1]~1 .lut_mask = 16'hC840;
defparam \ramif.ramload[1]~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y29_N20
cycloneive_lcell_comb \ramif.ramload[2]~2 (
// Equation(s):
// ramiframload_2 = (always1 & ((address_reg_a_0 & ((ram_block3a341))) # (!address_reg_a_0 & (ram_block3a210))))

	.dataa(\altsyncram_component|auto_generated|altsyncram1|address_reg_a [0]),
	.datab(always1),
	.datac(\altsyncram_component|auto_generated|altsyncram1|ram_block3a2~portadataout ),
	.datad(\altsyncram_component|auto_generated|altsyncram1|ram_block3a34~portadataout ),
	.cin(gnd),
	.combout(ramiframload_2),
	.cout());
// synopsys translate_off
defparam \ramif.ramload[2]~2 .lut_mask = 16'hC840;
defparam \ramif.ramload[2]~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y30_N6
cycloneive_lcell_comb \ramif.ramload[3]~3 (
// Equation(s):
// ramiframload_3 = (always1 & ((address_reg_a_0 & (ram_block3a351)) # (!address_reg_a_0 & ((ram_block3a310)))))

	.dataa(\altsyncram_component|auto_generated|altsyncram1|address_reg_a [0]),
	.datab(always1),
	.datac(\altsyncram_component|auto_generated|altsyncram1|ram_block3a35~portadataout ),
	.datad(\altsyncram_component|auto_generated|altsyncram1|ram_block3a3~portadataout ),
	.cin(gnd),
	.combout(ramiframload_3),
	.cout());
// synopsys translate_off
defparam \ramif.ramload[3]~3 .lut_mask = 16'hC480;
defparam \ramif.ramload[3]~3 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y33_N6
cycloneive_lcell_comb \ramif.ramload[4]~4 (
// Equation(s):
// ramiframload_4 = ((address_reg_a_0 & (ram_block3a361)) # (!address_reg_a_0 & ((ram_block3a410)))) # (!always1)

	.dataa(\altsyncram_component|auto_generated|altsyncram1|address_reg_a [0]),
	.datab(\altsyncram_component|auto_generated|altsyncram1|ram_block3a36~portadataout ),
	.datac(always1),
	.datad(\altsyncram_component|auto_generated|altsyncram1|ram_block3a4~portadataout ),
	.cin(gnd),
	.combout(ramiframload_4),
	.cout());
// synopsys translate_off
defparam \ramif.ramload[4]~4 .lut_mask = 16'hDF8F;
defparam \ramif.ramload[4]~4 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y30_N12
cycloneive_lcell_comb \ramif.ramload[5]~5 (
// Equation(s):
// ramiframload_5 = (always1 & ((address_reg_a_0 & ((ram_block3a371))) # (!address_reg_a_0 & (ram_block3a510))))

	.dataa(always1),
	.datab(\altsyncram_component|auto_generated|altsyncram1|address_reg_a [0]),
	.datac(\altsyncram_component|auto_generated|altsyncram1|ram_block3a5~portadataout ),
	.datad(\altsyncram_component|auto_generated|altsyncram1|ram_block3a37~portadataout ),
	.cin(gnd),
	.combout(ramiframload_5),
	.cout());
// synopsys translate_off
defparam \ramif.ramload[5]~5 .lut_mask = 16'hA820;
defparam \ramif.ramload[5]~5 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y30_N20
cycloneive_lcell_comb \ramif.ramload[6]~6 (
// Equation(s):
// ramiframload_6 = ((address_reg_a_0 & ((ram_block3a381))) # (!address_reg_a_0 & (ram_block3a64))) # (!always1)

	.dataa(\altsyncram_component|auto_generated|altsyncram1|address_reg_a [0]),
	.datab(always1),
	.datac(\altsyncram_component|auto_generated|altsyncram1|ram_block3a6~portadataout ),
	.datad(\altsyncram_component|auto_generated|altsyncram1|ram_block3a38~portadataout ),
	.cin(gnd),
	.combout(ramiframload_6),
	.cout());
// synopsys translate_off
defparam \ramif.ramload[6]~6 .lut_mask = 16'hFB73;
defparam \ramif.ramload[6]~6 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y30_N26
cycloneive_lcell_comb \ramif.ramload[7]~7 (
// Equation(s):
// ramiframload_7 = ((address_reg_a_0 & (ram_block3a391)) # (!address_reg_a_0 & ((ram_block3a71)))) # (!always1)

	.dataa(\altsyncram_component|auto_generated|altsyncram1|address_reg_a [0]),
	.datab(always1),
	.datac(\altsyncram_component|auto_generated|altsyncram1|ram_block3a39~portadataout ),
	.datad(\altsyncram_component|auto_generated|altsyncram1|ram_block3a7~portadataout ),
	.cin(gnd),
	.combout(ramiframload_7),
	.cout());
// synopsys translate_off
defparam \ramif.ramload[7]~7 .lut_mask = 16'hF7B3;
defparam \ramif.ramload[7]~7 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y29_N30
cycloneive_lcell_comb \ramif.ramload[8]~8 (
// Equation(s):
// ramiframload_8 = (always1 & ((address_reg_a_0 & (ram_block3a401)) # (!address_reg_a_0 & ((ram_block3a81)))))

	.dataa(\altsyncram_component|auto_generated|altsyncram1|address_reg_a [0]),
	.datab(always1),
	.datac(\altsyncram_component|auto_generated|altsyncram1|ram_block3a40~portadataout ),
	.datad(\altsyncram_component|auto_generated|altsyncram1|ram_block3a8~portadataout ),
	.cin(gnd),
	.combout(ramiframload_8),
	.cout());
// synopsys translate_off
defparam \ramif.ramload[8]~8 .lut_mask = 16'hC480;
defparam \ramif.ramload[8]~8 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y35_N16
cycloneive_lcell_comb \ramif.ramload[9]~9 (
// Equation(s):
// ramiframload_9 = ((address_reg_a_0 & ((ram_block3a412))) # (!address_reg_a_0 & (ram_block3a91))) # (!always1)

	.dataa(\altsyncram_component|auto_generated|altsyncram1|ram_block3a9~portadataout ),
	.datab(\altsyncram_component|auto_generated|altsyncram1|address_reg_a [0]),
	.datac(\altsyncram_component|auto_generated|altsyncram1|ram_block3a41~portadataout ),
	.datad(always1),
	.cin(gnd),
	.combout(ramiframload_9),
	.cout());
// synopsys translate_off
defparam \ramif.ramload[9]~9 .lut_mask = 16'hE2FF;
defparam \ramif.ramload[9]~9 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y30_N2
cycloneive_lcell_comb \ramif.ramload[10]~10 (
// Equation(s):
// ramiframload_10 = (always1 & ((address_reg_a_0 & ((ram_block3a421))) # (!address_reg_a_0 & (ram_block3a101))))

	.dataa(always1),
	.datab(\altsyncram_component|auto_generated|altsyncram1|address_reg_a [0]),
	.datac(\altsyncram_component|auto_generated|altsyncram1|ram_block3a10~portadataout ),
	.datad(\altsyncram_component|auto_generated|altsyncram1|ram_block3a42~portadataout ),
	.cin(gnd),
	.combout(ramiframload_10),
	.cout());
// synopsys translate_off
defparam \ramif.ramload[10]~10 .lut_mask = 16'hA820;
defparam \ramif.ramload[10]~10 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y29_N24
cycloneive_lcell_comb \ramif.ramload[11]~11 (
// Equation(s):
// ramiframload_11 = ((address_reg_a_0 & (ram_block3a431)) # (!address_reg_a_0 & ((ram_block3a112)))) # (!always1)

	.dataa(\altsyncram_component|auto_generated|altsyncram1|address_reg_a [0]),
	.datab(always1),
	.datac(\altsyncram_component|auto_generated|altsyncram1|ram_block3a43~portadataout ),
	.datad(\altsyncram_component|auto_generated|altsyncram1|ram_block3a11~portadataout ),
	.cin(gnd),
	.combout(ramiframload_11),
	.cout());
// synopsys translate_off
defparam \ramif.ramload[11]~11 .lut_mask = 16'hF7B3;
defparam \ramif.ramload[11]~11 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y34_N16
cycloneive_lcell_comb \ramif.ramload[12]~12 (
// Equation(s):
// ramiframload_12 = ((address_reg_a_0 & ((ram_block3a441))) # (!address_reg_a_0 & (ram_block3a121))) # (!always1)

	.dataa(\altsyncram_component|auto_generated|altsyncram1|address_reg_a [0]),
	.datab(always1),
	.datac(\altsyncram_component|auto_generated|altsyncram1|ram_block3a12~portadataout ),
	.datad(\altsyncram_component|auto_generated|altsyncram1|ram_block3a44~portadataout ),
	.cin(gnd),
	.combout(ramiframload_12),
	.cout());
// synopsys translate_off
defparam \ramif.ramload[12]~12 .lut_mask = 16'hFB73;
defparam \ramif.ramload[12]~12 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X50_Y33_N12
cycloneive_lcell_comb \ramif.ramload[13]~13 (
// Equation(s):
// ramiframload_13 = ((address_reg_a_0 & ((ram_block3a451))) # (!address_reg_a_0 & (ram_block3a131))) # (!always1)

	.dataa(\altsyncram_component|auto_generated|altsyncram1|address_reg_a [0]),
	.datab(always1),
	.datac(\altsyncram_component|auto_generated|altsyncram1|ram_block3a13~portadataout ),
	.datad(\altsyncram_component|auto_generated|altsyncram1|ram_block3a45~portadataout ),
	.cin(gnd),
	.combout(ramiframload_13),
	.cout());
// synopsys translate_off
defparam \ramif.ramload[13]~13 .lut_mask = 16'hFB73;
defparam \ramif.ramload[13]~13 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y30_N24
cycloneive_lcell_comb \ramif.ramload[14]~14 (
// Equation(s):
// ramiframload_14 = (always1 & ((address_reg_a_0 & (ram_block3a461)) # (!address_reg_a_0 & ((ram_block3a141)))))

	.dataa(\altsyncram_component|auto_generated|altsyncram1|address_reg_a [0]),
	.datab(always1),
	.datac(\altsyncram_component|auto_generated|altsyncram1|ram_block3a46~portadataout ),
	.datad(\altsyncram_component|auto_generated|altsyncram1|ram_block3a14~portadataout ),
	.cin(gnd),
	.combout(ramiframload_14),
	.cout());
// synopsys translate_off
defparam \ramif.ramload[14]~14 .lut_mask = 16'hC480;
defparam \ramif.ramload[14]~14 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y33_N0
cycloneive_lcell_comb \ramif.ramload[15]~15 (
// Equation(s):
// ramiframload_15 = ((address_reg_a_0 & ((ram_block3a471))) # (!address_reg_a_0 & (ram_block3a151))) # (!always1)

	.dataa(always1),
	.datab(\altsyncram_component|auto_generated|altsyncram1|address_reg_a [0]),
	.datac(\altsyncram_component|auto_generated|altsyncram1|ram_block3a15~portadataout ),
	.datad(\altsyncram_component|auto_generated|altsyncram1|ram_block3a47~portadataout ),
	.cin(gnd),
	.combout(ramiframload_15),
	.cout());
// synopsys translate_off
defparam \ramif.ramload[15]~15 .lut_mask = 16'hFD75;
defparam \ramif.ramload[15]~15 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y31_N28
cycloneive_lcell_comb \ramif.ramload[16]~16 (
// Equation(s):
// ramiframload_16 = ((address_reg_a_0 & (ram_block3a481)) # (!address_reg_a_0 & ((ram_block3a161)))) # (!always1)

	.dataa(always1),
	.datab(\altsyncram_component|auto_generated|altsyncram1|address_reg_a [0]),
	.datac(\altsyncram_component|auto_generated|altsyncram1|ram_block3a48~portadataout ),
	.datad(\altsyncram_component|auto_generated|altsyncram1|ram_block3a16~portadataout ),
	.cin(gnd),
	.combout(ramiframload_16),
	.cout());
// synopsys translate_off
defparam \ramif.ramload[16]~16 .lut_mask = 16'hF7D5;
defparam \ramif.ramload[16]~16 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y31_N14
cycloneive_lcell_comb \ramif.ramload[17]~17 (
// Equation(s):
// ramiframload_17 = (always1 & ((address_reg_a_0 & ((ram_block3a491))) # (!address_reg_a_0 & (ram_block3a171))))

	.dataa(always1),
	.datab(\altsyncram_component|auto_generated|altsyncram1|address_reg_a [0]),
	.datac(\altsyncram_component|auto_generated|altsyncram1|ram_block3a17~portadataout ),
	.datad(\altsyncram_component|auto_generated|altsyncram1|ram_block3a49~portadataout ),
	.cin(gnd),
	.combout(ramiframload_17),
	.cout());
// synopsys translate_off
defparam \ramif.ramload[17]~17 .lut_mask = 16'hA820;
defparam \ramif.ramload[17]~17 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y31_N16
cycloneive_lcell_comb \ramif.ramload[18]~18 (
// Equation(s):
// ramiframload_18 = (always1 & ((address_reg_a_0 & (ram_block3a501)) # (!address_reg_a_0 & ((ram_block3a181)))))

	.dataa(always1),
	.datab(\altsyncram_component|auto_generated|altsyncram1|address_reg_a [0]),
	.datac(\altsyncram_component|auto_generated|altsyncram1|ram_block3a50~portadataout ),
	.datad(\altsyncram_component|auto_generated|altsyncram1|ram_block3a18~portadataout ),
	.cin(gnd),
	.combout(ramiframload_18),
	.cout());
// synopsys translate_off
defparam \ramif.ramload[18]~18 .lut_mask = 16'hA280;
defparam \ramif.ramload[18]~18 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y33_N18
cycloneive_lcell_comb \ramif.ramload[19]~19 (
// Equation(s):
// ramiframload_19 = (always1 & ((address_reg_a_0 & (ram_block3a512)) # (!address_reg_a_0 & ((ram_block3a191)))))

	.dataa(always1),
	.datab(\altsyncram_component|auto_generated|altsyncram1|address_reg_a [0]),
	.datac(\altsyncram_component|auto_generated|altsyncram1|ram_block3a51~portadataout ),
	.datad(\altsyncram_component|auto_generated|altsyncram1|ram_block3a19~portadataout ),
	.cin(gnd),
	.combout(ramiframload_19),
	.cout());
// synopsys translate_off
defparam \ramif.ramload[19]~19 .lut_mask = 16'hA280;
defparam \ramif.ramload[19]~19 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y33_N16
cycloneive_lcell_comb \ramif.ramload[20]~20 (
// Equation(s):
// ramiframload_20 = ((address_reg_a_0 & ((ram_block3a521))) # (!address_reg_a_0 & (ram_block3a201))) # (!always1)

	.dataa(always1),
	.datab(\altsyncram_component|auto_generated|altsyncram1|address_reg_a [0]),
	.datac(\altsyncram_component|auto_generated|altsyncram1|ram_block3a20~portadataout ),
	.datad(\altsyncram_component|auto_generated|altsyncram1|ram_block3a52~portadataout ),
	.cin(gnd),
	.combout(ramiframload_20),
	.cout());
// synopsys translate_off
defparam \ramif.ramload[20]~20 .lut_mask = 16'hFD75;
defparam \ramif.ramload[20]~20 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y32_N16
cycloneive_lcell_comb \ramif.ramload[21]~21 (
// Equation(s):
// ramiframload_21 = (always1 & ((address_reg_a_0 & (ram_block3a531)) # (!address_reg_a_0 & ((ram_block3a212)))))

	.dataa(\altsyncram_component|auto_generated|altsyncram1|address_reg_a [0]),
	.datab(always1),
	.datac(\altsyncram_component|auto_generated|altsyncram1|ram_block3a53~portadataout ),
	.datad(\altsyncram_component|auto_generated|altsyncram1|ram_block3a21~portadataout ),
	.cin(gnd),
	.combout(ramiframload_21),
	.cout());
// synopsys translate_off
defparam \ramif.ramload[21]~21 .lut_mask = 16'hC480;
defparam \ramif.ramload[21]~21 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y32_N14
cycloneive_lcell_comb \ramif.ramload[22]~22 (
// Equation(s):
// ramiframload_22 = ((address_reg_a_0 & (ram_block3a541)) # (!address_reg_a_0 & ((ram_block3a221)))) # (!always1)

	.dataa(\altsyncram_component|auto_generated|altsyncram1|address_reg_a [0]),
	.datab(always1),
	.datac(\altsyncram_component|auto_generated|altsyncram1|ram_block3a54~portadataout ),
	.datad(\altsyncram_component|auto_generated|altsyncram1|ram_block3a22~portadataout ),
	.cin(gnd),
	.combout(ramiframload_22),
	.cout());
// synopsys translate_off
defparam \ramif.ramload[22]~22 .lut_mask = 16'hF7B3;
defparam \ramif.ramload[22]~22 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y32_N24
cycloneive_lcell_comb \ramif.ramload[23]~23 (
// Equation(s):
// ramiframload_23 = ((address_reg_a_0 & (ram_block3a551)) # (!address_reg_a_0 & ((ram_block3a231)))) # (!always1)

	.dataa(\altsyncram_component|auto_generated|altsyncram1|address_reg_a [0]),
	.datab(\altsyncram_component|auto_generated|altsyncram1|ram_block3a55~portadataout ),
	.datac(always1),
	.datad(\altsyncram_component|auto_generated|altsyncram1|ram_block3a23~portadataout ),
	.cin(gnd),
	.combout(ramiframload_23),
	.cout());
// synopsys translate_off
defparam \ramif.ramload[23]~23 .lut_mask = 16'hDF8F;
defparam \ramif.ramload[23]~23 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y32_N22
cycloneive_lcell_comb \ramif.ramload[24]~24 (
// Equation(s):
// ramiframload_24 = (always1 & ((address_reg_a_0 & ((ram_block3a561))) # (!address_reg_a_0 & (ram_block3a241))))

	.dataa(\altsyncram_component|auto_generated|altsyncram1|address_reg_a [0]),
	.datab(\altsyncram_component|auto_generated|altsyncram1|ram_block3a24~portadataout ),
	.datac(always1),
	.datad(\altsyncram_component|auto_generated|altsyncram1|ram_block3a56~portadataout ),
	.cin(gnd),
	.combout(ramiframload_24),
	.cout());
// synopsys translate_off
defparam \ramif.ramload[24]~24 .lut_mask = 16'hE040;
defparam \ramif.ramload[24]~24 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y33_N14
cycloneive_lcell_comb \ramif.ramload[25]~25 (
// Equation(s):
// ramiframload_25 = ((address_reg_a_0 & ((ram_block3a571))) # (!address_reg_a_0 & (ram_block3a251))) # (!always1)

	.dataa(always1),
	.datab(\altsyncram_component|auto_generated|altsyncram1|address_reg_a [0]),
	.datac(\altsyncram_component|auto_generated|altsyncram1|ram_block3a25~portadataout ),
	.datad(\altsyncram_component|auto_generated|altsyncram1|ram_block3a57~portadataout ),
	.cin(gnd),
	.combout(ramiframload_25),
	.cout());
// synopsys translate_off
defparam \ramif.ramload[25]~25 .lut_mask = 16'hFD75;
defparam \ramif.ramload[25]~25 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y30_N16
cycloneive_lcell_comb \ramif.ramload[26]~26 (
// Equation(s):
// ramiframload_26 = (always1 & ((address_reg_a_0 & (ram_block3a581)) # (!address_reg_a_0 & ((ram_block3a261)))))

	.dataa(always1),
	.datab(\altsyncram_component|auto_generated|altsyncram1|address_reg_a [0]),
	.datac(\altsyncram_component|auto_generated|altsyncram1|ram_block3a58~portadataout ),
	.datad(\altsyncram_component|auto_generated|altsyncram1|ram_block3a26~portadataout ),
	.cin(gnd),
	.combout(ramiframload_26),
	.cout());
// synopsys translate_off
defparam \ramif.ramload[26]~26 .lut_mask = 16'hA280;
defparam \ramif.ramload[26]~26 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y30_N22
cycloneive_lcell_comb \ramif.ramload[27]~27 (
// Equation(s):
// ramiframload_27 = ((address_reg_a_0 & (ram_block3a591)) # (!address_reg_a_0 & ((ram_block3a271)))) # (!always1)

	.dataa(\altsyncram_component|auto_generated|altsyncram1|address_reg_a [0]),
	.datab(always1),
	.datac(\altsyncram_component|auto_generated|altsyncram1|ram_block3a59~portadataout ),
	.datad(\altsyncram_component|auto_generated|altsyncram1|ram_block3a27~portadataout ),
	.cin(gnd),
	.combout(ramiframload_27),
	.cout());
// synopsys translate_off
defparam \ramif.ramload[27]~27 .lut_mask = 16'hF7B3;
defparam \ramif.ramload[27]~27 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y30_N10
cycloneive_lcell_comb \ramif.ramload[28]~28 (
// Equation(s):
// ramiframload_28 = ((address_reg_a_0 & (ram_block3a601)) # (!address_reg_a_0 & ((ram_block3a281)))) # (!always1)

	.dataa(always1),
	.datab(\altsyncram_component|auto_generated|altsyncram1|address_reg_a [0]),
	.datac(\altsyncram_component|auto_generated|altsyncram1|ram_block3a60~portadataout ),
	.datad(\altsyncram_component|auto_generated|altsyncram1|ram_block3a28~portadataout ),
	.cin(gnd),
	.combout(ramiframload_28),
	.cout());
// synopsys translate_off
defparam \ramif.ramload[28]~28 .lut_mask = 16'hF7D5;
defparam \ramif.ramload[28]~28 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y33_N20
cycloneive_lcell_comb \ramif.ramload[29]~29 (
// Equation(s):
// ramiframload_29 = ((address_reg_a_0 & ((ram_block3a611))) # (!address_reg_a_0 & (ram_block3a291))) # (!always1)

	.dataa(always1),
	.datab(\altsyncram_component|auto_generated|altsyncram1|address_reg_a [0]),
	.datac(\altsyncram_component|auto_generated|altsyncram1|ram_block3a29~portadataout ),
	.datad(\altsyncram_component|auto_generated|altsyncram1|ram_block3a61~portadataout ),
	.cin(gnd),
	.combout(ramiframload_29),
	.cout());
// synopsys translate_off
defparam \ramif.ramload[29]~29 .lut_mask = 16'hFD75;
defparam \ramif.ramload[29]~29 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y30_N12
cycloneive_lcell_comb \ramif.ramload[30]~30 (
// Equation(s):
// ramiframload_30 = (always1 & ((address_reg_a_0 & ((ram_block3a621))) # (!address_reg_a_0 & (ram_block3a301))))

	.dataa(\altsyncram_component|auto_generated|altsyncram1|address_reg_a [0]),
	.datab(always1),
	.datac(\altsyncram_component|auto_generated|altsyncram1|ram_block3a30~portadataout ),
	.datad(\altsyncram_component|auto_generated|altsyncram1|ram_block3a62~portadataout ),
	.cin(gnd),
	.combout(ramiframload_30),
	.cout());
// synopsys translate_off
defparam \ramif.ramload[30]~30 .lut_mask = 16'hC840;
defparam \ramif.ramload[30]~30 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y30_N10
cycloneive_lcell_comb \ramif.ramload[31]~31 (
// Equation(s):
// ramiframload_31 = ((address_reg_a_0 & (ram_block3a631)) # (!address_reg_a_0 & ((ram_block3a312)))) # (!always1)

	.dataa(\altsyncram_component|auto_generated|altsyncram1|address_reg_a [0]),
	.datab(\altsyncram_component|auto_generated|altsyncram1|ram_block3a63~portadataout ),
	.datac(\altsyncram_component|auto_generated|altsyncram1|ram_block3a31~portadataout ),
	.datad(always1),
	.cin(gnd),
	.combout(ramiframload_31),
	.cout());
// synopsys translate_off
defparam \ramif.ramload[31]~31 .lut_mask = 16'hD8FF;
defparam \ramif.ramload[31]~31 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y34_N18
cycloneive_lcell_comb \addr[7]~feeder (
// Equation(s):
// \addr[7]~feeder_combout  = \ramaddr~11_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(ramaddr6),
	.cin(gnd),
	.combout(\addr[7]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \addr[7]~feeder .lut_mask = 16'hFF00;
defparam \addr[7]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X54_Y34_N29
dffeas \en[1] (
	.clk(CLK),
	.d(\ramif.ramREN ),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~1_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(en[1]),
	.prn(vcc));
// synopsys translate_off
defparam \en[1] .is_wysiwyg = "true";
defparam \en[1] .power_up = "low";
// synopsys translate_on

// Location: FF_X54_Y34_N11
dffeas \en[0] (
	.clk(CLK),
	.d(\ramif.ramWEN ),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~1_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(en[0]),
	.prn(vcc));
// synopsys translate_off
defparam \en[0] .is_wysiwyg = "true";
defparam \en[0] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X54_Y34_N12
cycloneive_lcell_comb \always0~0 (
// Equation(s):
// \always0~0_combout  = (\ramWEN~0_combout  & ((en[1] $ (\ramREN~1_combout )) # (!en[0]))) # (!\ramWEN~0_combout  & ((en[0]) # (en[1] $ (\ramREN~1_combout ))))

	.dataa(\ramif.ramWEN ),
	.datab(en[1]),
	.datac(en[0]),
	.datad(\ramif.ramREN ),
	.cin(gnd),
	.combout(\always0~0_combout ),
	.cout());
// synopsys translate_off
defparam \always0~0 .lut_mask = 16'h7BDE;
defparam \always0~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y34_N26
cycloneive_lcell_comb \always0~1 (
// Equation(s):
// \always0~1_combout  = ((\always0~0_combout ) # ((\ramWEN~0_combout  & \ramREN~1_combout ))) # (!\Equal2~22_combout )

	.dataa(\ramif.ramWEN ),
	.datab(\Equal2~22_combout ),
	.datac(\always0~0_combout ),
	.datad(\ramif.ramREN ),
	.cin(gnd),
	.combout(\always0~1_combout ),
	.cout());
// synopsys translate_off
defparam \always0~1 .lut_mask = 16'hFBF3;
defparam \always0~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X55_Y34_N19
dffeas \addr[7] (
	.clk(CLK),
	.d(\addr[7]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~1_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(addr[7]),
	.prn(vcc));
// synopsys translate_off
defparam \addr[7] .is_wysiwyg = "true";
defparam \addr[7] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X55_Y34_N12
cycloneive_lcell_comb \addr[6]~feeder (
// Equation(s):
// \addr[6]~feeder_combout  = \ramaddr~13_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(ramaddr7),
	.cin(gnd),
	.combout(\addr[6]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \addr[6]~feeder .lut_mask = 16'hFF00;
defparam \addr[6]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X55_Y34_N13
dffeas \addr[6] (
	.clk(CLK),
	.d(\addr[6]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~1_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(addr[6]),
	.prn(vcc));
// synopsys translate_off
defparam \addr[6] .is_wysiwyg = "true";
defparam \addr[6] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X55_Y34_N8
cycloneive_lcell_comb \Equal2~5 (
// Equation(s):
// \Equal2~5_combout  = (\ramaddr~13_combout  & (addr[6] & (addr[7] $ (!\ramaddr~11_combout )))) # (!\ramaddr~13_combout  & (!addr[6] & (addr[7] $ (!\ramaddr~11_combout ))))

	.dataa(ramaddr7),
	.datab(addr[7]),
	.datac(addr[6]),
	.datad(ramaddr6),
	.cin(gnd),
	.combout(\Equal2~5_combout ),
	.cout());
// synopsys translate_off
defparam \Equal2~5 .lut_mask = 16'h8421;
defparam \Equal2~5 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y35_N16
cycloneive_lcell_comb \addr[2]~feeder (
// Equation(s):
// \addr[2]~feeder_combout  = \ramaddr~5_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(ramaddr3),
	.cin(gnd),
	.combout(\addr[2]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \addr[2]~feeder .lut_mask = 16'hFF00;
defparam \addr[2]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X54_Y35_N17
dffeas \addr[2] (
	.clk(CLK),
	.d(\addr[2]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~1_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(addr[2]),
	.prn(vcc));
// synopsys translate_off
defparam \addr[2] .is_wysiwyg = "true";
defparam \addr[2] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X54_Y35_N24
cycloneive_lcell_comb \Equal2~3 (
// Equation(s):
// \Equal2~3_combout  = (addr[3] & (\ramaddr~3_combout  & (addr[2] $ (!\ramaddr~5_combout )))) # (!addr[3] & (!\ramaddr~3_combout  & (addr[2] $ (!\ramaddr~5_combout ))))

	.dataa(addr[3]),
	.datab(addr[2]),
	.datac(ramaddr3),
	.datad(ramaddr2),
	.cin(gnd),
	.combout(\Equal2~3_combout ),
	.cout());
// synopsys translate_off
defparam \Equal2~3 .lut_mask = 16'h8241;
defparam \Equal2~3 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X49_Y34_N8
cycloneive_lcell_comb \addr[5]~feeder (
// Equation(s):
// \addr[5]~feeder_combout  = \ramaddr~7_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(ramaddr4),
	.cin(gnd),
	.combout(\addr[5]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \addr[5]~feeder .lut_mask = 16'hFF00;
defparam \addr[5]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X49_Y34_N9
dffeas \addr[5] (
	.clk(CLK),
	.d(\addr[5]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~1_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(addr[5]),
	.prn(vcc));
// synopsys translate_off
defparam \addr[5] .is_wysiwyg = "true";
defparam \addr[5] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X49_Y34_N10
cycloneive_lcell_comb \Equal2~4 (
// Equation(s):
// \Equal2~4_combout  = (addr[4] & (\ramaddr~9_combout  & (addr[5] $ (!\ramaddr~7_combout )))) # (!addr[4] & (!\ramaddr~9_combout  & (addr[5] $ (!\ramaddr~7_combout ))))

	.dataa(addr[4]),
	.datab(ramaddr5),
	.datac(addr[5]),
	.datad(ramaddr4),
	.cin(gnd),
	.combout(\Equal2~4_combout ),
	.cout());
// synopsys translate_off
defparam \Equal2~4 .lut_mask = 16'h9009;
defparam \Equal2~4 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y34_N30
cycloneive_lcell_comb \Equal2~6 (
// Equation(s):
// \Equal2~6_combout  = (\Equal2~2_combout  & (\Equal2~5_combout  & (\Equal2~3_combout  & \Equal2~4_combout )))

	.dataa(\Equal2~2_combout ),
	.datab(\Equal2~5_combout ),
	.datac(\Equal2~3_combout ),
	.datad(\Equal2~4_combout ),
	.cin(gnd),
	.combout(\Equal2~6_combout ),
	.cout());
// synopsys translate_off
defparam \Equal2~6 .lut_mask = 16'h8000;
defparam \Equal2~6 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X54_Y37_N13
dffeas \addr[10] (
	.clk(CLK),
	.d(ramaddr11),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~1_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(addr[10]),
	.prn(vcc));
// synopsys translate_off
defparam \addr[10] .is_wysiwyg = "true";
defparam \addr[10] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X54_Y37_N28
cycloneive_lcell_comb \Equal2~8 (
// Equation(s):
// \Equal2~8_combout  = (addr[11] & (\ramaddr~19_combout  & (addr[10] $ (!\ramaddr~21_combout )))) # (!addr[11] & (!\ramaddr~19_combout  & (addr[10] $ (!\ramaddr~21_combout ))))

	.dataa(addr[11]),
	.datab(addr[10]),
	.datac(ramaddr10),
	.datad(ramaddr11),
	.cin(gnd),
	.combout(\Equal2~8_combout ),
	.cout());
// synopsys translate_off
defparam \Equal2~8 .lut_mask = 16'h8421;
defparam \Equal2~8 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X54_Y33_N11
dffeas \addr[9] (
	.clk(CLK),
	.d(ramaddr8),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~1_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(addr[9]),
	.prn(vcc));
// synopsys translate_off
defparam \addr[9] .is_wysiwyg = "true";
defparam \addr[9] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X54_Y33_N26
cycloneive_lcell_comb \Equal2~7 (
// Equation(s):
// \Equal2~7_combout  = (addr[8] & (\ramaddr~17_combout  & (addr[9] $ (!\ramaddr~15_combout )))) # (!addr[8] & (!\ramaddr~17_combout  & (addr[9] $ (!\ramaddr~15_combout ))))

	.dataa(addr[8]),
	.datab(addr[9]),
	.datac(ramaddr9),
	.datad(ramaddr8),
	.cin(gnd),
	.combout(\Equal2~7_combout ),
	.cout());
// synopsys translate_off
defparam \Equal2~7 .lut_mask = 16'h8421;
defparam \Equal2~7 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y32_N4
cycloneive_lcell_comb \addr[12]~feeder (
// Equation(s):
// \addr[12]~feeder_combout  = \ramaddr~25_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(ramaddr13),
	.datad(gnd),
	.cin(gnd),
	.combout(\addr[12]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \addr[12]~feeder .lut_mask = 16'hF0F0;
defparam \addr[12]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X54_Y32_N5
dffeas \addr[12] (
	.clk(CLK),
	.d(\addr[12]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~1_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(addr[12]),
	.prn(vcc));
// synopsys translate_off
defparam \addr[12] .is_wysiwyg = "true";
defparam \addr[12] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X54_Y32_N20
cycloneive_lcell_comb \Equal2~9 (
// Equation(s):
// \Equal2~9_combout  = (addr[13] & (\ramaddr~23_combout  & (\ramaddr~25_combout  $ (!addr[12])))) # (!addr[13] & (!\ramaddr~23_combout  & (\ramaddr~25_combout  $ (!addr[12]))))

	.dataa(addr[13]),
	.datab(ramaddr13),
	.datac(addr[12]),
	.datad(ramaddr12),
	.cin(gnd),
	.combout(\Equal2~9_combout ),
	.cout());
// synopsys translate_off
defparam \Equal2~9 .lut_mask = 16'h8241;
defparam \Equal2~9 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y34_N24
cycloneive_lcell_comb \Equal2~11 (
// Equation(s):
// \Equal2~11_combout  = (\Equal2~10_combout  & (\Equal2~8_combout  & (\Equal2~7_combout  & \Equal2~9_combout )))

	.dataa(\Equal2~10_combout ),
	.datab(\Equal2~8_combout ),
	.datac(\Equal2~7_combout ),
	.datad(\Equal2~9_combout ),
	.cin(gnd),
	.combout(\Equal2~11_combout ),
	.cout());
// synopsys translate_off
defparam \Equal2~11 .lut_mask = 16'h8000;
defparam \Equal2~11 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X54_Y34_N17
dffeas \addr[26] (
	.clk(CLK),
	.d(\ramif.ramaddr [26]),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~1_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(addr[26]),
	.prn(vcc));
// synopsys translate_off
defparam \addr[26] .is_wysiwyg = "true";
defparam \addr[26] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X54_Y34_N4
cycloneive_lcell_comb \Equal2~18 (
// Equation(s):
// \Equal2~18_combout  = (addr[27] & (\ramaddr~51_combout  & (\ramaddr~53_combout  $ (!addr[26])))) # (!addr[27] & (!\ramaddr~51_combout  & (\ramaddr~53_combout  $ (!addr[26]))))

	.dataa(addr[27]),
	.datab(\ramif.ramaddr [26]),
	.datac(addr[26]),
	.datad(\ramif.ramaddr [27]),
	.cin(gnd),
	.combout(\Equal2~18_combout ),
	.cout());
// synopsys translate_off
defparam \Equal2~18 .lut_mask = 16'h8241;
defparam \Equal2~18 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X50_Y34_N13
dffeas \addr[29] (
	.clk(CLK),
	.d(\ramif.ramaddr [29]),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~1_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(addr[29]),
	.prn(vcc));
// synopsys translate_off
defparam \addr[29] .is_wysiwyg = "true";
defparam \addr[29] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X50_Y34_N28
cycloneive_lcell_comb \Equal2~19 (
// Equation(s):
// \Equal2~19_combout  = (addr[28] & (\ramaddr~57_combout  & (addr[29] $ (!\ramaddr~55_combout )))) # (!addr[28] & (!\ramaddr~57_combout  & (addr[29] $ (!\ramaddr~55_combout ))))

	.dataa(addr[28]),
	.datab(addr[29]),
	.datac(ramaddr19),
	.datad(\ramif.ramaddr [29]),
	.cin(gnd),
	.combout(\Equal2~19_combout ),
	.cout());
// synopsys translate_off
defparam \Equal2~19 .lut_mask = 16'h8421;
defparam \Equal2~19 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X53_Y34_N3
dffeas \addr[31] (
	.clk(CLK),
	.d(\ramif.ramaddr [31]),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~1_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(addr[31]),
	.prn(vcc));
// synopsys translate_off
defparam \addr[31] .is_wysiwyg = "true";
defparam \addr[31] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X53_Y34_N30
cycloneive_lcell_comb \Equal2~20 (
// Equation(s):
// \Equal2~20_combout  = (addr[30] & (\ramaddr~61_combout  & (\ramaddr~59_combout  $ (!addr[31])))) # (!addr[30] & (!\ramaddr~61_combout  & (\ramaddr~59_combout  $ (!addr[31]))))

	.dataa(addr[30]),
	.datab(\ramif.ramaddr [31]),
	.datac(addr[31]),
	.datad(\ramif.ramaddr [30]),
	.cin(gnd),
	.combout(\Equal2~20_combout ),
	.cout());
// synopsys translate_off
defparam \Equal2~20 .lut_mask = 16'h8241;
defparam \Equal2~20 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y34_N14
cycloneive_lcell_comb \Equal2~21 (
// Equation(s):
// \Equal2~21_combout  = (\Equal2~17_combout  & (\Equal2~18_combout  & (\Equal2~19_combout  & \Equal2~20_combout )))

	.dataa(\Equal2~17_combout ),
	.datab(\Equal2~18_combout ),
	.datac(\Equal2~19_combout ),
	.datad(\Equal2~20_combout ),
	.cin(gnd),
	.combout(\Equal2~21_combout ),
	.cout());
// synopsys translate_off
defparam \Equal2~21 .lut_mask = 16'h8000;
defparam \Equal2~21 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X53_Y34_N19
dffeas \addr[23] (
	.clk(CLK),
	.d(\ramif.ramaddr [23]),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~1_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(addr[23]),
	.prn(vcc));
// synopsys translate_off
defparam \addr[23] .is_wysiwyg = "true";
defparam \addr[23] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X53_Y34_N4
cycloneive_lcell_comb \Equal2~15 (
// Equation(s):
// \Equal2~15_combout  = (addr[22] & (\ramaddr~45_combout  & (addr[23] $ (!\ramaddr~43_combout )))) # (!addr[22] & (!\ramaddr~45_combout  & (addr[23] $ (!\ramaddr~43_combout ))))

	.dataa(addr[22]),
	.datab(addr[23]),
	.datac(\ramif.ramaddr [22]),
	.datad(\ramif.ramaddr [23]),
	.cin(gnd),
	.combout(\Equal2~15_combout ),
	.cout());
// synopsys translate_off
defparam \Equal2~15 .lut_mask = 16'h8421;
defparam \Equal2~15 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X53_Y34_N11
dffeas \addr[21] (
	.clk(CLK),
	.d(\ramif.ramaddr [21]),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~1_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(addr[21]),
	.prn(vcc));
// synopsys translate_off
defparam \addr[21] .is_wysiwyg = "true";
defparam \addr[21] .power_up = "low";
// synopsys translate_on

// Location: FF_X53_Y34_N1
dffeas \addr[20] (
	.clk(CLK),
	.d(\ramif.ramaddr [20]),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~1_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(addr[20]),
	.prn(vcc));
// synopsys translate_off
defparam \addr[20] .is_wysiwyg = "true";
defparam \addr[20] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X53_Y34_N26
cycloneive_lcell_comb \Equal2~14 (
// Equation(s):
// \Equal2~14_combout  = (\ramaddr~39_combout  & (addr[21] & (addr[20] $ (!\ramaddr~41_combout )))) # (!\ramaddr~39_combout  & (!addr[21] & (addr[20] $ (!\ramaddr~41_combout ))))

	.dataa(\ramif.ramaddr [21]),
	.datab(addr[21]),
	.datac(addr[20]),
	.datad(\ramif.ramaddr [20]),
	.cin(gnd),
	.combout(\Equal2~14_combout ),
	.cout());
// synopsys translate_off
defparam \Equal2~14 .lut_mask = 16'h9009;
defparam \Equal2~14 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X50_Y34_N11
dffeas \addr[17] (
	.clk(CLK),
	.d(\ramif.ramaddr [17]),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~1_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(addr[17]),
	.prn(vcc));
// synopsys translate_off
defparam \addr[17] .is_wysiwyg = "true";
defparam \addr[17] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X50_Y34_N24
cycloneive_lcell_comb \Equal2~12 (
// Equation(s):
// \Equal2~12_combout  = (addr[16] & (\ramaddr~33_combout  & (addr[17] $ (!\ramaddr~31_combout )))) # (!addr[16] & (!\ramaddr~33_combout  & (addr[17] $ (!\ramaddr~31_combout ))))

	.dataa(addr[16]),
	.datab(\ramif.ramaddr [16]),
	.datac(addr[17]),
	.datad(\ramif.ramaddr [17]),
	.cin(gnd),
	.combout(\Equal2~12_combout ),
	.cout());
// synopsys translate_off
defparam \Equal2~12 .lut_mask = 16'h9009;
defparam \Equal2~12 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y34_N18
cycloneive_lcell_comb \Equal2~16 (
// Equation(s):
// \Equal2~16_combout  = (\Equal2~13_combout  & (\Equal2~15_combout  & (\Equal2~14_combout  & \Equal2~12_combout )))

	.dataa(\Equal2~13_combout ),
	.datab(\Equal2~15_combout ),
	.datac(\Equal2~14_combout ),
	.datad(\Equal2~12_combout ),
	.cin(gnd),
	.combout(\Equal2~16_combout ),
	.cout());
// synopsys translate_off
defparam \Equal2~16 .lut_mask = 16'h8000;
defparam \Equal2~16 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y34_N0
cycloneive_lcell_comb \Equal2~22 (
// Equation(s):
// \Equal2~22_combout  = (\Equal2~6_combout  & (\Equal2~11_combout  & (\Equal2~21_combout  & \Equal2~16_combout )))

	.dataa(\Equal2~6_combout ),
	.datab(\Equal2~11_combout ),
	.datac(\Equal2~21_combout ),
	.datad(\Equal2~16_combout ),
	.cin(gnd),
	.combout(\Equal2~22_combout ),
	.cout());
// synopsys translate_off
defparam \Equal2~22 .lut_mask = 16'h8000;
defparam \Equal2~22 .sum_lutc_input = "datac";
// synopsys translate_on

endmodule

module altsyncram_1 (
	ram_block3a32,
	ram_block3a0,
	ram_block3a33,
	ram_block3a1,
	ram_block3a34,
	ram_block3a2,
	ram_block3a35,
	ram_block3a3,
	ram_block3a36,
	ram_block3a4,
	ram_block3a37,
	ram_block3a5,
	ram_block3a38,
	ram_block3a6,
	ram_block3a39,
	ram_block3a7,
	ram_block3a40,
	ram_block3a8,
	ram_block3a41,
	ram_block3a9,
	ram_block3a42,
	ram_block3a10,
	ram_block3a43,
	ram_block3a11,
	ram_block3a44,
	ram_block3a12,
	ram_block3a45,
	ram_block3a13,
	ram_block3a46,
	ram_block3a14,
	ram_block3a47,
	ram_block3a15,
	ram_block3a48,
	ram_block3a16,
	ram_block3a49,
	ram_block3a17,
	ram_block3a50,
	ram_block3a18,
	ram_block3a51,
	ram_block3a19,
	ram_block3a52,
	ram_block3a20,
	ram_block3a53,
	ram_block3a21,
	ram_block3a54,
	ram_block3a22,
	ram_block3a55,
	ram_block3a23,
	ram_block3a56,
	ram_block3a24,
	ram_block3a57,
	ram_block3a25,
	ram_block3a58,
	ram_block3a26,
	ram_block3a59,
	ram_block3a27,
	ram_block3a60,
	ram_block3a28,
	ram_block3a61,
	ram_block3a29,
	ram_block3a62,
	ram_block3a30,
	ram_block3a63,
	ram_block3a31,
	is_in_use_reg,
	address_reg_a_0,
	address_a,
	ramaddr,
	ramWEN,
	always1,
	ir_loaded_address_reg_0,
	ir_loaded_address_reg_1,
	ir_loaded_address_reg_2,
	ir_loaded_address_reg_3,
	tdo,
	data_a,
	altera_internal_jtag,
	state_4,
	irf_reg_0_1,
	irf_reg_1_1,
	irf_reg_2_1,
	irf_reg_3_1,
	irf_reg_4_1,
	node_ena_1,
	clr_reg,
	virtual_ir_scan_reg,
	state_3,
	state_5,
	state_8,
	altera_internal_jtag1,
	clock0,
	devpor,
	devclrn,
	devoe);
output 	ram_block3a32;
output 	ram_block3a0;
output 	ram_block3a33;
output 	ram_block3a1;
output 	ram_block3a34;
output 	ram_block3a2;
output 	ram_block3a35;
output 	ram_block3a3;
output 	ram_block3a36;
output 	ram_block3a4;
output 	ram_block3a37;
output 	ram_block3a5;
output 	ram_block3a38;
output 	ram_block3a6;
output 	ram_block3a39;
output 	ram_block3a7;
output 	ram_block3a40;
output 	ram_block3a8;
output 	ram_block3a41;
output 	ram_block3a9;
output 	ram_block3a42;
output 	ram_block3a10;
output 	ram_block3a43;
output 	ram_block3a11;
output 	ram_block3a44;
output 	ram_block3a12;
output 	ram_block3a45;
output 	ram_block3a13;
output 	ram_block3a46;
output 	ram_block3a14;
output 	ram_block3a47;
output 	ram_block3a15;
output 	ram_block3a48;
output 	ram_block3a16;
output 	ram_block3a49;
output 	ram_block3a17;
output 	ram_block3a50;
output 	ram_block3a18;
output 	ram_block3a51;
output 	ram_block3a19;
output 	ram_block3a52;
output 	ram_block3a20;
output 	ram_block3a53;
output 	ram_block3a21;
output 	ram_block3a54;
output 	ram_block3a22;
output 	ram_block3a55;
output 	ram_block3a23;
output 	ram_block3a56;
output 	ram_block3a24;
output 	ram_block3a57;
output 	ram_block3a25;
output 	ram_block3a58;
output 	ram_block3a26;
output 	ram_block3a59;
output 	ram_block3a27;
output 	ram_block3a60;
output 	ram_block3a28;
output 	ram_block3a61;
output 	ram_block3a29;
output 	ram_block3a62;
output 	ram_block3a30;
output 	ram_block3a63;
output 	ram_block3a31;
output 	is_in_use_reg;
output 	address_reg_a_0;
input 	[13:0] address_a;
input 	ramaddr;
input 	ramWEN;
input 	always1;
output 	ir_loaded_address_reg_0;
output 	ir_loaded_address_reg_1;
output 	ir_loaded_address_reg_2;
output 	ir_loaded_address_reg_3;
output 	tdo;
input 	[31:0] data_a;
input 	altera_internal_jtag;
input 	state_4;
input 	irf_reg_0_1;
input 	irf_reg_1_1;
input 	irf_reg_2_1;
input 	irf_reg_3_1;
input 	irf_reg_4_1;
input 	node_ena_1;
input 	clr_reg;
input 	virtual_ir_scan_reg;
input 	state_3;
input 	state_5;
input 	state_8;
input 	altera_internal_jtag1;
input 	clock0;

// Design Ports Information

input 	devpor;
input 	devclrn;
input 	devoe;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
assign unknown = 1'bx;



altsyncram_99f1 auto_generated(
	.ram_block3a32(ram_block3a32),
	.ram_block3a0(ram_block3a0),
	.ram_block3a33(ram_block3a33),
	.ram_block3a1(ram_block3a1),
	.ram_block3a34(ram_block3a34),
	.ram_block3a2(ram_block3a2),
	.ram_block3a35(ram_block3a35),
	.ram_block3a3(ram_block3a3),
	.ram_block3a36(ram_block3a36),
	.ram_block3a4(ram_block3a4),
	.ram_block3a37(ram_block3a37),
	.ram_block3a5(ram_block3a5),
	.ram_block3a38(ram_block3a38),
	.ram_block3a6(ram_block3a6),
	.ram_block3a39(ram_block3a39),
	.ram_block3a7(ram_block3a7),
	.ram_block3a40(ram_block3a40),
	.ram_block3a8(ram_block3a8),
	.ram_block3a41(ram_block3a41),
	.ram_block3a9(ram_block3a9),
	.ram_block3a42(ram_block3a42),
	.ram_block3a10(ram_block3a10),
	.ram_block3a43(ram_block3a43),
	.ram_block3a11(ram_block3a11),
	.ram_block3a44(ram_block3a44),
	.ram_block3a12(ram_block3a12),
	.ram_block3a45(ram_block3a45),
	.ram_block3a13(ram_block3a13),
	.ram_block3a46(ram_block3a46),
	.ram_block3a14(ram_block3a14),
	.ram_block3a47(ram_block3a47),
	.ram_block3a15(ram_block3a15),
	.ram_block3a48(ram_block3a48),
	.ram_block3a16(ram_block3a16),
	.ram_block3a49(ram_block3a49),
	.ram_block3a17(ram_block3a17),
	.ram_block3a50(ram_block3a50),
	.ram_block3a18(ram_block3a18),
	.ram_block3a51(ram_block3a51),
	.ram_block3a19(ram_block3a19),
	.ram_block3a52(ram_block3a52),
	.ram_block3a20(ram_block3a20),
	.ram_block3a53(ram_block3a53),
	.ram_block3a21(ram_block3a21),
	.ram_block3a54(ram_block3a54),
	.ram_block3a22(ram_block3a22),
	.ram_block3a55(ram_block3a55),
	.ram_block3a23(ram_block3a23),
	.ram_block3a56(ram_block3a56),
	.ram_block3a24(ram_block3a24),
	.ram_block3a57(ram_block3a57),
	.ram_block3a25(ram_block3a25),
	.ram_block3a58(ram_block3a58),
	.ram_block3a26(ram_block3a26),
	.ram_block3a59(ram_block3a59),
	.ram_block3a27(ram_block3a27),
	.ram_block3a60(ram_block3a60),
	.ram_block3a28(ram_block3a28),
	.ram_block3a61(ram_block3a61),
	.ram_block3a29(ram_block3a29),
	.ram_block3a62(ram_block3a62),
	.ram_block3a30(ram_block3a30),
	.ram_block3a63(ram_block3a63),
	.ram_block3a31(ram_block3a31),
	.is_in_use_reg(is_in_use_reg),
	.address_reg_a_0(address_reg_a_0),
	.address_a({address_a[13],address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.ramaddr(ramaddr),
	.ramWEN(ramWEN),
	.always1(always1),
	.ir_loaded_address_reg_0(ir_loaded_address_reg_0),
	.ir_loaded_address_reg_1(ir_loaded_address_reg_1),
	.ir_loaded_address_reg_2(ir_loaded_address_reg_2),
	.ir_loaded_address_reg_3(ir_loaded_address_reg_3),
	.tdo(tdo),
	.data_a({data_a[31],data_a[30],data_a[29],data_a[28],data_a[27],data_a[26],data_a[25],data_a[24],data_a[23],data_a[22],data_a[21],data_a[20],data_a[19],data_a[18],data_a[17],data_a[16],data_a[15],data_a[14],data_a[13],data_a[12],data_a[11],data_a[10],data_a[9],data_a[8],data_a[7],data_a[6],data_a[5],data_a[4],data_a[3],data_a[2],data_a[1],data_a[0]}),
	.altera_internal_jtag(altera_internal_jtag),
	.state_4(state_4),
	.irf_reg_0_1(irf_reg_0_1),
	.irf_reg_1_1(irf_reg_1_1),
	.irf_reg_2_1(irf_reg_2_1),
	.irf_reg_3_1(irf_reg_3_1),
	.irf_reg_4_1(irf_reg_4_1),
	.node_ena_1(node_ena_1),
	.clr_reg(clr_reg),
	.virtual_ir_scan_reg(virtual_ir_scan_reg),
	.state_3(state_3),
	.state_5(state_5),
	.state_8(state_8),
	.altera_internal_jtag1(altera_internal_jtag1),
	.clock0(clock0),
	.devpor(devpor),
	.devclrn(devclrn),
	.devoe(devoe));

endmodule

module altsyncram_99f1 (
	ram_block3a32,
	ram_block3a0,
	ram_block3a33,
	ram_block3a1,
	ram_block3a34,
	ram_block3a2,
	ram_block3a35,
	ram_block3a3,
	ram_block3a36,
	ram_block3a4,
	ram_block3a37,
	ram_block3a5,
	ram_block3a38,
	ram_block3a6,
	ram_block3a39,
	ram_block3a7,
	ram_block3a40,
	ram_block3a8,
	ram_block3a41,
	ram_block3a9,
	ram_block3a42,
	ram_block3a10,
	ram_block3a43,
	ram_block3a11,
	ram_block3a44,
	ram_block3a12,
	ram_block3a45,
	ram_block3a13,
	ram_block3a46,
	ram_block3a14,
	ram_block3a47,
	ram_block3a15,
	ram_block3a48,
	ram_block3a16,
	ram_block3a49,
	ram_block3a17,
	ram_block3a50,
	ram_block3a18,
	ram_block3a51,
	ram_block3a19,
	ram_block3a52,
	ram_block3a20,
	ram_block3a53,
	ram_block3a21,
	ram_block3a54,
	ram_block3a22,
	ram_block3a55,
	ram_block3a23,
	ram_block3a56,
	ram_block3a24,
	ram_block3a57,
	ram_block3a25,
	ram_block3a58,
	ram_block3a26,
	ram_block3a59,
	ram_block3a27,
	ram_block3a60,
	ram_block3a28,
	ram_block3a61,
	ram_block3a29,
	ram_block3a62,
	ram_block3a30,
	ram_block3a63,
	ram_block3a31,
	is_in_use_reg,
	address_reg_a_0,
	address_a,
	ramaddr,
	ramWEN,
	always1,
	ir_loaded_address_reg_0,
	ir_loaded_address_reg_1,
	ir_loaded_address_reg_2,
	ir_loaded_address_reg_3,
	tdo,
	data_a,
	altera_internal_jtag,
	state_4,
	irf_reg_0_1,
	irf_reg_1_1,
	irf_reg_2_1,
	irf_reg_3_1,
	irf_reg_4_1,
	node_ena_1,
	clr_reg,
	virtual_ir_scan_reg,
	state_3,
	state_5,
	state_8,
	altera_internal_jtag1,
	clock0,
	devpor,
	devclrn,
	devoe);
output 	ram_block3a32;
output 	ram_block3a0;
output 	ram_block3a33;
output 	ram_block3a1;
output 	ram_block3a34;
output 	ram_block3a2;
output 	ram_block3a35;
output 	ram_block3a3;
output 	ram_block3a36;
output 	ram_block3a4;
output 	ram_block3a37;
output 	ram_block3a5;
output 	ram_block3a38;
output 	ram_block3a6;
output 	ram_block3a39;
output 	ram_block3a7;
output 	ram_block3a40;
output 	ram_block3a8;
output 	ram_block3a41;
output 	ram_block3a9;
output 	ram_block3a42;
output 	ram_block3a10;
output 	ram_block3a43;
output 	ram_block3a11;
output 	ram_block3a44;
output 	ram_block3a12;
output 	ram_block3a45;
output 	ram_block3a13;
output 	ram_block3a46;
output 	ram_block3a14;
output 	ram_block3a47;
output 	ram_block3a15;
output 	ram_block3a48;
output 	ram_block3a16;
output 	ram_block3a49;
output 	ram_block3a17;
output 	ram_block3a50;
output 	ram_block3a18;
output 	ram_block3a51;
output 	ram_block3a19;
output 	ram_block3a52;
output 	ram_block3a20;
output 	ram_block3a53;
output 	ram_block3a21;
output 	ram_block3a54;
output 	ram_block3a22;
output 	ram_block3a55;
output 	ram_block3a23;
output 	ram_block3a56;
output 	ram_block3a24;
output 	ram_block3a57;
output 	ram_block3a25;
output 	ram_block3a58;
output 	ram_block3a26;
output 	ram_block3a59;
output 	ram_block3a27;
output 	ram_block3a60;
output 	ram_block3a28;
output 	ram_block3a61;
output 	ram_block3a29;
output 	ram_block3a62;
output 	ram_block3a30;
output 	ram_block3a63;
output 	ram_block3a31;
output 	is_in_use_reg;
output 	address_reg_a_0;
input 	[13:0] address_a;
input 	ramaddr;
input 	ramWEN;
input 	always1;
output 	ir_loaded_address_reg_0;
output 	ir_loaded_address_reg_1;
output 	ir_loaded_address_reg_2;
output 	ir_loaded_address_reg_3;
output 	tdo;
input 	[31:0] data_a;
input 	altera_internal_jtag;
input 	state_4;
input 	irf_reg_0_1;
input 	irf_reg_1_1;
input 	irf_reg_2_1;
input 	irf_reg_3_1;
input 	irf_reg_4_1;
input 	node_ena_1;
input 	clr_reg;
input 	virtual_ir_scan_reg;
input 	state_3;
input 	state_5;
input 	state_8;
input 	altera_internal_jtag1;
input 	clock0;

// Design Ports Information

input 	devpor;
input 	devclrn;
input 	devoe;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
assign unknown = 1'bx;

wire \altsyncram1|ram_block3a32~PORTBDATAOUT0 ;
wire \altsyncram1|ram_block3a0~PORTBDATAOUT0 ;
wire \altsyncram1|ram_block3a33~PORTBDATAOUT0 ;
wire \altsyncram1|ram_block3a1~PORTBDATAOUT0 ;
wire \altsyncram1|ram_block3a34~PORTBDATAOUT0 ;
wire \altsyncram1|ram_block3a2~PORTBDATAOUT0 ;
wire \altsyncram1|ram_block3a35~PORTBDATAOUT0 ;
wire \altsyncram1|ram_block3a3~PORTBDATAOUT0 ;
wire \altsyncram1|ram_block3a36~PORTBDATAOUT0 ;
wire \altsyncram1|ram_block3a4~PORTBDATAOUT0 ;
wire \altsyncram1|ram_block3a37~PORTBDATAOUT0 ;
wire \altsyncram1|ram_block3a5~PORTBDATAOUT0 ;
wire \altsyncram1|ram_block3a38~PORTBDATAOUT0 ;
wire \altsyncram1|ram_block3a6~PORTBDATAOUT0 ;
wire \altsyncram1|ram_block3a39~PORTBDATAOUT0 ;
wire \altsyncram1|ram_block3a7~PORTBDATAOUT0 ;
wire \altsyncram1|ram_block3a40~PORTBDATAOUT0 ;
wire \altsyncram1|ram_block3a8~PORTBDATAOUT0 ;
wire \altsyncram1|ram_block3a41~PORTBDATAOUT0 ;
wire \altsyncram1|ram_block3a9~PORTBDATAOUT0 ;
wire \altsyncram1|ram_block3a42~PORTBDATAOUT0 ;
wire \altsyncram1|ram_block3a10~PORTBDATAOUT0 ;
wire \altsyncram1|ram_block3a43~PORTBDATAOUT0 ;
wire \altsyncram1|ram_block3a11~PORTBDATAOUT0 ;
wire \altsyncram1|ram_block3a44~PORTBDATAOUT0 ;
wire \altsyncram1|ram_block3a12~PORTBDATAOUT0 ;
wire \altsyncram1|ram_block3a45~PORTBDATAOUT0 ;
wire \altsyncram1|ram_block3a13~PORTBDATAOUT0 ;
wire \altsyncram1|ram_block3a46~PORTBDATAOUT0 ;
wire \altsyncram1|ram_block3a14~PORTBDATAOUT0 ;
wire \altsyncram1|ram_block3a47~PORTBDATAOUT0 ;
wire \altsyncram1|ram_block3a15~PORTBDATAOUT0 ;
wire \altsyncram1|ram_block3a48~PORTBDATAOUT0 ;
wire \altsyncram1|ram_block3a16~PORTBDATAOUT0 ;
wire \altsyncram1|ram_block3a49~PORTBDATAOUT0 ;
wire \altsyncram1|ram_block3a17~PORTBDATAOUT0 ;
wire \altsyncram1|ram_block3a50~PORTBDATAOUT0 ;
wire \altsyncram1|ram_block3a18~PORTBDATAOUT0 ;
wire \altsyncram1|ram_block3a51~PORTBDATAOUT0 ;
wire \altsyncram1|ram_block3a19~PORTBDATAOUT0 ;
wire \altsyncram1|ram_block3a52~PORTBDATAOUT0 ;
wire \altsyncram1|ram_block3a20~PORTBDATAOUT0 ;
wire \altsyncram1|ram_block3a53~PORTBDATAOUT0 ;
wire \altsyncram1|ram_block3a21~PORTBDATAOUT0 ;
wire \altsyncram1|ram_block3a54~PORTBDATAOUT0 ;
wire \altsyncram1|ram_block3a22~PORTBDATAOUT0 ;
wire \altsyncram1|ram_block3a55~PORTBDATAOUT0 ;
wire \altsyncram1|ram_block3a23~PORTBDATAOUT0 ;
wire \altsyncram1|ram_block3a56~PORTBDATAOUT0 ;
wire \altsyncram1|ram_block3a24~PORTBDATAOUT0 ;
wire \altsyncram1|ram_block3a57~PORTBDATAOUT0 ;
wire \altsyncram1|ram_block3a25~PORTBDATAOUT0 ;
wire \altsyncram1|ram_block3a58~PORTBDATAOUT0 ;
wire \altsyncram1|ram_block3a26~PORTBDATAOUT0 ;
wire \altsyncram1|ram_block3a59~PORTBDATAOUT0 ;
wire \altsyncram1|ram_block3a27~PORTBDATAOUT0 ;
wire \altsyncram1|ram_block3a60~PORTBDATAOUT0 ;
wire \altsyncram1|ram_block3a28~PORTBDATAOUT0 ;
wire \altsyncram1|ram_block3a61~PORTBDATAOUT0 ;
wire \altsyncram1|ram_block3a29~PORTBDATAOUT0 ;
wire \altsyncram1|ram_block3a62~PORTBDATAOUT0 ;
wire \altsyncram1|ram_block3a30~PORTBDATAOUT0 ;
wire \altsyncram1|ram_block3a63~PORTBDATAOUT0 ;
wire \altsyncram1|ram_block3a31~PORTBDATAOUT0 ;
wire \mgl_prim2|sdr~0_combout ;
wire [0:0] \altsyncram1|address_reg_b ;
wire [31:0] \mgl_prim2|ram_rom_data_reg ;
wire [13:0] \mgl_prim2|ram_rom_addr_reg ;


sld_mod_ram_rom mgl_prim2(
	.ram_block3a32(\altsyncram1|ram_block3a32~PORTBDATAOUT0 ),
	.ram_block3a0(\altsyncram1|ram_block3a0~PORTBDATAOUT0 ),
	.ram_block3a33(\altsyncram1|ram_block3a33~PORTBDATAOUT0 ),
	.ram_block3a1(\altsyncram1|ram_block3a1~PORTBDATAOUT0 ),
	.ram_block3a34(\altsyncram1|ram_block3a34~PORTBDATAOUT0 ),
	.ram_block3a2(\altsyncram1|ram_block3a2~PORTBDATAOUT0 ),
	.ram_block3a35(\altsyncram1|ram_block3a35~PORTBDATAOUT0 ),
	.ram_block3a3(\altsyncram1|ram_block3a3~PORTBDATAOUT0 ),
	.ram_block3a36(\altsyncram1|ram_block3a36~PORTBDATAOUT0 ),
	.ram_block3a4(\altsyncram1|ram_block3a4~PORTBDATAOUT0 ),
	.ram_block3a37(\altsyncram1|ram_block3a37~PORTBDATAOUT0 ),
	.ram_block3a5(\altsyncram1|ram_block3a5~PORTBDATAOUT0 ),
	.ram_block3a38(\altsyncram1|ram_block3a38~PORTBDATAOUT0 ),
	.ram_block3a6(\altsyncram1|ram_block3a6~PORTBDATAOUT0 ),
	.ram_block3a39(\altsyncram1|ram_block3a39~PORTBDATAOUT0 ),
	.ram_block3a7(\altsyncram1|ram_block3a7~PORTBDATAOUT0 ),
	.ram_block3a40(\altsyncram1|ram_block3a40~PORTBDATAOUT0 ),
	.ram_block3a8(\altsyncram1|ram_block3a8~PORTBDATAOUT0 ),
	.ram_block3a41(\altsyncram1|ram_block3a41~PORTBDATAOUT0 ),
	.ram_block3a9(\altsyncram1|ram_block3a9~PORTBDATAOUT0 ),
	.ram_block3a42(\altsyncram1|ram_block3a42~PORTBDATAOUT0 ),
	.ram_block3a10(\altsyncram1|ram_block3a10~PORTBDATAOUT0 ),
	.ram_block3a43(\altsyncram1|ram_block3a43~PORTBDATAOUT0 ),
	.ram_block3a11(\altsyncram1|ram_block3a11~PORTBDATAOUT0 ),
	.ram_block3a44(\altsyncram1|ram_block3a44~PORTBDATAOUT0 ),
	.ram_block3a12(\altsyncram1|ram_block3a12~PORTBDATAOUT0 ),
	.ram_block3a45(\altsyncram1|ram_block3a45~PORTBDATAOUT0 ),
	.ram_block3a13(\altsyncram1|ram_block3a13~PORTBDATAOUT0 ),
	.ram_block3a46(\altsyncram1|ram_block3a46~PORTBDATAOUT0 ),
	.ram_block3a14(\altsyncram1|ram_block3a14~PORTBDATAOUT0 ),
	.ram_block3a47(\altsyncram1|ram_block3a47~PORTBDATAOUT0 ),
	.ram_block3a15(\altsyncram1|ram_block3a15~PORTBDATAOUT0 ),
	.ram_block3a48(\altsyncram1|ram_block3a48~PORTBDATAOUT0 ),
	.ram_block3a16(\altsyncram1|ram_block3a16~PORTBDATAOUT0 ),
	.ram_block3a49(\altsyncram1|ram_block3a49~PORTBDATAOUT0 ),
	.ram_block3a17(\altsyncram1|ram_block3a17~PORTBDATAOUT0 ),
	.ram_block3a50(\altsyncram1|ram_block3a50~PORTBDATAOUT0 ),
	.ram_block3a18(\altsyncram1|ram_block3a18~PORTBDATAOUT0 ),
	.ram_block3a51(\altsyncram1|ram_block3a51~PORTBDATAOUT0 ),
	.ram_block3a19(\altsyncram1|ram_block3a19~PORTBDATAOUT0 ),
	.ram_block3a52(\altsyncram1|ram_block3a52~PORTBDATAOUT0 ),
	.ram_block3a20(\altsyncram1|ram_block3a20~PORTBDATAOUT0 ),
	.ram_block3a53(\altsyncram1|ram_block3a53~PORTBDATAOUT0 ),
	.ram_block3a21(\altsyncram1|ram_block3a21~PORTBDATAOUT0 ),
	.ram_block3a54(\altsyncram1|ram_block3a54~PORTBDATAOUT0 ),
	.ram_block3a22(\altsyncram1|ram_block3a22~PORTBDATAOUT0 ),
	.ram_block3a55(\altsyncram1|ram_block3a55~PORTBDATAOUT0 ),
	.ram_block3a23(\altsyncram1|ram_block3a23~PORTBDATAOUT0 ),
	.ram_block3a56(\altsyncram1|ram_block3a56~PORTBDATAOUT0 ),
	.ram_block3a24(\altsyncram1|ram_block3a24~PORTBDATAOUT0 ),
	.ram_block3a57(\altsyncram1|ram_block3a57~PORTBDATAOUT0 ),
	.ram_block3a25(\altsyncram1|ram_block3a25~PORTBDATAOUT0 ),
	.ram_block3a58(\altsyncram1|ram_block3a58~PORTBDATAOUT0 ),
	.ram_block3a26(\altsyncram1|ram_block3a26~PORTBDATAOUT0 ),
	.ram_block3a59(\altsyncram1|ram_block3a59~PORTBDATAOUT0 ),
	.ram_block3a27(\altsyncram1|ram_block3a27~PORTBDATAOUT0 ),
	.ram_block3a60(\altsyncram1|ram_block3a60~PORTBDATAOUT0 ),
	.ram_block3a28(\altsyncram1|ram_block3a28~PORTBDATAOUT0 ),
	.ram_block3a61(\altsyncram1|ram_block3a61~PORTBDATAOUT0 ),
	.ram_block3a29(\altsyncram1|ram_block3a29~PORTBDATAOUT0 ),
	.ram_block3a62(\altsyncram1|ram_block3a62~PORTBDATAOUT0 ),
	.ram_block3a30(\altsyncram1|ram_block3a30~PORTBDATAOUT0 ),
	.ram_block3a63(\altsyncram1|ram_block3a63~PORTBDATAOUT0 ),
	.ram_block3a31(\altsyncram1|ram_block3a31~PORTBDATAOUT0 ),
	.is_in_use_reg1(is_in_use_reg),
	.ram_rom_data_reg_0(\mgl_prim2|ram_rom_data_reg [0]),
	.ram_rom_addr_reg_13(\mgl_prim2|ram_rom_addr_reg [13]),
	.ram_rom_addr_reg_0(\mgl_prim2|ram_rom_addr_reg [0]),
	.ram_rom_addr_reg_1(\mgl_prim2|ram_rom_addr_reg [1]),
	.ram_rom_addr_reg_2(\mgl_prim2|ram_rom_addr_reg [2]),
	.ram_rom_addr_reg_3(\mgl_prim2|ram_rom_addr_reg [3]),
	.ram_rom_addr_reg_4(\mgl_prim2|ram_rom_addr_reg [4]),
	.ram_rom_addr_reg_5(\mgl_prim2|ram_rom_addr_reg [5]),
	.ram_rom_addr_reg_6(\mgl_prim2|ram_rom_addr_reg [6]),
	.ram_rom_addr_reg_7(\mgl_prim2|ram_rom_addr_reg [7]),
	.ram_rom_addr_reg_8(\mgl_prim2|ram_rom_addr_reg [8]),
	.ram_rom_addr_reg_9(\mgl_prim2|ram_rom_addr_reg [9]),
	.ram_rom_addr_reg_10(\mgl_prim2|ram_rom_addr_reg [10]),
	.ram_rom_addr_reg_11(\mgl_prim2|ram_rom_addr_reg [11]),
	.ram_rom_addr_reg_12(\mgl_prim2|ram_rom_addr_reg [12]),
	.ram_rom_data_reg_1(\mgl_prim2|ram_rom_data_reg [1]),
	.ram_rom_data_reg_2(\mgl_prim2|ram_rom_data_reg [2]),
	.ram_rom_data_reg_3(\mgl_prim2|ram_rom_data_reg [3]),
	.ram_rom_data_reg_4(\mgl_prim2|ram_rom_data_reg [4]),
	.ram_rom_data_reg_5(\mgl_prim2|ram_rom_data_reg [5]),
	.ram_rom_data_reg_6(\mgl_prim2|ram_rom_data_reg [6]),
	.ram_rom_data_reg_7(\mgl_prim2|ram_rom_data_reg [7]),
	.ram_rom_data_reg_8(\mgl_prim2|ram_rom_data_reg [8]),
	.ram_rom_data_reg_9(\mgl_prim2|ram_rom_data_reg [9]),
	.ram_rom_data_reg_10(\mgl_prim2|ram_rom_data_reg [10]),
	.ram_rom_data_reg_11(\mgl_prim2|ram_rom_data_reg [11]),
	.ram_rom_data_reg_12(\mgl_prim2|ram_rom_data_reg [12]),
	.ram_rom_data_reg_13(\mgl_prim2|ram_rom_data_reg [13]),
	.ram_rom_data_reg_14(\mgl_prim2|ram_rom_data_reg [14]),
	.ram_rom_data_reg_15(\mgl_prim2|ram_rom_data_reg [15]),
	.ram_rom_data_reg_16(\mgl_prim2|ram_rom_data_reg [16]),
	.ram_rom_data_reg_17(\mgl_prim2|ram_rom_data_reg [17]),
	.ram_rom_data_reg_18(\mgl_prim2|ram_rom_data_reg [18]),
	.ram_rom_data_reg_19(\mgl_prim2|ram_rom_data_reg [19]),
	.ram_rom_data_reg_20(\mgl_prim2|ram_rom_data_reg [20]),
	.ram_rom_data_reg_21(\mgl_prim2|ram_rom_data_reg [21]),
	.ram_rom_data_reg_22(\mgl_prim2|ram_rom_data_reg [22]),
	.ram_rom_data_reg_23(\mgl_prim2|ram_rom_data_reg [23]),
	.ram_rom_data_reg_24(\mgl_prim2|ram_rom_data_reg [24]),
	.ram_rom_data_reg_25(\mgl_prim2|ram_rom_data_reg [25]),
	.ram_rom_data_reg_26(\mgl_prim2|ram_rom_data_reg [26]),
	.ram_rom_data_reg_27(\mgl_prim2|ram_rom_data_reg [27]),
	.ram_rom_data_reg_28(\mgl_prim2|ram_rom_data_reg [28]),
	.ram_rom_data_reg_29(\mgl_prim2|ram_rom_data_reg [29]),
	.ram_rom_data_reg_30(\mgl_prim2|ram_rom_data_reg [30]),
	.ram_rom_data_reg_31(\mgl_prim2|ram_rom_data_reg [31]),
	.ir_loaded_address_reg_0(ir_loaded_address_reg_0),
	.ir_loaded_address_reg_1(ir_loaded_address_reg_1),
	.ir_loaded_address_reg_2(ir_loaded_address_reg_2),
	.ir_loaded_address_reg_3(ir_loaded_address_reg_3),
	.tdo(tdo),
	.sdr(\mgl_prim2|sdr~0_combout ),
	.address_reg_b_0(\altsyncram1|address_reg_b [0]),
	.altera_internal_jtag(altera_internal_jtag),
	.state_4(state_4),
	.ir_in({gnd,irf_reg_3_1,gnd,gnd,irf_reg_0_1}),
	.irf_reg_1_1(irf_reg_1_1),
	.irf_reg_2_1(irf_reg_2_1),
	.irf_reg_4_1(irf_reg_4_1),
	.node_ena_1(node_ena_1),
	.clr(clr_reg),
	.virtual_ir_scan_reg(virtual_ir_scan_reg),
	.state_3(state_3),
	.state_5(state_5),
	.state_8(state_8),
	.raw_tck(altera_internal_jtag1),
	.devpor(devpor),
	.devclrn(devclrn),
	.devoe(devoe));

altsyncram_fta2 altsyncram1(
	.ram_block3a321(ram_block3a32),
	.ram_block3a322(\altsyncram1|ram_block3a32~PORTBDATAOUT0 ),
	.ram_block3a01(ram_block3a0),
	.ram_block3a02(\altsyncram1|ram_block3a0~PORTBDATAOUT0 ),
	.ram_block3a331(ram_block3a33),
	.ram_block3a332(\altsyncram1|ram_block3a33~PORTBDATAOUT0 ),
	.ram_block3a110(ram_block3a1),
	.ram_block3a111(\altsyncram1|ram_block3a1~PORTBDATAOUT0 ),
	.ram_block3a341(ram_block3a34),
	.ram_block3a342(\altsyncram1|ram_block3a34~PORTBDATAOUT0 ),
	.ram_block3a210(ram_block3a2),
	.ram_block3a211(\altsyncram1|ram_block3a2~PORTBDATAOUT0 ),
	.ram_block3a351(ram_block3a35),
	.ram_block3a352(\altsyncram1|ram_block3a35~PORTBDATAOUT0 ),
	.ram_block3a310(ram_block3a3),
	.ram_block3a311(\altsyncram1|ram_block3a3~PORTBDATAOUT0 ),
	.ram_block3a361(ram_block3a36),
	.ram_block3a362(\altsyncram1|ram_block3a36~PORTBDATAOUT0 ),
	.ram_block3a410(ram_block3a4),
	.ram_block3a411(\altsyncram1|ram_block3a4~PORTBDATAOUT0 ),
	.ram_block3a371(ram_block3a37),
	.ram_block3a372(\altsyncram1|ram_block3a37~PORTBDATAOUT0 ),
	.ram_block3a510(ram_block3a5),
	.ram_block3a511(\altsyncram1|ram_block3a5~PORTBDATAOUT0 ),
	.ram_block3a381(ram_block3a38),
	.ram_block3a382(\altsyncram1|ram_block3a38~PORTBDATAOUT0 ),
	.ram_block3a64(ram_block3a6),
	.ram_block3a65(\altsyncram1|ram_block3a6~PORTBDATAOUT0 ),
	.ram_block3a391(ram_block3a39),
	.ram_block3a392(\altsyncram1|ram_block3a39~PORTBDATAOUT0 ),
	.ram_block3a71(ram_block3a7),
	.ram_block3a72(\altsyncram1|ram_block3a7~PORTBDATAOUT0 ),
	.ram_block3a401(ram_block3a40),
	.ram_block3a402(\altsyncram1|ram_block3a40~PORTBDATAOUT0 ),
	.ram_block3a81(ram_block3a8),
	.ram_block3a82(\altsyncram1|ram_block3a8~PORTBDATAOUT0 ),
	.ram_block3a412(ram_block3a41),
	.ram_block3a413(\altsyncram1|ram_block3a41~PORTBDATAOUT0 ),
	.ram_block3a91(ram_block3a9),
	.ram_block3a92(\altsyncram1|ram_block3a9~PORTBDATAOUT0 ),
	.ram_block3a421(ram_block3a42),
	.ram_block3a422(\altsyncram1|ram_block3a42~PORTBDATAOUT0 ),
	.ram_block3a101(ram_block3a10),
	.ram_block3a102(\altsyncram1|ram_block3a10~PORTBDATAOUT0 ),
	.ram_block3a431(ram_block3a43),
	.ram_block3a432(\altsyncram1|ram_block3a43~PORTBDATAOUT0 ),
	.ram_block3a112(ram_block3a11),
	.ram_block3a113(\altsyncram1|ram_block3a11~PORTBDATAOUT0 ),
	.ram_block3a441(ram_block3a44),
	.ram_block3a442(\altsyncram1|ram_block3a44~PORTBDATAOUT0 ),
	.ram_block3a121(ram_block3a12),
	.ram_block3a122(\altsyncram1|ram_block3a12~PORTBDATAOUT0 ),
	.ram_block3a451(ram_block3a45),
	.ram_block3a452(\altsyncram1|ram_block3a45~PORTBDATAOUT0 ),
	.ram_block3a131(ram_block3a13),
	.ram_block3a132(\altsyncram1|ram_block3a13~PORTBDATAOUT0 ),
	.ram_block3a461(ram_block3a46),
	.ram_block3a462(\altsyncram1|ram_block3a46~PORTBDATAOUT0 ),
	.ram_block3a141(ram_block3a14),
	.ram_block3a142(\altsyncram1|ram_block3a14~PORTBDATAOUT0 ),
	.ram_block3a471(ram_block3a47),
	.ram_block3a472(\altsyncram1|ram_block3a47~PORTBDATAOUT0 ),
	.ram_block3a151(ram_block3a15),
	.ram_block3a152(\altsyncram1|ram_block3a15~PORTBDATAOUT0 ),
	.ram_block3a481(ram_block3a48),
	.ram_block3a482(\altsyncram1|ram_block3a48~PORTBDATAOUT0 ),
	.ram_block3a161(ram_block3a16),
	.ram_block3a162(\altsyncram1|ram_block3a16~PORTBDATAOUT0 ),
	.ram_block3a491(ram_block3a49),
	.ram_block3a492(\altsyncram1|ram_block3a49~PORTBDATAOUT0 ),
	.ram_block3a171(ram_block3a17),
	.ram_block3a172(\altsyncram1|ram_block3a17~PORTBDATAOUT0 ),
	.ram_block3a501(ram_block3a50),
	.ram_block3a502(\altsyncram1|ram_block3a50~PORTBDATAOUT0 ),
	.ram_block3a181(ram_block3a18),
	.ram_block3a182(\altsyncram1|ram_block3a18~PORTBDATAOUT0 ),
	.ram_block3a512(ram_block3a51),
	.ram_block3a513(\altsyncram1|ram_block3a51~PORTBDATAOUT0 ),
	.ram_block3a191(ram_block3a19),
	.ram_block3a192(\altsyncram1|ram_block3a19~PORTBDATAOUT0 ),
	.ram_block3a521(ram_block3a52),
	.ram_block3a522(\altsyncram1|ram_block3a52~PORTBDATAOUT0 ),
	.ram_block3a201(ram_block3a20),
	.ram_block3a202(\altsyncram1|ram_block3a20~PORTBDATAOUT0 ),
	.ram_block3a531(ram_block3a53),
	.ram_block3a532(\altsyncram1|ram_block3a53~PORTBDATAOUT0 ),
	.ram_block3a212(ram_block3a21),
	.ram_block3a213(\altsyncram1|ram_block3a21~PORTBDATAOUT0 ),
	.ram_block3a541(ram_block3a54),
	.ram_block3a542(\altsyncram1|ram_block3a54~PORTBDATAOUT0 ),
	.ram_block3a221(ram_block3a22),
	.ram_block3a222(\altsyncram1|ram_block3a22~PORTBDATAOUT0 ),
	.ram_block3a551(ram_block3a55),
	.ram_block3a552(\altsyncram1|ram_block3a55~PORTBDATAOUT0 ),
	.ram_block3a231(ram_block3a23),
	.ram_block3a232(\altsyncram1|ram_block3a23~PORTBDATAOUT0 ),
	.ram_block3a561(ram_block3a56),
	.ram_block3a562(\altsyncram1|ram_block3a56~PORTBDATAOUT0 ),
	.ram_block3a241(ram_block3a24),
	.ram_block3a242(\altsyncram1|ram_block3a24~PORTBDATAOUT0 ),
	.ram_block3a571(ram_block3a57),
	.ram_block3a572(\altsyncram1|ram_block3a57~PORTBDATAOUT0 ),
	.ram_block3a251(ram_block3a25),
	.ram_block3a252(\altsyncram1|ram_block3a25~PORTBDATAOUT0 ),
	.ram_block3a581(ram_block3a58),
	.ram_block3a582(\altsyncram1|ram_block3a58~PORTBDATAOUT0 ),
	.ram_block3a261(ram_block3a26),
	.ram_block3a262(\altsyncram1|ram_block3a26~PORTBDATAOUT0 ),
	.ram_block3a591(ram_block3a59),
	.ram_block3a592(\altsyncram1|ram_block3a59~PORTBDATAOUT0 ),
	.ram_block3a271(ram_block3a27),
	.ram_block3a272(\altsyncram1|ram_block3a27~PORTBDATAOUT0 ),
	.ram_block3a601(ram_block3a60),
	.ram_block3a602(\altsyncram1|ram_block3a60~PORTBDATAOUT0 ),
	.ram_block3a281(ram_block3a28),
	.ram_block3a282(\altsyncram1|ram_block3a28~PORTBDATAOUT0 ),
	.ram_block3a611(ram_block3a61),
	.ram_block3a612(\altsyncram1|ram_block3a61~PORTBDATAOUT0 ),
	.ram_block3a291(ram_block3a29),
	.ram_block3a292(\altsyncram1|ram_block3a29~PORTBDATAOUT0 ),
	.ram_block3a621(ram_block3a62),
	.ram_block3a622(\altsyncram1|ram_block3a62~PORTBDATAOUT0 ),
	.ram_block3a301(ram_block3a30),
	.ram_block3a302(\altsyncram1|ram_block3a30~PORTBDATAOUT0 ),
	.ram_block3a631(ram_block3a63),
	.ram_block3a632(\altsyncram1|ram_block3a63~PORTBDATAOUT0 ),
	.ram_block3a312(ram_block3a31),
	.ram_block3a313(\altsyncram1|ram_block3a31~PORTBDATAOUT0 ),
	.data_b({\mgl_prim2|ram_rom_data_reg [31],\mgl_prim2|ram_rom_data_reg [30],\mgl_prim2|ram_rom_data_reg [29],\mgl_prim2|ram_rom_data_reg [28],\mgl_prim2|ram_rom_data_reg [27],\mgl_prim2|ram_rom_data_reg [26],\mgl_prim2|ram_rom_data_reg [25],\mgl_prim2|ram_rom_data_reg [24],\mgl_prim2|ram_rom_data_reg [23],
\mgl_prim2|ram_rom_data_reg [22],\mgl_prim2|ram_rom_data_reg [21],\mgl_prim2|ram_rom_data_reg [20],\mgl_prim2|ram_rom_data_reg [19],\mgl_prim2|ram_rom_data_reg [18],\mgl_prim2|ram_rom_data_reg [17],\mgl_prim2|ram_rom_data_reg [16],\mgl_prim2|ram_rom_data_reg [15],\mgl_prim2|ram_rom_data_reg [14],
\mgl_prim2|ram_rom_data_reg [13],\mgl_prim2|ram_rom_data_reg [12],\mgl_prim2|ram_rom_data_reg [11],\mgl_prim2|ram_rom_data_reg [10],\mgl_prim2|ram_rom_data_reg [9],\mgl_prim2|ram_rom_data_reg [8],\mgl_prim2|ram_rom_data_reg [7],\mgl_prim2|ram_rom_data_reg [6],\mgl_prim2|ram_rom_data_reg [5],
\mgl_prim2|ram_rom_data_reg [4],\mgl_prim2|ram_rom_data_reg [3],\mgl_prim2|ram_rom_data_reg [2],\mgl_prim2|ram_rom_data_reg [1],\mgl_prim2|ram_rom_data_reg [0]}),
	.ram_rom_addr_reg_13(\mgl_prim2|ram_rom_addr_reg [13]),
	.address_b({gnd,\mgl_prim2|ram_rom_addr_reg [12],\mgl_prim2|ram_rom_addr_reg [11],\mgl_prim2|ram_rom_addr_reg [10],\mgl_prim2|ram_rom_addr_reg [9],\mgl_prim2|ram_rom_addr_reg [8],\mgl_prim2|ram_rom_addr_reg [7],\mgl_prim2|ram_rom_addr_reg [6],\mgl_prim2|ram_rom_addr_reg [5],\mgl_prim2|ram_rom_addr_reg [4],
\mgl_prim2|ram_rom_addr_reg [3],\mgl_prim2|ram_rom_addr_reg [2],\mgl_prim2|ram_rom_addr_reg [1],\mgl_prim2|ram_rom_addr_reg [0]}),
	.address_reg_a_0(address_reg_a_0),
	.address_a({address_a[13],address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.ramaddr(ramaddr),
	.ramWEN(ramWEN),
	.always1(always1),
	.sdr(\mgl_prim2|sdr~0_combout ),
	.data_a({data_a[31],data_a[30],data_a[29],data_a[28],data_a[27],data_a[26],data_a[25],data_a[24],data_a[23],data_a[22],data_a[21],data_a[20],data_a[19],data_a[18],data_a[17],data_a[16],data_a[15],data_a[14],data_a[13],data_a[12],data_a[11],data_a[10],data_a[9],data_a[8],data_a[7],data_a[6],data_a[5],data_a[4],data_a[3],data_a[2],data_a[1],data_a[0]}),
	.address_reg_b_0(\altsyncram1|address_reg_b [0]),
	.irf_reg_2_1(irf_reg_2_1),
	.state_5(state_5),
	.clock1(altera_internal_jtag1),
	.clock0(clock0),
	.devpor(devpor),
	.devclrn(devclrn),
	.devoe(devoe));

endmodule

module altsyncram_fta2 (
	ram_block3a321,
	ram_block3a322,
	ram_block3a01,
	ram_block3a02,
	ram_block3a331,
	ram_block3a332,
	ram_block3a110,
	ram_block3a111,
	ram_block3a341,
	ram_block3a342,
	ram_block3a210,
	ram_block3a211,
	ram_block3a351,
	ram_block3a352,
	ram_block3a310,
	ram_block3a311,
	ram_block3a361,
	ram_block3a362,
	ram_block3a410,
	ram_block3a411,
	ram_block3a371,
	ram_block3a372,
	ram_block3a510,
	ram_block3a511,
	ram_block3a381,
	ram_block3a382,
	ram_block3a64,
	ram_block3a65,
	ram_block3a391,
	ram_block3a392,
	ram_block3a71,
	ram_block3a72,
	ram_block3a401,
	ram_block3a402,
	ram_block3a81,
	ram_block3a82,
	ram_block3a412,
	ram_block3a413,
	ram_block3a91,
	ram_block3a92,
	ram_block3a421,
	ram_block3a422,
	ram_block3a101,
	ram_block3a102,
	ram_block3a431,
	ram_block3a432,
	ram_block3a112,
	ram_block3a113,
	ram_block3a441,
	ram_block3a442,
	ram_block3a121,
	ram_block3a122,
	ram_block3a451,
	ram_block3a452,
	ram_block3a131,
	ram_block3a132,
	ram_block3a461,
	ram_block3a462,
	ram_block3a141,
	ram_block3a142,
	ram_block3a471,
	ram_block3a472,
	ram_block3a151,
	ram_block3a152,
	ram_block3a481,
	ram_block3a482,
	ram_block3a161,
	ram_block3a162,
	ram_block3a491,
	ram_block3a492,
	ram_block3a171,
	ram_block3a172,
	ram_block3a501,
	ram_block3a502,
	ram_block3a181,
	ram_block3a182,
	ram_block3a512,
	ram_block3a513,
	ram_block3a191,
	ram_block3a192,
	ram_block3a521,
	ram_block3a522,
	ram_block3a201,
	ram_block3a202,
	ram_block3a531,
	ram_block3a532,
	ram_block3a212,
	ram_block3a213,
	ram_block3a541,
	ram_block3a542,
	ram_block3a221,
	ram_block3a222,
	ram_block3a551,
	ram_block3a552,
	ram_block3a231,
	ram_block3a232,
	ram_block3a561,
	ram_block3a562,
	ram_block3a241,
	ram_block3a242,
	ram_block3a571,
	ram_block3a572,
	ram_block3a251,
	ram_block3a252,
	ram_block3a581,
	ram_block3a582,
	ram_block3a261,
	ram_block3a262,
	ram_block3a591,
	ram_block3a592,
	ram_block3a271,
	ram_block3a272,
	ram_block3a601,
	ram_block3a602,
	ram_block3a281,
	ram_block3a282,
	ram_block3a611,
	ram_block3a612,
	ram_block3a291,
	ram_block3a292,
	ram_block3a621,
	ram_block3a622,
	ram_block3a301,
	ram_block3a302,
	ram_block3a631,
	ram_block3a632,
	ram_block3a312,
	ram_block3a313,
	data_b,
	ram_rom_addr_reg_13,
	address_b,
	address_reg_a_0,
	address_a,
	ramaddr,
	ramWEN,
	always1,
	sdr,
	data_a,
	address_reg_b_0,
	irf_reg_2_1,
	state_5,
	clock1,
	clock0,
	devpor,
	devclrn,
	devoe);
output 	ram_block3a321;
output 	ram_block3a322;
output 	ram_block3a01;
output 	ram_block3a02;
output 	ram_block3a331;
output 	ram_block3a332;
output 	ram_block3a110;
output 	ram_block3a111;
output 	ram_block3a341;
output 	ram_block3a342;
output 	ram_block3a210;
output 	ram_block3a211;
output 	ram_block3a351;
output 	ram_block3a352;
output 	ram_block3a310;
output 	ram_block3a311;
output 	ram_block3a361;
output 	ram_block3a362;
output 	ram_block3a410;
output 	ram_block3a411;
output 	ram_block3a371;
output 	ram_block3a372;
output 	ram_block3a510;
output 	ram_block3a511;
output 	ram_block3a381;
output 	ram_block3a382;
output 	ram_block3a64;
output 	ram_block3a65;
output 	ram_block3a391;
output 	ram_block3a392;
output 	ram_block3a71;
output 	ram_block3a72;
output 	ram_block3a401;
output 	ram_block3a402;
output 	ram_block3a81;
output 	ram_block3a82;
output 	ram_block3a412;
output 	ram_block3a413;
output 	ram_block3a91;
output 	ram_block3a92;
output 	ram_block3a421;
output 	ram_block3a422;
output 	ram_block3a101;
output 	ram_block3a102;
output 	ram_block3a431;
output 	ram_block3a432;
output 	ram_block3a112;
output 	ram_block3a113;
output 	ram_block3a441;
output 	ram_block3a442;
output 	ram_block3a121;
output 	ram_block3a122;
output 	ram_block3a451;
output 	ram_block3a452;
output 	ram_block3a131;
output 	ram_block3a132;
output 	ram_block3a461;
output 	ram_block3a462;
output 	ram_block3a141;
output 	ram_block3a142;
output 	ram_block3a471;
output 	ram_block3a472;
output 	ram_block3a151;
output 	ram_block3a152;
output 	ram_block3a481;
output 	ram_block3a482;
output 	ram_block3a161;
output 	ram_block3a162;
output 	ram_block3a491;
output 	ram_block3a492;
output 	ram_block3a171;
output 	ram_block3a172;
output 	ram_block3a501;
output 	ram_block3a502;
output 	ram_block3a181;
output 	ram_block3a182;
output 	ram_block3a512;
output 	ram_block3a513;
output 	ram_block3a191;
output 	ram_block3a192;
output 	ram_block3a521;
output 	ram_block3a522;
output 	ram_block3a201;
output 	ram_block3a202;
output 	ram_block3a531;
output 	ram_block3a532;
output 	ram_block3a212;
output 	ram_block3a213;
output 	ram_block3a541;
output 	ram_block3a542;
output 	ram_block3a221;
output 	ram_block3a222;
output 	ram_block3a551;
output 	ram_block3a552;
output 	ram_block3a231;
output 	ram_block3a232;
output 	ram_block3a561;
output 	ram_block3a562;
output 	ram_block3a241;
output 	ram_block3a242;
output 	ram_block3a571;
output 	ram_block3a572;
output 	ram_block3a251;
output 	ram_block3a252;
output 	ram_block3a581;
output 	ram_block3a582;
output 	ram_block3a261;
output 	ram_block3a262;
output 	ram_block3a591;
output 	ram_block3a592;
output 	ram_block3a271;
output 	ram_block3a272;
output 	ram_block3a601;
output 	ram_block3a602;
output 	ram_block3a281;
output 	ram_block3a282;
output 	ram_block3a611;
output 	ram_block3a612;
output 	ram_block3a291;
output 	ram_block3a292;
output 	ram_block3a621;
output 	ram_block3a622;
output 	ram_block3a301;
output 	ram_block3a302;
output 	ram_block3a631;
output 	ram_block3a632;
output 	ram_block3a312;
output 	ram_block3a313;
input 	[31:0] data_b;
input 	ram_rom_addr_reg_13;
input 	[13:0] address_b;
output 	address_reg_a_0;
input 	[13:0] address_a;
input 	ramaddr;
input 	ramWEN;
input 	always1;
input 	sdr;
input 	[31:0] data_a;
output 	address_reg_b_0;
input 	irf_reg_2_1;
input 	state_5;
input 	clock1;
input 	clock0;

// Design Ports Information

input 	devpor;
input 	devclrn;
input 	devoe;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
assign unknown = 1'bx;

wire \decode4|eq_node[1]~0_combout ;
wire \decode5|eq_node[1]~0_combout ;
wire \decode4|eq_node[0]~1_combout ;
wire \decode5|eq_node[0]~1_combout ;
wire \address_reg_b[0]~feeder_combout ;

wire [0:0] ram_block3a32_PORTADATAOUT_bus;
wire [0:0] ram_block3a32_PORTBDATAOUT_bus;
wire [0:0] ram_block3a0_PORTADATAOUT_bus;
wire [0:0] ram_block3a0_PORTBDATAOUT_bus;
wire [0:0] ram_block3a33_PORTADATAOUT_bus;
wire [0:0] ram_block3a33_PORTBDATAOUT_bus;
wire [0:0] ram_block3a1_PORTADATAOUT_bus;
wire [0:0] ram_block3a1_PORTBDATAOUT_bus;
wire [0:0] ram_block3a34_PORTADATAOUT_bus;
wire [0:0] ram_block3a34_PORTBDATAOUT_bus;
wire [0:0] ram_block3a2_PORTADATAOUT_bus;
wire [0:0] ram_block3a2_PORTBDATAOUT_bus;
wire [0:0] ram_block3a35_PORTADATAOUT_bus;
wire [0:0] ram_block3a35_PORTBDATAOUT_bus;
wire [0:0] ram_block3a3_PORTADATAOUT_bus;
wire [0:0] ram_block3a3_PORTBDATAOUT_bus;
wire [0:0] ram_block3a36_PORTADATAOUT_bus;
wire [0:0] ram_block3a36_PORTBDATAOUT_bus;
wire [0:0] ram_block3a4_PORTADATAOUT_bus;
wire [0:0] ram_block3a4_PORTBDATAOUT_bus;
wire [0:0] ram_block3a37_PORTADATAOUT_bus;
wire [0:0] ram_block3a37_PORTBDATAOUT_bus;
wire [0:0] ram_block3a5_PORTADATAOUT_bus;
wire [0:0] ram_block3a5_PORTBDATAOUT_bus;
wire [0:0] ram_block3a38_PORTADATAOUT_bus;
wire [0:0] ram_block3a38_PORTBDATAOUT_bus;
wire [0:0] ram_block3a6_PORTADATAOUT_bus;
wire [0:0] ram_block3a6_PORTBDATAOUT_bus;
wire [0:0] ram_block3a39_PORTADATAOUT_bus;
wire [0:0] ram_block3a39_PORTBDATAOUT_bus;
wire [0:0] ram_block3a7_PORTADATAOUT_bus;
wire [0:0] ram_block3a7_PORTBDATAOUT_bus;
wire [0:0] ram_block3a40_PORTADATAOUT_bus;
wire [0:0] ram_block3a40_PORTBDATAOUT_bus;
wire [0:0] ram_block3a8_PORTADATAOUT_bus;
wire [0:0] ram_block3a8_PORTBDATAOUT_bus;
wire [0:0] ram_block3a41_PORTADATAOUT_bus;
wire [0:0] ram_block3a41_PORTBDATAOUT_bus;
wire [0:0] ram_block3a9_PORTADATAOUT_bus;
wire [0:0] ram_block3a9_PORTBDATAOUT_bus;
wire [0:0] ram_block3a42_PORTADATAOUT_bus;
wire [0:0] ram_block3a42_PORTBDATAOUT_bus;
wire [0:0] ram_block3a10_PORTADATAOUT_bus;
wire [0:0] ram_block3a10_PORTBDATAOUT_bus;
wire [0:0] ram_block3a43_PORTADATAOUT_bus;
wire [0:0] ram_block3a43_PORTBDATAOUT_bus;
wire [0:0] ram_block3a11_PORTADATAOUT_bus;
wire [0:0] ram_block3a11_PORTBDATAOUT_bus;
wire [0:0] ram_block3a44_PORTADATAOUT_bus;
wire [0:0] ram_block3a44_PORTBDATAOUT_bus;
wire [0:0] ram_block3a12_PORTADATAOUT_bus;
wire [0:0] ram_block3a12_PORTBDATAOUT_bus;
wire [0:0] ram_block3a45_PORTADATAOUT_bus;
wire [0:0] ram_block3a45_PORTBDATAOUT_bus;
wire [0:0] ram_block3a13_PORTADATAOUT_bus;
wire [0:0] ram_block3a13_PORTBDATAOUT_bus;
wire [0:0] ram_block3a46_PORTADATAOUT_bus;
wire [0:0] ram_block3a46_PORTBDATAOUT_bus;
wire [0:0] ram_block3a14_PORTADATAOUT_bus;
wire [0:0] ram_block3a14_PORTBDATAOUT_bus;
wire [0:0] ram_block3a47_PORTADATAOUT_bus;
wire [0:0] ram_block3a47_PORTBDATAOUT_bus;
wire [0:0] ram_block3a15_PORTADATAOUT_bus;
wire [0:0] ram_block3a15_PORTBDATAOUT_bus;
wire [0:0] ram_block3a48_PORTADATAOUT_bus;
wire [0:0] ram_block3a48_PORTBDATAOUT_bus;
wire [0:0] ram_block3a16_PORTADATAOUT_bus;
wire [0:0] ram_block3a16_PORTBDATAOUT_bus;
wire [0:0] ram_block3a49_PORTADATAOUT_bus;
wire [0:0] ram_block3a49_PORTBDATAOUT_bus;
wire [0:0] ram_block3a17_PORTADATAOUT_bus;
wire [0:0] ram_block3a17_PORTBDATAOUT_bus;
wire [0:0] ram_block3a50_PORTADATAOUT_bus;
wire [0:0] ram_block3a50_PORTBDATAOUT_bus;
wire [0:0] ram_block3a18_PORTADATAOUT_bus;
wire [0:0] ram_block3a18_PORTBDATAOUT_bus;
wire [0:0] ram_block3a51_PORTADATAOUT_bus;
wire [0:0] ram_block3a51_PORTBDATAOUT_bus;
wire [0:0] ram_block3a19_PORTADATAOUT_bus;
wire [0:0] ram_block3a19_PORTBDATAOUT_bus;
wire [0:0] ram_block3a52_PORTADATAOUT_bus;
wire [0:0] ram_block3a52_PORTBDATAOUT_bus;
wire [0:0] ram_block3a20_PORTADATAOUT_bus;
wire [0:0] ram_block3a20_PORTBDATAOUT_bus;
wire [0:0] ram_block3a53_PORTADATAOUT_bus;
wire [0:0] ram_block3a53_PORTBDATAOUT_bus;
wire [0:0] ram_block3a21_PORTADATAOUT_bus;
wire [0:0] ram_block3a21_PORTBDATAOUT_bus;
wire [0:0] ram_block3a54_PORTADATAOUT_bus;
wire [0:0] ram_block3a54_PORTBDATAOUT_bus;
wire [0:0] ram_block3a22_PORTADATAOUT_bus;
wire [0:0] ram_block3a22_PORTBDATAOUT_bus;
wire [0:0] ram_block3a55_PORTADATAOUT_bus;
wire [0:0] ram_block3a55_PORTBDATAOUT_bus;
wire [0:0] ram_block3a23_PORTADATAOUT_bus;
wire [0:0] ram_block3a23_PORTBDATAOUT_bus;
wire [0:0] ram_block3a56_PORTADATAOUT_bus;
wire [0:0] ram_block3a56_PORTBDATAOUT_bus;
wire [0:0] ram_block3a24_PORTADATAOUT_bus;
wire [0:0] ram_block3a24_PORTBDATAOUT_bus;
wire [0:0] ram_block3a57_PORTADATAOUT_bus;
wire [0:0] ram_block3a57_PORTBDATAOUT_bus;
wire [0:0] ram_block3a25_PORTADATAOUT_bus;
wire [0:0] ram_block3a25_PORTBDATAOUT_bus;
wire [0:0] ram_block3a58_PORTADATAOUT_bus;
wire [0:0] ram_block3a58_PORTBDATAOUT_bus;
wire [0:0] ram_block3a26_PORTADATAOUT_bus;
wire [0:0] ram_block3a26_PORTBDATAOUT_bus;
wire [0:0] ram_block3a59_PORTADATAOUT_bus;
wire [0:0] ram_block3a59_PORTBDATAOUT_bus;
wire [0:0] ram_block3a27_PORTADATAOUT_bus;
wire [0:0] ram_block3a27_PORTBDATAOUT_bus;
wire [0:0] ram_block3a60_PORTADATAOUT_bus;
wire [0:0] ram_block3a60_PORTBDATAOUT_bus;
wire [0:0] ram_block3a28_PORTADATAOUT_bus;
wire [0:0] ram_block3a28_PORTBDATAOUT_bus;
wire [0:0] ram_block3a61_PORTADATAOUT_bus;
wire [0:0] ram_block3a61_PORTBDATAOUT_bus;
wire [0:0] ram_block3a29_PORTADATAOUT_bus;
wire [0:0] ram_block3a29_PORTBDATAOUT_bus;
wire [0:0] ram_block3a62_PORTADATAOUT_bus;
wire [0:0] ram_block3a62_PORTBDATAOUT_bus;
wire [0:0] ram_block3a30_PORTADATAOUT_bus;
wire [0:0] ram_block3a30_PORTBDATAOUT_bus;
wire [0:0] ram_block3a63_PORTADATAOUT_bus;
wire [0:0] ram_block3a63_PORTBDATAOUT_bus;
wire [0:0] ram_block3a31_PORTADATAOUT_bus;
wire [0:0] ram_block3a31_PORTBDATAOUT_bus;

assign ram_block3a321 = ram_block3a32_PORTADATAOUT_bus[0];

assign ram_block3a322 = ram_block3a32_PORTBDATAOUT_bus[0];

assign ram_block3a01 = ram_block3a0_PORTADATAOUT_bus[0];

assign ram_block3a02 = ram_block3a0_PORTBDATAOUT_bus[0];

assign ram_block3a331 = ram_block3a33_PORTADATAOUT_bus[0];

assign ram_block3a332 = ram_block3a33_PORTBDATAOUT_bus[0];

assign ram_block3a110 = ram_block3a1_PORTADATAOUT_bus[0];

assign ram_block3a111 = ram_block3a1_PORTBDATAOUT_bus[0];

assign ram_block3a341 = ram_block3a34_PORTADATAOUT_bus[0];

assign ram_block3a342 = ram_block3a34_PORTBDATAOUT_bus[0];

assign ram_block3a210 = ram_block3a2_PORTADATAOUT_bus[0];

assign ram_block3a211 = ram_block3a2_PORTBDATAOUT_bus[0];

assign ram_block3a351 = ram_block3a35_PORTADATAOUT_bus[0];

assign ram_block3a352 = ram_block3a35_PORTBDATAOUT_bus[0];

assign ram_block3a310 = ram_block3a3_PORTADATAOUT_bus[0];

assign ram_block3a311 = ram_block3a3_PORTBDATAOUT_bus[0];

assign ram_block3a361 = ram_block3a36_PORTADATAOUT_bus[0];

assign ram_block3a362 = ram_block3a36_PORTBDATAOUT_bus[0];

assign ram_block3a410 = ram_block3a4_PORTADATAOUT_bus[0];

assign ram_block3a411 = ram_block3a4_PORTBDATAOUT_bus[0];

assign ram_block3a371 = ram_block3a37_PORTADATAOUT_bus[0];

assign ram_block3a372 = ram_block3a37_PORTBDATAOUT_bus[0];

assign ram_block3a510 = ram_block3a5_PORTADATAOUT_bus[0];

assign ram_block3a511 = ram_block3a5_PORTBDATAOUT_bus[0];

assign ram_block3a381 = ram_block3a38_PORTADATAOUT_bus[0];

assign ram_block3a382 = ram_block3a38_PORTBDATAOUT_bus[0];

assign ram_block3a64 = ram_block3a6_PORTADATAOUT_bus[0];

assign ram_block3a65 = ram_block3a6_PORTBDATAOUT_bus[0];

assign ram_block3a391 = ram_block3a39_PORTADATAOUT_bus[0];

assign ram_block3a392 = ram_block3a39_PORTBDATAOUT_bus[0];

assign ram_block3a71 = ram_block3a7_PORTADATAOUT_bus[0];

assign ram_block3a72 = ram_block3a7_PORTBDATAOUT_bus[0];

assign ram_block3a401 = ram_block3a40_PORTADATAOUT_bus[0];

assign ram_block3a402 = ram_block3a40_PORTBDATAOUT_bus[0];

assign ram_block3a81 = ram_block3a8_PORTADATAOUT_bus[0];

assign ram_block3a82 = ram_block3a8_PORTBDATAOUT_bus[0];

assign ram_block3a412 = ram_block3a41_PORTADATAOUT_bus[0];

assign ram_block3a413 = ram_block3a41_PORTBDATAOUT_bus[0];

assign ram_block3a91 = ram_block3a9_PORTADATAOUT_bus[0];

assign ram_block3a92 = ram_block3a9_PORTBDATAOUT_bus[0];

assign ram_block3a421 = ram_block3a42_PORTADATAOUT_bus[0];

assign ram_block3a422 = ram_block3a42_PORTBDATAOUT_bus[0];

assign ram_block3a101 = ram_block3a10_PORTADATAOUT_bus[0];

assign ram_block3a102 = ram_block3a10_PORTBDATAOUT_bus[0];

assign ram_block3a431 = ram_block3a43_PORTADATAOUT_bus[0];

assign ram_block3a432 = ram_block3a43_PORTBDATAOUT_bus[0];

assign ram_block3a112 = ram_block3a11_PORTADATAOUT_bus[0];

assign ram_block3a113 = ram_block3a11_PORTBDATAOUT_bus[0];

assign ram_block3a441 = ram_block3a44_PORTADATAOUT_bus[0];

assign ram_block3a442 = ram_block3a44_PORTBDATAOUT_bus[0];

assign ram_block3a121 = ram_block3a12_PORTADATAOUT_bus[0];

assign ram_block3a122 = ram_block3a12_PORTBDATAOUT_bus[0];

assign ram_block3a451 = ram_block3a45_PORTADATAOUT_bus[0];

assign ram_block3a452 = ram_block3a45_PORTBDATAOUT_bus[0];

assign ram_block3a131 = ram_block3a13_PORTADATAOUT_bus[0];

assign ram_block3a132 = ram_block3a13_PORTBDATAOUT_bus[0];

assign ram_block3a461 = ram_block3a46_PORTADATAOUT_bus[0];

assign ram_block3a462 = ram_block3a46_PORTBDATAOUT_bus[0];

assign ram_block3a141 = ram_block3a14_PORTADATAOUT_bus[0];

assign ram_block3a142 = ram_block3a14_PORTBDATAOUT_bus[0];

assign ram_block3a471 = ram_block3a47_PORTADATAOUT_bus[0];

assign ram_block3a472 = ram_block3a47_PORTBDATAOUT_bus[0];

assign ram_block3a151 = ram_block3a15_PORTADATAOUT_bus[0];

assign ram_block3a152 = ram_block3a15_PORTBDATAOUT_bus[0];

assign ram_block3a481 = ram_block3a48_PORTADATAOUT_bus[0];

assign ram_block3a482 = ram_block3a48_PORTBDATAOUT_bus[0];

assign ram_block3a161 = ram_block3a16_PORTADATAOUT_bus[0];

assign ram_block3a162 = ram_block3a16_PORTBDATAOUT_bus[0];

assign ram_block3a491 = ram_block3a49_PORTADATAOUT_bus[0];

assign ram_block3a492 = ram_block3a49_PORTBDATAOUT_bus[0];

assign ram_block3a171 = ram_block3a17_PORTADATAOUT_bus[0];

assign ram_block3a172 = ram_block3a17_PORTBDATAOUT_bus[0];

assign ram_block3a501 = ram_block3a50_PORTADATAOUT_bus[0];

assign ram_block3a502 = ram_block3a50_PORTBDATAOUT_bus[0];

assign ram_block3a181 = ram_block3a18_PORTADATAOUT_bus[0];

assign ram_block3a182 = ram_block3a18_PORTBDATAOUT_bus[0];

assign ram_block3a512 = ram_block3a51_PORTADATAOUT_bus[0];

assign ram_block3a513 = ram_block3a51_PORTBDATAOUT_bus[0];

assign ram_block3a191 = ram_block3a19_PORTADATAOUT_bus[0];

assign ram_block3a192 = ram_block3a19_PORTBDATAOUT_bus[0];

assign ram_block3a521 = ram_block3a52_PORTADATAOUT_bus[0];

assign ram_block3a522 = ram_block3a52_PORTBDATAOUT_bus[0];

assign ram_block3a201 = ram_block3a20_PORTADATAOUT_bus[0];

assign ram_block3a202 = ram_block3a20_PORTBDATAOUT_bus[0];

assign ram_block3a531 = ram_block3a53_PORTADATAOUT_bus[0];

assign ram_block3a532 = ram_block3a53_PORTBDATAOUT_bus[0];

assign ram_block3a212 = ram_block3a21_PORTADATAOUT_bus[0];

assign ram_block3a213 = ram_block3a21_PORTBDATAOUT_bus[0];

assign ram_block3a541 = ram_block3a54_PORTADATAOUT_bus[0];

assign ram_block3a542 = ram_block3a54_PORTBDATAOUT_bus[0];

assign ram_block3a221 = ram_block3a22_PORTADATAOUT_bus[0];

assign ram_block3a222 = ram_block3a22_PORTBDATAOUT_bus[0];

assign ram_block3a551 = ram_block3a55_PORTADATAOUT_bus[0];

assign ram_block3a552 = ram_block3a55_PORTBDATAOUT_bus[0];

assign ram_block3a231 = ram_block3a23_PORTADATAOUT_bus[0];

assign ram_block3a232 = ram_block3a23_PORTBDATAOUT_bus[0];

assign ram_block3a561 = ram_block3a56_PORTADATAOUT_bus[0];

assign ram_block3a562 = ram_block3a56_PORTBDATAOUT_bus[0];

assign ram_block3a241 = ram_block3a24_PORTADATAOUT_bus[0];

assign ram_block3a242 = ram_block3a24_PORTBDATAOUT_bus[0];

assign ram_block3a571 = ram_block3a57_PORTADATAOUT_bus[0];

assign ram_block3a572 = ram_block3a57_PORTBDATAOUT_bus[0];

assign ram_block3a251 = ram_block3a25_PORTADATAOUT_bus[0];

assign ram_block3a252 = ram_block3a25_PORTBDATAOUT_bus[0];

assign ram_block3a581 = ram_block3a58_PORTADATAOUT_bus[0];

assign ram_block3a582 = ram_block3a58_PORTBDATAOUT_bus[0];

assign ram_block3a261 = ram_block3a26_PORTADATAOUT_bus[0];

assign ram_block3a262 = ram_block3a26_PORTBDATAOUT_bus[0];

assign ram_block3a591 = ram_block3a59_PORTADATAOUT_bus[0];

assign ram_block3a592 = ram_block3a59_PORTBDATAOUT_bus[0];

assign ram_block3a271 = ram_block3a27_PORTADATAOUT_bus[0];

assign ram_block3a272 = ram_block3a27_PORTBDATAOUT_bus[0];

assign ram_block3a601 = ram_block3a60_PORTADATAOUT_bus[0];

assign ram_block3a602 = ram_block3a60_PORTBDATAOUT_bus[0];

assign ram_block3a281 = ram_block3a28_PORTADATAOUT_bus[0];

assign ram_block3a282 = ram_block3a28_PORTBDATAOUT_bus[0];

assign ram_block3a611 = ram_block3a61_PORTADATAOUT_bus[0];

assign ram_block3a612 = ram_block3a61_PORTBDATAOUT_bus[0];

assign ram_block3a291 = ram_block3a29_PORTADATAOUT_bus[0];

assign ram_block3a292 = ram_block3a29_PORTBDATAOUT_bus[0];

assign ram_block3a621 = ram_block3a62_PORTADATAOUT_bus[0];

assign ram_block3a622 = ram_block3a62_PORTBDATAOUT_bus[0];

assign ram_block3a301 = ram_block3a30_PORTADATAOUT_bus[0];

assign ram_block3a302 = ram_block3a30_PORTBDATAOUT_bus[0];

assign ram_block3a631 = ram_block3a63_PORTADATAOUT_bus[0];

assign ram_block3a632 = ram_block3a63_PORTBDATAOUT_bus[0];

assign ram_block3a312 = ram_block3a31_PORTADATAOUT_bus[0];

assign ram_block3a313 = ram_block3a31_PORTBDATAOUT_bus[0];

decode_jsa_1 decode5(
	.ram_rom_addr_reg_13(ram_rom_addr_reg_13),
	.sdr(sdr),
	.eq_node_1(\decode5|eq_node[1]~0_combout ),
	.eq_node_0(\decode5|eq_node[0]~1_combout ),
	.irf_reg_2_1(irf_reg_2_1),
	.state_5(state_5),
	.devpor(devpor),
	.devclrn(devclrn),
	.devoe(devoe));

decode_jsa decode4(
	.ramaddr(ramaddr),
	.ramWEN(ramWEN),
	.always1(always1),
	.eq_node_1(\decode4|eq_node[1]~0_combout ),
	.eq_node_0(\decode4|eq_node[0]~1_combout ),
	.devpor(devpor),
	.devclrn(devclrn),
	.devoe(devoe));

// Location: M9K_X51_Y37_N0
cycloneive_ram_block ram_block3a32(
	.portawe(\decode4|eq_node[1]~0_combout ),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(\decode5|eq_node[1]~0_combout ),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock1),
	.ena0(!ramaddr),
	.ena1(ram_rom_addr_reg_13),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({data_a[0]}),
	.portaaddr({address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain({data_b[0]}),
	.portbaddr({address_b[12],address_b[11],address_b[10],address_b[9],address_b[8],address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.devclrn(devclrn),
	.devpor(devpor),
	.portadataout(ram_block3a32_PORTADATAOUT_bus),
	.portbdataout(ram_block3a32_PORTBDATAOUT_bus));
// synopsys translate_off
defparam ram_block3a32.clk0_core_clock_enable = "ena0";
defparam ram_block3a32.clk1_core_clock_enable = "ena1";
defparam ram_block3a32.data_interleave_offset_in_bits = 1;
defparam ram_block3a32.data_interleave_width_in_bits = 1;
defparam ram_block3a32.init_file = "meminit.hex";
defparam ram_block3a32.init_file_layout = "port_a";
defparam ram_block3a32.logical_ram_name = "ram:RAM|altsyncram:altsyncram_component|altsyncram_99f1:auto_generated|altsyncram_fta2:altsyncram1|ALTSYNCRAM";
defparam ram_block3a32.mixed_port_feed_through_mode = "dont_care";
defparam ram_block3a32.operation_mode = "bidir_dual_port";
defparam ram_block3a32.port_a_address_clear = "none";
defparam ram_block3a32.port_a_address_width = 13;
defparam ram_block3a32.port_a_byte_enable_clock = "none";
defparam ram_block3a32.port_a_data_out_clear = "none";
defparam ram_block3a32.port_a_data_out_clock = "none";
defparam ram_block3a32.port_a_data_width = 1;
defparam ram_block3a32.port_a_first_address = 0;
defparam ram_block3a32.port_a_first_bit_number = 0;
defparam ram_block3a32.port_a_last_address = 8191;
defparam ram_block3a32.port_a_logical_ram_depth = 16384;
defparam ram_block3a32.port_a_logical_ram_width = 32;
defparam ram_block3a32.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block3a32.port_b_address_clear = "none";
defparam ram_block3a32.port_b_address_clock = "clock1";
defparam ram_block3a32.port_b_address_width = 13;
defparam ram_block3a32.port_b_data_in_clock = "clock1";
defparam ram_block3a32.port_b_data_out_clear = "none";
defparam ram_block3a32.port_b_data_out_clock = "none";
defparam ram_block3a32.port_b_data_width = 1;
defparam ram_block3a32.port_b_first_address = 0;
defparam ram_block3a32.port_b_first_bit_number = 0;
defparam ram_block3a32.port_b_last_address = 8191;
defparam ram_block3a32.port_b_logical_ram_depth = 16384;
defparam ram_block3a32.port_b_logical_ram_width = 32;
defparam ram_block3a32.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block3a32.port_b_read_enable_clock = "clock1";
defparam ram_block3a32.port_b_write_enable_clock = "clock1";
defparam ram_block3a32.ram_block_type = "M9K";
defparam ram_block3a32.mem_init3 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a32.mem_init2 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a32.mem_init1 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a32.mem_init0 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
// synopsys translate_on

// Location: M9K_X51_Y33_N0
cycloneive_ram_block ram_block3a0(
	.portawe(\decode4|eq_node[0]~1_combout ),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(\decode5|eq_node[0]~1_combout ),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock1),
	.ena0(ramaddr),
	.ena1(!ram_rom_addr_reg_13),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({data_a[0]}),
	.portaaddr({address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain({data_b[0]}),
	.portbaddr({address_b[12],address_b[11],address_b[10],address_b[9],address_b[8],address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.devclrn(devclrn),
	.devpor(devpor),
	.portadataout(ram_block3a0_PORTADATAOUT_bus),
	.portbdataout(ram_block3a0_PORTBDATAOUT_bus));
// synopsys translate_off
defparam ram_block3a0.clk0_core_clock_enable = "ena0";
defparam ram_block3a0.clk1_core_clock_enable = "ena1";
defparam ram_block3a0.data_interleave_offset_in_bits = 1;
defparam ram_block3a0.data_interleave_width_in_bits = 1;
defparam ram_block3a0.init_file = "meminit.hex";
defparam ram_block3a0.init_file_layout = "port_a";
defparam ram_block3a0.logical_ram_name = "ram:RAM|altsyncram:altsyncram_component|altsyncram_99f1:auto_generated|altsyncram_fta2:altsyncram1|ALTSYNCRAM";
defparam ram_block3a0.mixed_port_feed_through_mode = "dont_care";
defparam ram_block3a0.operation_mode = "bidir_dual_port";
defparam ram_block3a0.port_a_address_clear = "none";
defparam ram_block3a0.port_a_address_width = 13;
defparam ram_block3a0.port_a_byte_enable_clock = "none";
defparam ram_block3a0.port_a_data_out_clear = "none";
defparam ram_block3a0.port_a_data_out_clock = "none";
defparam ram_block3a0.port_a_data_width = 1;
defparam ram_block3a0.port_a_first_address = 0;
defparam ram_block3a0.port_a_first_bit_number = 0;
defparam ram_block3a0.port_a_last_address = 8191;
defparam ram_block3a0.port_a_logical_ram_depth = 16384;
defparam ram_block3a0.port_a_logical_ram_width = 32;
defparam ram_block3a0.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block3a0.port_b_address_clear = "none";
defparam ram_block3a0.port_b_address_clock = "clock1";
defparam ram_block3a0.port_b_address_width = 13;
defparam ram_block3a0.port_b_data_in_clock = "clock1";
defparam ram_block3a0.port_b_data_out_clear = "none";
defparam ram_block3a0.port_b_data_out_clock = "none";
defparam ram_block3a0.port_b_data_width = 1;
defparam ram_block3a0.port_b_first_address = 0;
defparam ram_block3a0.port_b_first_bit_number = 0;
defparam ram_block3a0.port_b_last_address = 8191;
defparam ram_block3a0.port_b_logical_ram_depth = 16384;
defparam ram_block3a0.port_b_logical_ram_width = 32;
defparam ram_block3a0.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block3a0.port_b_read_enable_clock = "clock1";
defparam ram_block3a0.port_b_write_enable_clock = "clock1";
defparam ram_block3a0.ram_block_type = "M9K";
defparam ram_block3a0.mem_init3 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a0.mem_init2 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a0.mem_init1 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a0.mem_init0 = 2048'h0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001802C7EA14A7EF95C00000000000000000000000000000A242111E008528F7260;
// synopsys translate_on

// Location: M9K_X51_Y25_N0
cycloneive_ram_block ram_block3a33(
	.portawe(\decode4|eq_node[1]~0_combout ),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(\decode5|eq_node[1]~0_combout ),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock1),
	.ena0(!ramaddr),
	.ena1(ram_rom_addr_reg_13),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({data_a[1]}),
	.portaaddr({address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain({data_b[1]}),
	.portbaddr({address_b[12],address_b[11],address_b[10],address_b[9],address_b[8],address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.devclrn(devclrn),
	.devpor(devpor),
	.portadataout(ram_block3a33_PORTADATAOUT_bus),
	.portbdataout(ram_block3a33_PORTBDATAOUT_bus));
// synopsys translate_off
defparam ram_block3a33.clk0_core_clock_enable = "ena0";
defparam ram_block3a33.clk1_core_clock_enable = "ena1";
defparam ram_block3a33.data_interleave_offset_in_bits = 1;
defparam ram_block3a33.data_interleave_width_in_bits = 1;
defparam ram_block3a33.init_file = "meminit.hex";
defparam ram_block3a33.init_file_layout = "port_a";
defparam ram_block3a33.logical_ram_name = "ram:RAM|altsyncram:altsyncram_component|altsyncram_99f1:auto_generated|altsyncram_fta2:altsyncram1|ALTSYNCRAM";
defparam ram_block3a33.mixed_port_feed_through_mode = "dont_care";
defparam ram_block3a33.operation_mode = "bidir_dual_port";
defparam ram_block3a33.port_a_address_clear = "none";
defparam ram_block3a33.port_a_address_width = 13;
defparam ram_block3a33.port_a_byte_enable_clock = "none";
defparam ram_block3a33.port_a_data_out_clear = "none";
defparam ram_block3a33.port_a_data_out_clock = "none";
defparam ram_block3a33.port_a_data_width = 1;
defparam ram_block3a33.port_a_first_address = 0;
defparam ram_block3a33.port_a_first_bit_number = 1;
defparam ram_block3a33.port_a_last_address = 8191;
defparam ram_block3a33.port_a_logical_ram_depth = 16384;
defparam ram_block3a33.port_a_logical_ram_width = 32;
defparam ram_block3a33.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block3a33.port_b_address_clear = "none";
defparam ram_block3a33.port_b_address_clock = "clock1";
defparam ram_block3a33.port_b_address_width = 13;
defparam ram_block3a33.port_b_data_in_clock = "clock1";
defparam ram_block3a33.port_b_data_out_clear = "none";
defparam ram_block3a33.port_b_data_out_clock = "none";
defparam ram_block3a33.port_b_data_width = 1;
defparam ram_block3a33.port_b_first_address = 0;
defparam ram_block3a33.port_b_first_bit_number = 1;
defparam ram_block3a33.port_b_last_address = 8191;
defparam ram_block3a33.port_b_logical_ram_depth = 16384;
defparam ram_block3a33.port_b_logical_ram_width = 32;
defparam ram_block3a33.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block3a33.port_b_read_enable_clock = "clock1";
defparam ram_block3a33.port_b_write_enable_clock = "clock1";
defparam ram_block3a33.ram_block_type = "M9K";
defparam ram_block3a33.mem_init3 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a33.mem_init2 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a33.mem_init1 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a33.mem_init0 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
// synopsys translate_on

// Location: M9K_X37_Y25_N0
cycloneive_ram_block ram_block3a1(
	.portawe(\decode4|eq_node[0]~1_combout ),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(\decode5|eq_node[0]~1_combout ),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock1),
	.ena0(ramaddr),
	.ena1(!ram_rom_addr_reg_13),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({data_a[1]}),
	.portaaddr({address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain({data_b[1]}),
	.portbaddr({address_b[12],address_b[11],address_b[10],address_b[9],address_b[8],address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.devclrn(devclrn),
	.devpor(devpor),
	.portadataout(ram_block3a1_PORTADATAOUT_bus),
	.portbdataout(ram_block3a1_PORTBDATAOUT_bus));
// synopsys translate_off
defparam ram_block3a1.clk0_core_clock_enable = "ena0";
defparam ram_block3a1.clk1_core_clock_enable = "ena1";
defparam ram_block3a1.data_interleave_offset_in_bits = 1;
defparam ram_block3a1.data_interleave_width_in_bits = 1;
defparam ram_block3a1.init_file = "meminit.hex";
defparam ram_block3a1.init_file_layout = "port_a";
defparam ram_block3a1.logical_ram_name = "ram:RAM|altsyncram:altsyncram_component|altsyncram_99f1:auto_generated|altsyncram_fta2:altsyncram1|ALTSYNCRAM";
defparam ram_block3a1.mixed_port_feed_through_mode = "dont_care";
defparam ram_block3a1.operation_mode = "bidir_dual_port";
defparam ram_block3a1.port_a_address_clear = "none";
defparam ram_block3a1.port_a_address_width = 13;
defparam ram_block3a1.port_a_byte_enable_clock = "none";
defparam ram_block3a1.port_a_data_out_clear = "none";
defparam ram_block3a1.port_a_data_out_clock = "none";
defparam ram_block3a1.port_a_data_width = 1;
defparam ram_block3a1.port_a_first_address = 0;
defparam ram_block3a1.port_a_first_bit_number = 1;
defparam ram_block3a1.port_a_last_address = 8191;
defparam ram_block3a1.port_a_logical_ram_depth = 16384;
defparam ram_block3a1.port_a_logical_ram_width = 32;
defparam ram_block3a1.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block3a1.port_b_address_clear = "none";
defparam ram_block3a1.port_b_address_clock = "clock1";
defparam ram_block3a1.port_b_address_width = 13;
defparam ram_block3a1.port_b_data_in_clock = "clock1";
defparam ram_block3a1.port_b_data_out_clear = "none";
defparam ram_block3a1.port_b_data_out_clock = "none";
defparam ram_block3a1.port_b_data_width = 1;
defparam ram_block3a1.port_b_first_address = 0;
defparam ram_block3a1.port_b_first_bit_number = 1;
defparam ram_block3a1.port_b_last_address = 8191;
defparam ram_block3a1.port_b_logical_ram_depth = 16384;
defparam ram_block3a1.port_b_logical_ram_width = 32;
defparam ram_block3a1.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block3a1.port_b_read_enable_clock = "clock1";
defparam ram_block3a1.port_b_write_enable_clock = "clock1";
defparam ram_block3a1.ram_block_type = "M9K";
defparam ram_block3a1.mem_init3 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a1.mem_init2 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a1.mem_init1 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a1.mem_init0 = 2048'h0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001D4AE6429116B3C8A000000000000000000000000000012242108900D12808390;
// synopsys translate_on

// Location: M9K_X51_Y23_N0
cycloneive_ram_block ram_block3a34(
	.portawe(\decode4|eq_node[1]~0_combout ),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(\decode5|eq_node[1]~0_combout ),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock1),
	.ena0(!ramaddr),
	.ena1(ram_rom_addr_reg_13),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({data_a[2]}),
	.portaaddr({address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain({data_b[2]}),
	.portbaddr({address_b[12],address_b[11],address_b[10],address_b[9],address_b[8],address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.devclrn(devclrn),
	.devpor(devpor),
	.portadataout(ram_block3a34_PORTADATAOUT_bus),
	.portbdataout(ram_block3a34_PORTBDATAOUT_bus));
// synopsys translate_off
defparam ram_block3a34.clk0_core_clock_enable = "ena0";
defparam ram_block3a34.clk1_core_clock_enable = "ena1";
defparam ram_block3a34.data_interleave_offset_in_bits = 1;
defparam ram_block3a34.data_interleave_width_in_bits = 1;
defparam ram_block3a34.init_file = "meminit.hex";
defparam ram_block3a34.init_file_layout = "port_a";
defparam ram_block3a34.logical_ram_name = "ram:RAM|altsyncram:altsyncram_component|altsyncram_99f1:auto_generated|altsyncram_fta2:altsyncram1|ALTSYNCRAM";
defparam ram_block3a34.mixed_port_feed_through_mode = "dont_care";
defparam ram_block3a34.operation_mode = "bidir_dual_port";
defparam ram_block3a34.port_a_address_clear = "none";
defparam ram_block3a34.port_a_address_width = 13;
defparam ram_block3a34.port_a_byte_enable_clock = "none";
defparam ram_block3a34.port_a_data_out_clear = "none";
defparam ram_block3a34.port_a_data_out_clock = "none";
defparam ram_block3a34.port_a_data_width = 1;
defparam ram_block3a34.port_a_first_address = 0;
defparam ram_block3a34.port_a_first_bit_number = 2;
defparam ram_block3a34.port_a_last_address = 8191;
defparam ram_block3a34.port_a_logical_ram_depth = 16384;
defparam ram_block3a34.port_a_logical_ram_width = 32;
defparam ram_block3a34.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block3a34.port_b_address_clear = "none";
defparam ram_block3a34.port_b_address_clock = "clock1";
defparam ram_block3a34.port_b_address_width = 13;
defparam ram_block3a34.port_b_data_in_clock = "clock1";
defparam ram_block3a34.port_b_data_out_clear = "none";
defparam ram_block3a34.port_b_data_out_clock = "none";
defparam ram_block3a34.port_b_data_width = 1;
defparam ram_block3a34.port_b_first_address = 0;
defparam ram_block3a34.port_b_first_bit_number = 2;
defparam ram_block3a34.port_b_last_address = 8191;
defparam ram_block3a34.port_b_logical_ram_depth = 16384;
defparam ram_block3a34.port_b_logical_ram_width = 32;
defparam ram_block3a34.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block3a34.port_b_read_enable_clock = "clock1";
defparam ram_block3a34.port_b_write_enable_clock = "clock1";
defparam ram_block3a34.ram_block_type = "M9K";
defparam ram_block3a34.mem_init3 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a34.mem_init2 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a34.mem_init1 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a34.mem_init0 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
// synopsys translate_on

// Location: M9K_X64_Y25_N0
cycloneive_ram_block ram_block3a2(
	.portawe(\decode4|eq_node[0]~1_combout ),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(\decode5|eq_node[0]~1_combout ),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock1),
	.ena0(ramaddr),
	.ena1(!ram_rom_addr_reg_13),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({data_a[2]}),
	.portaaddr({address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain({data_b[2]}),
	.portbaddr({address_b[12],address_b[11],address_b[10],address_b[9],address_b[8],address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.devclrn(devclrn),
	.devpor(devpor),
	.portadataout(ram_block3a2_PORTADATAOUT_bus),
	.portbdataout(ram_block3a2_PORTBDATAOUT_bus));
// synopsys translate_off
defparam ram_block3a2.clk0_core_clock_enable = "ena0";
defparam ram_block3a2.clk1_core_clock_enable = "ena1";
defparam ram_block3a2.data_interleave_offset_in_bits = 1;
defparam ram_block3a2.data_interleave_width_in_bits = 1;
defparam ram_block3a2.init_file = "meminit.hex";
defparam ram_block3a2.init_file_layout = "port_a";
defparam ram_block3a2.logical_ram_name = "ram:RAM|altsyncram:altsyncram_component|altsyncram_99f1:auto_generated|altsyncram_fta2:altsyncram1|ALTSYNCRAM";
defparam ram_block3a2.mixed_port_feed_through_mode = "dont_care";
defparam ram_block3a2.operation_mode = "bidir_dual_port";
defparam ram_block3a2.port_a_address_clear = "none";
defparam ram_block3a2.port_a_address_width = 13;
defparam ram_block3a2.port_a_byte_enable_clock = "none";
defparam ram_block3a2.port_a_data_out_clear = "none";
defparam ram_block3a2.port_a_data_out_clock = "none";
defparam ram_block3a2.port_a_data_width = 1;
defparam ram_block3a2.port_a_first_address = 0;
defparam ram_block3a2.port_a_first_bit_number = 2;
defparam ram_block3a2.port_a_last_address = 8191;
defparam ram_block3a2.port_a_logical_ram_depth = 16384;
defparam ram_block3a2.port_a_logical_ram_width = 32;
defparam ram_block3a2.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block3a2.port_b_address_clear = "none";
defparam ram_block3a2.port_b_address_clock = "clock1";
defparam ram_block3a2.port_b_address_width = 13;
defparam ram_block3a2.port_b_data_in_clock = "clock1";
defparam ram_block3a2.port_b_data_out_clear = "none";
defparam ram_block3a2.port_b_data_out_clock = "none";
defparam ram_block3a2.port_b_data_width = 1;
defparam ram_block3a2.port_b_first_address = 0;
defparam ram_block3a2.port_b_first_bit_number = 2;
defparam ram_block3a2.port_b_last_address = 8191;
defparam ram_block3a2.port_b_logical_ram_depth = 16384;
defparam ram_block3a2.port_b_logical_ram_width = 32;
defparam ram_block3a2.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block3a2.port_b_read_enable_clock = "clock1";
defparam ram_block3a2.port_b_write_enable_clock = "clock1";
defparam ram_block3a2.ram_block_type = "M9K";
defparam ram_block3a2.mem_init3 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a2.mem_init2 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a2.mem_init1 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a2.mem_init0 = 2048'h0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000961CA470728D97800000000000000000000000000000172E7BD1C323272F6867;
// synopsys translate_on

// Location: M9K_X51_Y30_N0
cycloneive_ram_block ram_block3a35(
	.portawe(\decode4|eq_node[1]~0_combout ),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(\decode5|eq_node[1]~0_combout ),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock1),
	.ena0(!ramaddr),
	.ena1(ram_rom_addr_reg_13),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({data_a[3]}),
	.portaaddr({address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain({data_b[3]}),
	.portbaddr({address_b[12],address_b[11],address_b[10],address_b[9],address_b[8],address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.devclrn(devclrn),
	.devpor(devpor),
	.portadataout(ram_block3a35_PORTADATAOUT_bus),
	.portbdataout(ram_block3a35_PORTBDATAOUT_bus));
// synopsys translate_off
defparam ram_block3a35.clk0_core_clock_enable = "ena0";
defparam ram_block3a35.clk1_core_clock_enable = "ena1";
defparam ram_block3a35.data_interleave_offset_in_bits = 1;
defparam ram_block3a35.data_interleave_width_in_bits = 1;
defparam ram_block3a35.init_file = "meminit.hex";
defparam ram_block3a35.init_file_layout = "port_a";
defparam ram_block3a35.logical_ram_name = "ram:RAM|altsyncram:altsyncram_component|altsyncram_99f1:auto_generated|altsyncram_fta2:altsyncram1|ALTSYNCRAM";
defparam ram_block3a35.mixed_port_feed_through_mode = "dont_care";
defparam ram_block3a35.operation_mode = "bidir_dual_port";
defparam ram_block3a35.port_a_address_clear = "none";
defparam ram_block3a35.port_a_address_width = 13;
defparam ram_block3a35.port_a_byte_enable_clock = "none";
defparam ram_block3a35.port_a_data_out_clear = "none";
defparam ram_block3a35.port_a_data_out_clock = "none";
defparam ram_block3a35.port_a_data_width = 1;
defparam ram_block3a35.port_a_first_address = 0;
defparam ram_block3a35.port_a_first_bit_number = 3;
defparam ram_block3a35.port_a_last_address = 8191;
defparam ram_block3a35.port_a_logical_ram_depth = 16384;
defparam ram_block3a35.port_a_logical_ram_width = 32;
defparam ram_block3a35.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block3a35.port_b_address_clear = "none";
defparam ram_block3a35.port_b_address_clock = "clock1";
defparam ram_block3a35.port_b_address_width = 13;
defparam ram_block3a35.port_b_data_in_clock = "clock1";
defparam ram_block3a35.port_b_data_out_clear = "none";
defparam ram_block3a35.port_b_data_out_clock = "none";
defparam ram_block3a35.port_b_data_width = 1;
defparam ram_block3a35.port_b_first_address = 0;
defparam ram_block3a35.port_b_first_bit_number = 3;
defparam ram_block3a35.port_b_last_address = 8191;
defparam ram_block3a35.port_b_logical_ram_depth = 16384;
defparam ram_block3a35.port_b_logical_ram_width = 32;
defparam ram_block3a35.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block3a35.port_b_read_enable_clock = "clock1";
defparam ram_block3a35.port_b_write_enable_clock = "clock1";
defparam ram_block3a35.ram_block_type = "M9K";
defparam ram_block3a35.mem_init3 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a35.mem_init2 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a35.mem_init1 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a35.mem_init0 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
// synopsys translate_on

// Location: M9K_X51_Y31_N0
cycloneive_ram_block ram_block3a3(
	.portawe(\decode4|eq_node[0]~1_combout ),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(\decode5|eq_node[0]~1_combout ),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock1),
	.ena0(ramaddr),
	.ena1(!ram_rom_addr_reg_13),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({data_a[3]}),
	.portaaddr({address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain({data_b[3]}),
	.portbaddr({address_b[12],address_b[11],address_b[10],address_b[9],address_b[8],address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.devclrn(devclrn),
	.devpor(devpor),
	.portadataout(ram_block3a3_PORTADATAOUT_bus),
	.portbdataout(ram_block3a3_PORTBDATAOUT_bus));
// synopsys translate_off
defparam ram_block3a3.clk0_core_clock_enable = "ena0";
defparam ram_block3a3.clk1_core_clock_enable = "ena1";
defparam ram_block3a3.data_interleave_offset_in_bits = 1;
defparam ram_block3a3.data_interleave_width_in_bits = 1;
defparam ram_block3a3.init_file = "meminit.hex";
defparam ram_block3a3.init_file_layout = "port_a";
defparam ram_block3a3.logical_ram_name = "ram:RAM|altsyncram:altsyncram_component|altsyncram_99f1:auto_generated|altsyncram_fta2:altsyncram1|ALTSYNCRAM";
defparam ram_block3a3.mixed_port_feed_through_mode = "dont_care";
defparam ram_block3a3.operation_mode = "bidir_dual_port";
defparam ram_block3a3.port_a_address_clear = "none";
defparam ram_block3a3.port_a_address_width = 13;
defparam ram_block3a3.port_a_byte_enable_clock = "none";
defparam ram_block3a3.port_a_data_out_clear = "none";
defparam ram_block3a3.port_a_data_out_clock = "none";
defparam ram_block3a3.port_a_data_width = 1;
defparam ram_block3a3.port_a_first_address = 0;
defparam ram_block3a3.port_a_first_bit_number = 3;
defparam ram_block3a3.port_a_last_address = 8191;
defparam ram_block3a3.port_a_logical_ram_depth = 16384;
defparam ram_block3a3.port_a_logical_ram_width = 32;
defparam ram_block3a3.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block3a3.port_b_address_clear = "none";
defparam ram_block3a3.port_b_address_clock = "clock1";
defparam ram_block3a3.port_b_address_width = 13;
defparam ram_block3a3.port_b_data_in_clock = "clock1";
defparam ram_block3a3.port_b_data_out_clear = "none";
defparam ram_block3a3.port_b_data_out_clock = "none";
defparam ram_block3a3.port_b_data_width = 1;
defparam ram_block3a3.port_b_first_address = 0;
defparam ram_block3a3.port_b_first_bit_number = 3;
defparam ram_block3a3.port_b_last_address = 8191;
defparam ram_block3a3.port_b_logical_ram_depth = 16384;
defparam ram_block3a3.port_b_logical_ram_width = 32;
defparam ram_block3a3.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block3a3.port_b_read_enable_clock = "clock1";
defparam ram_block3a3.port_b_write_enable_clock = "clock1";
defparam ram_block3a3.ram_block_type = "M9K";
defparam ram_block3a3.mem_init3 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a3.mem_init2 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a3.mem_init1 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a3.mem_init0 = 2048'h000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000009F20E64C2468E52000000000000000000000000000022346308C62632A08083;
// synopsys translate_on

// Location: M9K_X51_Y28_N0
cycloneive_ram_block ram_block3a36(
	.portawe(\decode4|eq_node[1]~0_combout ),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(\decode5|eq_node[1]~0_combout ),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock1),
	.ena0(!ramaddr),
	.ena1(ram_rom_addr_reg_13),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({data_a[4]}),
	.portaaddr({address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain({data_b[4]}),
	.portbaddr({address_b[12],address_b[11],address_b[10],address_b[9],address_b[8],address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.devclrn(devclrn),
	.devpor(devpor),
	.portadataout(ram_block3a36_PORTADATAOUT_bus),
	.portbdataout(ram_block3a36_PORTBDATAOUT_bus));
// synopsys translate_off
defparam ram_block3a36.clk0_core_clock_enable = "ena0";
defparam ram_block3a36.clk1_core_clock_enable = "ena1";
defparam ram_block3a36.data_interleave_offset_in_bits = 1;
defparam ram_block3a36.data_interleave_width_in_bits = 1;
defparam ram_block3a36.init_file = "meminit.hex";
defparam ram_block3a36.init_file_layout = "port_a";
defparam ram_block3a36.logical_ram_name = "ram:RAM|altsyncram:altsyncram_component|altsyncram_99f1:auto_generated|altsyncram_fta2:altsyncram1|ALTSYNCRAM";
defparam ram_block3a36.mixed_port_feed_through_mode = "dont_care";
defparam ram_block3a36.operation_mode = "bidir_dual_port";
defparam ram_block3a36.port_a_address_clear = "none";
defparam ram_block3a36.port_a_address_width = 13;
defparam ram_block3a36.port_a_byte_enable_clock = "none";
defparam ram_block3a36.port_a_data_out_clear = "none";
defparam ram_block3a36.port_a_data_out_clock = "none";
defparam ram_block3a36.port_a_data_width = 1;
defparam ram_block3a36.port_a_first_address = 0;
defparam ram_block3a36.port_a_first_bit_number = 4;
defparam ram_block3a36.port_a_last_address = 8191;
defparam ram_block3a36.port_a_logical_ram_depth = 16384;
defparam ram_block3a36.port_a_logical_ram_width = 32;
defparam ram_block3a36.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block3a36.port_b_address_clear = "none";
defparam ram_block3a36.port_b_address_clock = "clock1";
defparam ram_block3a36.port_b_address_width = 13;
defparam ram_block3a36.port_b_data_in_clock = "clock1";
defparam ram_block3a36.port_b_data_out_clear = "none";
defparam ram_block3a36.port_b_data_out_clock = "none";
defparam ram_block3a36.port_b_data_width = 1;
defparam ram_block3a36.port_b_first_address = 0;
defparam ram_block3a36.port_b_first_bit_number = 4;
defparam ram_block3a36.port_b_last_address = 8191;
defparam ram_block3a36.port_b_logical_ram_depth = 16384;
defparam ram_block3a36.port_b_logical_ram_width = 32;
defparam ram_block3a36.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block3a36.port_b_read_enable_clock = "clock1";
defparam ram_block3a36.port_b_write_enable_clock = "clock1";
defparam ram_block3a36.ram_block_type = "M9K";
defparam ram_block3a36.mem_init3 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a36.mem_init2 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a36.mem_init1 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a36.mem_init0 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
// synopsys translate_on

// Location: M9K_X51_Y27_N0
cycloneive_ram_block ram_block3a4(
	.portawe(\decode4|eq_node[0]~1_combout ),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(\decode5|eq_node[0]~1_combout ),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock1),
	.ena0(ramaddr),
	.ena1(!ram_rom_addr_reg_13),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({data_a[4]}),
	.portaaddr({address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain({data_b[4]}),
	.portbaddr({address_b[12],address_b[11],address_b[10],address_b[9],address_b[8],address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.devclrn(devclrn),
	.devpor(devpor),
	.portadataout(ram_block3a4_PORTADATAOUT_bus),
	.portbdataout(ram_block3a4_PORTBDATAOUT_bus));
// synopsys translate_off
defparam ram_block3a4.clk0_core_clock_enable = "ena0";
defparam ram_block3a4.clk1_core_clock_enable = "ena1";
defparam ram_block3a4.data_interleave_offset_in_bits = 1;
defparam ram_block3a4.data_interleave_width_in_bits = 1;
defparam ram_block3a4.init_file = "meminit.hex";
defparam ram_block3a4.init_file_layout = "port_a";
defparam ram_block3a4.logical_ram_name = "ram:RAM|altsyncram:altsyncram_component|altsyncram_99f1:auto_generated|altsyncram_fta2:altsyncram1|ALTSYNCRAM";
defparam ram_block3a4.mixed_port_feed_through_mode = "dont_care";
defparam ram_block3a4.operation_mode = "bidir_dual_port";
defparam ram_block3a4.port_a_address_clear = "none";
defparam ram_block3a4.port_a_address_width = 13;
defparam ram_block3a4.port_a_byte_enable_clock = "none";
defparam ram_block3a4.port_a_data_out_clear = "none";
defparam ram_block3a4.port_a_data_out_clock = "none";
defparam ram_block3a4.port_a_data_width = 1;
defparam ram_block3a4.port_a_first_address = 0;
defparam ram_block3a4.port_a_first_bit_number = 4;
defparam ram_block3a4.port_a_last_address = 8191;
defparam ram_block3a4.port_a_logical_ram_depth = 16384;
defparam ram_block3a4.port_a_logical_ram_width = 32;
defparam ram_block3a4.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block3a4.port_b_address_clear = "none";
defparam ram_block3a4.port_b_address_clock = "clock1";
defparam ram_block3a4.port_b_address_width = 13;
defparam ram_block3a4.port_b_data_in_clock = "clock1";
defparam ram_block3a4.port_b_data_out_clear = "none";
defparam ram_block3a4.port_b_data_out_clock = "none";
defparam ram_block3a4.port_b_data_width = 1;
defparam ram_block3a4.port_b_first_address = 0;
defparam ram_block3a4.port_b_first_bit_number = 4;
defparam ram_block3a4.port_b_last_address = 8191;
defparam ram_block3a4.port_b_logical_ram_depth = 16384;
defparam ram_block3a4.port_b_logical_ram_width = 32;
defparam ram_block3a4.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block3a4.port_b_read_enable_clock = "clock1";
defparam ram_block3a4.port_b_write_enable_clock = "clock1";
defparam ram_block3a4.ram_block_type = "M9K";
defparam ram_block3a4.mem_init3 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a4.mem_init2 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a4.mem_init1 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a4.mem_init0 = 2048'h000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000060B81842D24565BE000000000000000000000000000002242101022202208083;
// synopsys translate_on

// Location: M9K_X51_Y36_N0
cycloneive_ram_block ram_block3a37(
	.portawe(\decode4|eq_node[1]~0_combout ),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(\decode5|eq_node[1]~0_combout ),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock1),
	.ena0(!ramaddr),
	.ena1(ram_rom_addr_reg_13),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({data_a[5]}),
	.portaaddr({address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain({data_b[5]}),
	.portbaddr({address_b[12],address_b[11],address_b[10],address_b[9],address_b[8],address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.devclrn(devclrn),
	.devpor(devpor),
	.portadataout(ram_block3a37_PORTADATAOUT_bus),
	.portbdataout(ram_block3a37_PORTBDATAOUT_bus));
// synopsys translate_off
defparam ram_block3a37.clk0_core_clock_enable = "ena0";
defparam ram_block3a37.clk1_core_clock_enable = "ena1";
defparam ram_block3a37.data_interleave_offset_in_bits = 1;
defparam ram_block3a37.data_interleave_width_in_bits = 1;
defparam ram_block3a37.init_file = "meminit.hex";
defparam ram_block3a37.init_file_layout = "port_a";
defparam ram_block3a37.logical_ram_name = "ram:RAM|altsyncram:altsyncram_component|altsyncram_99f1:auto_generated|altsyncram_fta2:altsyncram1|ALTSYNCRAM";
defparam ram_block3a37.mixed_port_feed_through_mode = "dont_care";
defparam ram_block3a37.operation_mode = "bidir_dual_port";
defparam ram_block3a37.port_a_address_clear = "none";
defparam ram_block3a37.port_a_address_width = 13;
defparam ram_block3a37.port_a_byte_enable_clock = "none";
defparam ram_block3a37.port_a_data_out_clear = "none";
defparam ram_block3a37.port_a_data_out_clock = "none";
defparam ram_block3a37.port_a_data_width = 1;
defparam ram_block3a37.port_a_first_address = 0;
defparam ram_block3a37.port_a_first_bit_number = 5;
defparam ram_block3a37.port_a_last_address = 8191;
defparam ram_block3a37.port_a_logical_ram_depth = 16384;
defparam ram_block3a37.port_a_logical_ram_width = 32;
defparam ram_block3a37.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block3a37.port_b_address_clear = "none";
defparam ram_block3a37.port_b_address_clock = "clock1";
defparam ram_block3a37.port_b_address_width = 13;
defparam ram_block3a37.port_b_data_in_clock = "clock1";
defparam ram_block3a37.port_b_data_out_clear = "none";
defparam ram_block3a37.port_b_data_out_clock = "none";
defparam ram_block3a37.port_b_data_width = 1;
defparam ram_block3a37.port_b_first_address = 0;
defparam ram_block3a37.port_b_first_bit_number = 5;
defparam ram_block3a37.port_b_last_address = 8191;
defparam ram_block3a37.port_b_logical_ram_depth = 16384;
defparam ram_block3a37.port_b_logical_ram_width = 32;
defparam ram_block3a37.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block3a37.port_b_read_enable_clock = "clock1";
defparam ram_block3a37.port_b_write_enable_clock = "clock1";
defparam ram_block3a37.ram_block_type = "M9K";
defparam ram_block3a37.mem_init3 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a37.mem_init2 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a37.mem_init1 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a37.mem_init0 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
// synopsys translate_on

// Location: M9K_X51_Y39_N0
cycloneive_ram_block ram_block3a5(
	.portawe(\decode4|eq_node[0]~1_combout ),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(\decode5|eq_node[0]~1_combout ),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock1),
	.ena0(ramaddr),
	.ena1(!ram_rom_addr_reg_13),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({data_a[5]}),
	.portaaddr({address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain({data_b[5]}),
	.portbaddr({address_b[12],address_b[11],address_b[10],address_b[9],address_b[8],address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.devclrn(devclrn),
	.devpor(devpor),
	.portadataout(ram_block3a5_PORTADATAOUT_bus),
	.portbdataout(ram_block3a5_PORTBDATAOUT_bus));
// synopsys translate_off
defparam ram_block3a5.clk0_core_clock_enable = "ena0";
defparam ram_block3a5.clk1_core_clock_enable = "ena1";
defparam ram_block3a5.data_interleave_offset_in_bits = 1;
defparam ram_block3a5.data_interleave_width_in_bits = 1;
defparam ram_block3a5.init_file = "meminit.hex";
defparam ram_block3a5.init_file_layout = "port_a";
defparam ram_block3a5.logical_ram_name = "ram:RAM|altsyncram:altsyncram_component|altsyncram_99f1:auto_generated|altsyncram_fta2:altsyncram1|ALTSYNCRAM";
defparam ram_block3a5.mixed_port_feed_through_mode = "dont_care";
defparam ram_block3a5.operation_mode = "bidir_dual_port";
defparam ram_block3a5.port_a_address_clear = "none";
defparam ram_block3a5.port_a_address_width = 13;
defparam ram_block3a5.port_a_byte_enable_clock = "none";
defparam ram_block3a5.port_a_data_out_clear = "none";
defparam ram_block3a5.port_a_data_out_clock = "none";
defparam ram_block3a5.port_a_data_width = 1;
defparam ram_block3a5.port_a_first_address = 0;
defparam ram_block3a5.port_a_first_bit_number = 5;
defparam ram_block3a5.port_a_last_address = 8191;
defparam ram_block3a5.port_a_logical_ram_depth = 16384;
defparam ram_block3a5.port_a_logical_ram_width = 32;
defparam ram_block3a5.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block3a5.port_b_address_clear = "none";
defparam ram_block3a5.port_b_address_clock = "clock1";
defparam ram_block3a5.port_b_address_width = 13;
defparam ram_block3a5.port_b_data_in_clock = "clock1";
defparam ram_block3a5.port_b_data_out_clear = "none";
defparam ram_block3a5.port_b_data_out_clock = "none";
defparam ram_block3a5.port_b_data_width = 1;
defparam ram_block3a5.port_b_first_address = 0;
defparam ram_block3a5.port_b_first_bit_number = 5;
defparam ram_block3a5.port_b_last_address = 8191;
defparam ram_block3a5.port_b_logical_ram_depth = 16384;
defparam ram_block3a5.port_b_logical_ram_width = 32;
defparam ram_block3a5.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block3a5.port_b_read_enable_clock = "clock1";
defparam ram_block3a5.port_b_write_enable_clock = "clock1";
defparam ram_block3a5.ram_block_type = "M9K";
defparam ram_block3a5.mem_init3 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a5.mem_init2 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a5.mem_init1 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a5.mem_init0 = 2048'h000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000056414512D6B00448000000000000000000000000000002246308006652AF7263;
// synopsys translate_on

// Location: M9K_X51_Y29_N0
cycloneive_ram_block ram_block3a38(
	.portawe(\decode4|eq_node[1]~0_combout ),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(\decode5|eq_node[1]~0_combout ),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock1),
	.ena0(!ramaddr),
	.ena1(ram_rom_addr_reg_13),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({data_a[6]}),
	.portaaddr({address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain({data_b[6]}),
	.portbaddr({address_b[12],address_b[11],address_b[10],address_b[9],address_b[8],address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.devclrn(devclrn),
	.devpor(devpor),
	.portadataout(ram_block3a38_PORTADATAOUT_bus),
	.portbdataout(ram_block3a38_PORTBDATAOUT_bus));
// synopsys translate_off
defparam ram_block3a38.clk0_core_clock_enable = "ena0";
defparam ram_block3a38.clk1_core_clock_enable = "ena1";
defparam ram_block3a38.data_interleave_offset_in_bits = 1;
defparam ram_block3a38.data_interleave_width_in_bits = 1;
defparam ram_block3a38.init_file = "meminit.hex";
defparam ram_block3a38.init_file_layout = "port_a";
defparam ram_block3a38.logical_ram_name = "ram:RAM|altsyncram:altsyncram_component|altsyncram_99f1:auto_generated|altsyncram_fta2:altsyncram1|ALTSYNCRAM";
defparam ram_block3a38.mixed_port_feed_through_mode = "dont_care";
defparam ram_block3a38.operation_mode = "bidir_dual_port";
defparam ram_block3a38.port_a_address_clear = "none";
defparam ram_block3a38.port_a_address_width = 13;
defparam ram_block3a38.port_a_byte_enable_clock = "none";
defparam ram_block3a38.port_a_data_out_clear = "none";
defparam ram_block3a38.port_a_data_out_clock = "none";
defparam ram_block3a38.port_a_data_width = 1;
defparam ram_block3a38.port_a_first_address = 0;
defparam ram_block3a38.port_a_first_bit_number = 6;
defparam ram_block3a38.port_a_last_address = 8191;
defparam ram_block3a38.port_a_logical_ram_depth = 16384;
defparam ram_block3a38.port_a_logical_ram_width = 32;
defparam ram_block3a38.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block3a38.port_b_address_clear = "none";
defparam ram_block3a38.port_b_address_clock = "clock1";
defparam ram_block3a38.port_b_address_width = 13;
defparam ram_block3a38.port_b_data_in_clock = "clock1";
defparam ram_block3a38.port_b_data_out_clear = "none";
defparam ram_block3a38.port_b_data_out_clock = "none";
defparam ram_block3a38.port_b_data_width = 1;
defparam ram_block3a38.port_b_first_address = 0;
defparam ram_block3a38.port_b_first_bit_number = 6;
defparam ram_block3a38.port_b_last_address = 8191;
defparam ram_block3a38.port_b_logical_ram_depth = 16384;
defparam ram_block3a38.port_b_logical_ram_width = 32;
defparam ram_block3a38.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block3a38.port_b_read_enable_clock = "clock1";
defparam ram_block3a38.port_b_write_enable_clock = "clock1";
defparam ram_block3a38.ram_block_type = "M9K";
defparam ram_block3a38.mem_init3 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a38.mem_init2 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a38.mem_init1 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a38.mem_init0 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
// synopsys translate_on

// Location: M9K_X37_Y29_N0
cycloneive_ram_block ram_block3a6(
	.portawe(\decode4|eq_node[0]~1_combout ),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(\decode5|eq_node[0]~1_combout ),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock1),
	.ena0(ramaddr),
	.ena1(!ram_rom_addr_reg_13),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({data_a[6]}),
	.portaaddr({address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain({data_b[6]}),
	.portbaddr({address_b[12],address_b[11],address_b[10],address_b[9],address_b[8],address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.devclrn(devclrn),
	.devpor(devpor),
	.portadataout(ram_block3a6_PORTADATAOUT_bus),
	.portbdataout(ram_block3a6_PORTBDATAOUT_bus));
// synopsys translate_off
defparam ram_block3a6.clk0_core_clock_enable = "ena0";
defparam ram_block3a6.clk1_core_clock_enable = "ena1";
defparam ram_block3a6.data_interleave_offset_in_bits = 1;
defparam ram_block3a6.data_interleave_width_in_bits = 1;
defparam ram_block3a6.init_file = "meminit.hex";
defparam ram_block3a6.init_file_layout = "port_a";
defparam ram_block3a6.logical_ram_name = "ram:RAM|altsyncram:altsyncram_component|altsyncram_99f1:auto_generated|altsyncram_fta2:altsyncram1|ALTSYNCRAM";
defparam ram_block3a6.mixed_port_feed_through_mode = "dont_care";
defparam ram_block3a6.operation_mode = "bidir_dual_port";
defparam ram_block3a6.port_a_address_clear = "none";
defparam ram_block3a6.port_a_address_width = 13;
defparam ram_block3a6.port_a_byte_enable_clock = "none";
defparam ram_block3a6.port_a_data_out_clear = "none";
defparam ram_block3a6.port_a_data_out_clock = "none";
defparam ram_block3a6.port_a_data_width = 1;
defparam ram_block3a6.port_a_first_address = 0;
defparam ram_block3a6.port_a_first_bit_number = 6;
defparam ram_block3a6.port_a_last_address = 8191;
defparam ram_block3a6.port_a_logical_ram_depth = 16384;
defparam ram_block3a6.port_a_logical_ram_width = 32;
defparam ram_block3a6.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block3a6.port_b_address_clear = "none";
defparam ram_block3a6.port_b_address_clock = "clock1";
defparam ram_block3a6.port_b_address_width = 13;
defparam ram_block3a6.port_b_data_in_clock = "clock1";
defparam ram_block3a6.port_b_data_out_clear = "none";
defparam ram_block3a6.port_b_data_out_clock = "none";
defparam ram_block3a6.port_b_data_width = 1;
defparam ram_block3a6.port_b_first_address = 0;
defparam ram_block3a6.port_b_first_bit_number = 6;
defparam ram_block3a6.port_b_last_address = 8191;
defparam ram_block3a6.port_b_logical_ram_depth = 16384;
defparam ram_block3a6.port_b_logical_ram_width = 32;
defparam ram_block3a6.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block3a6.port_b_read_enable_clock = "clock1";
defparam ram_block3a6.port_b_write_enable_clock = "clock1";
defparam ram_block3a6.ram_block_type = "M9K";
defparam ram_block3a6.mem_init3 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a6.mem_init2 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a6.mem_init1 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a6.mem_init0 = 2048'h0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001003088D801A0F827000000000000000000000000000012042100402202200113;
// synopsys translate_on

// Location: M9K_X51_Y32_N0
cycloneive_ram_block ram_block3a39(
	.portawe(\decode4|eq_node[1]~0_combout ),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(\decode5|eq_node[1]~0_combout ),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock1),
	.ena0(!ramaddr),
	.ena1(ram_rom_addr_reg_13),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({data_a[7]}),
	.portaaddr({address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain({data_b[7]}),
	.portbaddr({address_b[12],address_b[11],address_b[10],address_b[9],address_b[8],address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.devclrn(devclrn),
	.devpor(devpor),
	.portadataout(ram_block3a39_PORTADATAOUT_bus),
	.portbdataout(ram_block3a39_PORTBDATAOUT_bus));
// synopsys translate_off
defparam ram_block3a39.clk0_core_clock_enable = "ena0";
defparam ram_block3a39.clk1_core_clock_enable = "ena1";
defparam ram_block3a39.data_interleave_offset_in_bits = 1;
defparam ram_block3a39.data_interleave_width_in_bits = 1;
defparam ram_block3a39.init_file = "meminit.hex";
defparam ram_block3a39.init_file_layout = "port_a";
defparam ram_block3a39.logical_ram_name = "ram:RAM|altsyncram:altsyncram_component|altsyncram_99f1:auto_generated|altsyncram_fta2:altsyncram1|ALTSYNCRAM";
defparam ram_block3a39.mixed_port_feed_through_mode = "dont_care";
defparam ram_block3a39.operation_mode = "bidir_dual_port";
defparam ram_block3a39.port_a_address_clear = "none";
defparam ram_block3a39.port_a_address_width = 13;
defparam ram_block3a39.port_a_byte_enable_clock = "none";
defparam ram_block3a39.port_a_data_out_clear = "none";
defparam ram_block3a39.port_a_data_out_clock = "none";
defparam ram_block3a39.port_a_data_width = 1;
defparam ram_block3a39.port_a_first_address = 0;
defparam ram_block3a39.port_a_first_bit_number = 7;
defparam ram_block3a39.port_a_last_address = 8191;
defparam ram_block3a39.port_a_logical_ram_depth = 16384;
defparam ram_block3a39.port_a_logical_ram_width = 32;
defparam ram_block3a39.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block3a39.port_b_address_clear = "none";
defparam ram_block3a39.port_b_address_clock = "clock1";
defparam ram_block3a39.port_b_address_width = 13;
defparam ram_block3a39.port_b_data_in_clock = "clock1";
defparam ram_block3a39.port_b_data_out_clear = "none";
defparam ram_block3a39.port_b_data_out_clock = "none";
defparam ram_block3a39.port_b_data_width = 1;
defparam ram_block3a39.port_b_first_address = 0;
defparam ram_block3a39.port_b_first_bit_number = 7;
defparam ram_block3a39.port_b_last_address = 8191;
defparam ram_block3a39.port_b_logical_ram_depth = 16384;
defparam ram_block3a39.port_b_logical_ram_width = 32;
defparam ram_block3a39.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block3a39.port_b_read_enable_clock = "clock1";
defparam ram_block3a39.port_b_write_enable_clock = "clock1";
defparam ram_block3a39.ram_block_type = "M9K";
defparam ram_block3a39.mem_init3 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a39.mem_init2 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a39.mem_init1 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a39.mem_init0 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
// synopsys translate_on

// Location: M9K_X37_Y28_N0
cycloneive_ram_block ram_block3a7(
	.portawe(\decode4|eq_node[0]~1_combout ),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(\decode5|eq_node[0]~1_combout ),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock1),
	.ena0(ramaddr),
	.ena1(!ram_rom_addr_reg_13),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({data_a[7]}),
	.portaaddr({address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain({data_b[7]}),
	.portbaddr({address_b[12],address_b[11],address_b[10],address_b[9],address_b[8],address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.devclrn(devclrn),
	.devpor(devpor),
	.portadataout(ram_block3a7_PORTADATAOUT_bus),
	.portbdataout(ram_block3a7_PORTBDATAOUT_bus));
// synopsys translate_off
defparam ram_block3a7.clk0_core_clock_enable = "ena0";
defparam ram_block3a7.clk1_core_clock_enable = "ena1";
defparam ram_block3a7.data_interleave_offset_in_bits = 1;
defparam ram_block3a7.data_interleave_width_in_bits = 1;
defparam ram_block3a7.init_file = "meminit.hex";
defparam ram_block3a7.init_file_layout = "port_a";
defparam ram_block3a7.logical_ram_name = "ram:RAM|altsyncram:altsyncram_component|altsyncram_99f1:auto_generated|altsyncram_fta2:altsyncram1|ALTSYNCRAM";
defparam ram_block3a7.mixed_port_feed_through_mode = "dont_care";
defparam ram_block3a7.operation_mode = "bidir_dual_port";
defparam ram_block3a7.port_a_address_clear = "none";
defparam ram_block3a7.port_a_address_width = 13;
defparam ram_block3a7.port_a_byte_enable_clock = "none";
defparam ram_block3a7.port_a_data_out_clear = "none";
defparam ram_block3a7.port_a_data_out_clock = "none";
defparam ram_block3a7.port_a_data_width = 1;
defparam ram_block3a7.port_a_first_address = 0;
defparam ram_block3a7.port_a_first_bit_number = 7;
defparam ram_block3a7.port_a_last_address = 8191;
defparam ram_block3a7.port_a_logical_ram_depth = 16384;
defparam ram_block3a7.port_a_logical_ram_width = 32;
defparam ram_block3a7.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block3a7.port_b_address_clear = "none";
defparam ram_block3a7.port_b_address_clock = "clock1";
defparam ram_block3a7.port_b_address_width = 13;
defparam ram_block3a7.port_b_data_in_clock = "clock1";
defparam ram_block3a7.port_b_data_out_clear = "none";
defparam ram_block3a7.port_b_data_out_clock = "none";
defparam ram_block3a7.port_b_data_width = 1;
defparam ram_block3a7.port_b_first_address = 0;
defparam ram_block3a7.port_b_first_bit_number = 7;
defparam ram_block3a7.port_b_last_address = 8191;
defparam ram_block3a7.port_b_logical_ram_depth = 16384;
defparam ram_block3a7.port_b_logical_ram_width = 32;
defparam ram_block3a7.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block3a7.port_b_read_enable_clock = "clock1";
defparam ram_block3a7.port_b_write_enable_clock = "clock1";
defparam ram_block3a7.ram_block_type = "M9K";
defparam ram_block3a7.mem_init3 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a7.mem_init2 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a7.mem_init1 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a7.mem_init0 = 2048'h0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000204210000220A200403;
// synopsys translate_on

// Location: M9K_X37_Y23_N0
cycloneive_ram_block ram_block3a40(
	.portawe(\decode4|eq_node[1]~0_combout ),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(\decode5|eq_node[1]~0_combout ),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock1),
	.ena0(!ramaddr),
	.ena1(ram_rom_addr_reg_13),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({data_a[8]}),
	.portaaddr({address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain({data_b[8]}),
	.portbaddr({address_b[12],address_b[11],address_b[10],address_b[9],address_b[8],address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.devclrn(devclrn),
	.devpor(devpor),
	.portadataout(ram_block3a40_PORTADATAOUT_bus),
	.portbdataout(ram_block3a40_PORTBDATAOUT_bus));
// synopsys translate_off
defparam ram_block3a40.clk0_core_clock_enable = "ena0";
defparam ram_block3a40.clk1_core_clock_enable = "ena1";
defparam ram_block3a40.data_interleave_offset_in_bits = 1;
defparam ram_block3a40.data_interleave_width_in_bits = 1;
defparam ram_block3a40.init_file = "meminit.hex";
defparam ram_block3a40.init_file_layout = "port_a";
defparam ram_block3a40.logical_ram_name = "ram:RAM|altsyncram:altsyncram_component|altsyncram_99f1:auto_generated|altsyncram_fta2:altsyncram1|ALTSYNCRAM";
defparam ram_block3a40.mixed_port_feed_through_mode = "dont_care";
defparam ram_block3a40.operation_mode = "bidir_dual_port";
defparam ram_block3a40.port_a_address_clear = "none";
defparam ram_block3a40.port_a_address_width = 13;
defparam ram_block3a40.port_a_byte_enable_clock = "none";
defparam ram_block3a40.port_a_data_out_clear = "none";
defparam ram_block3a40.port_a_data_out_clock = "none";
defparam ram_block3a40.port_a_data_width = 1;
defparam ram_block3a40.port_a_first_address = 0;
defparam ram_block3a40.port_a_first_bit_number = 8;
defparam ram_block3a40.port_a_last_address = 8191;
defparam ram_block3a40.port_a_logical_ram_depth = 16384;
defparam ram_block3a40.port_a_logical_ram_width = 32;
defparam ram_block3a40.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block3a40.port_b_address_clear = "none";
defparam ram_block3a40.port_b_address_clock = "clock1";
defparam ram_block3a40.port_b_address_width = 13;
defparam ram_block3a40.port_b_data_in_clock = "clock1";
defparam ram_block3a40.port_b_data_out_clear = "none";
defparam ram_block3a40.port_b_data_out_clock = "none";
defparam ram_block3a40.port_b_data_width = 1;
defparam ram_block3a40.port_b_first_address = 0;
defparam ram_block3a40.port_b_first_bit_number = 8;
defparam ram_block3a40.port_b_last_address = 8191;
defparam ram_block3a40.port_b_logical_ram_depth = 16384;
defparam ram_block3a40.port_b_logical_ram_width = 32;
defparam ram_block3a40.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block3a40.port_b_read_enable_clock = "clock1";
defparam ram_block3a40.port_b_write_enable_clock = "clock1";
defparam ram_block3a40.ram_block_type = "M9K";
defparam ram_block3a40.mem_init3 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a40.mem_init2 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a40.mem_init1 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a40.mem_init0 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
// synopsys translate_on

// Location: M9K_X37_Y26_N0
cycloneive_ram_block ram_block3a8(
	.portawe(\decode4|eq_node[0]~1_combout ),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(\decode5|eq_node[0]~1_combout ),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock1),
	.ena0(ramaddr),
	.ena1(!ram_rom_addr_reg_13),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({data_a[8]}),
	.portaaddr({address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain({data_b[8]}),
	.portbaddr({address_b[12],address_b[11],address_b[10],address_b[9],address_b[8],address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.devclrn(devclrn),
	.devpor(devpor),
	.portadataout(ram_block3a8_PORTADATAOUT_bus),
	.portbdataout(ram_block3a8_PORTBDATAOUT_bus));
// synopsys translate_off
defparam ram_block3a8.clk0_core_clock_enable = "ena0";
defparam ram_block3a8.clk1_core_clock_enable = "ena1";
defparam ram_block3a8.data_interleave_offset_in_bits = 1;
defparam ram_block3a8.data_interleave_width_in_bits = 1;
defparam ram_block3a8.init_file = "meminit.hex";
defparam ram_block3a8.init_file_layout = "port_a";
defparam ram_block3a8.logical_ram_name = "ram:RAM|altsyncram:altsyncram_component|altsyncram_99f1:auto_generated|altsyncram_fta2:altsyncram1|ALTSYNCRAM";
defparam ram_block3a8.mixed_port_feed_through_mode = "dont_care";
defparam ram_block3a8.operation_mode = "bidir_dual_port";
defparam ram_block3a8.port_a_address_clear = "none";
defparam ram_block3a8.port_a_address_width = 13;
defparam ram_block3a8.port_a_byte_enable_clock = "none";
defparam ram_block3a8.port_a_data_out_clear = "none";
defparam ram_block3a8.port_a_data_out_clock = "none";
defparam ram_block3a8.port_a_data_width = 1;
defparam ram_block3a8.port_a_first_address = 0;
defparam ram_block3a8.port_a_first_bit_number = 8;
defparam ram_block3a8.port_a_last_address = 8191;
defparam ram_block3a8.port_a_logical_ram_depth = 16384;
defparam ram_block3a8.port_a_logical_ram_width = 32;
defparam ram_block3a8.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block3a8.port_b_address_clear = "none";
defparam ram_block3a8.port_b_address_clock = "clock1";
defparam ram_block3a8.port_b_address_width = 13;
defparam ram_block3a8.port_b_data_in_clock = "clock1";
defparam ram_block3a8.port_b_data_out_clear = "none";
defparam ram_block3a8.port_b_data_out_clock = "none";
defparam ram_block3a8.port_b_data_width = 1;
defparam ram_block3a8.port_b_first_address = 0;
defparam ram_block3a8.port_b_first_bit_number = 8;
defparam ram_block3a8.port_b_last_address = 8191;
defparam ram_block3a8.port_b_logical_ram_depth = 16384;
defparam ram_block3a8.port_b_logical_ram_width = 32;
defparam ram_block3a8.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block3a8.port_b_read_enable_clock = "clock1";
defparam ram_block3a8.port_b_write_enable_clock = "clock1";
defparam ram_block3a8.ram_block_type = "M9K";
defparam ram_block3a8.mem_init3 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a8.mem_init2 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a8.mem_init1 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a8.mem_init0 = 2048'h0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000204210000220220080F;
// synopsys translate_on

// Location: M9K_X37_Y35_N0
cycloneive_ram_block ram_block3a41(
	.portawe(\decode4|eq_node[1]~0_combout ),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(\decode5|eq_node[1]~0_combout ),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock1),
	.ena0(!ramaddr),
	.ena1(ram_rom_addr_reg_13),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({data_a[9]}),
	.portaaddr({address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain({data_b[9]}),
	.portbaddr({address_b[12],address_b[11],address_b[10],address_b[9],address_b[8],address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.devclrn(devclrn),
	.devpor(devpor),
	.portadataout(ram_block3a41_PORTADATAOUT_bus),
	.portbdataout(ram_block3a41_PORTBDATAOUT_bus));
// synopsys translate_off
defparam ram_block3a41.clk0_core_clock_enable = "ena0";
defparam ram_block3a41.clk1_core_clock_enable = "ena1";
defparam ram_block3a41.data_interleave_offset_in_bits = 1;
defparam ram_block3a41.data_interleave_width_in_bits = 1;
defparam ram_block3a41.init_file = "meminit.hex";
defparam ram_block3a41.init_file_layout = "port_a";
defparam ram_block3a41.logical_ram_name = "ram:RAM|altsyncram:altsyncram_component|altsyncram_99f1:auto_generated|altsyncram_fta2:altsyncram1|ALTSYNCRAM";
defparam ram_block3a41.mixed_port_feed_through_mode = "dont_care";
defparam ram_block3a41.operation_mode = "bidir_dual_port";
defparam ram_block3a41.port_a_address_clear = "none";
defparam ram_block3a41.port_a_address_width = 13;
defparam ram_block3a41.port_a_byte_enable_clock = "none";
defparam ram_block3a41.port_a_data_out_clear = "none";
defparam ram_block3a41.port_a_data_out_clock = "none";
defparam ram_block3a41.port_a_data_width = 1;
defparam ram_block3a41.port_a_first_address = 0;
defparam ram_block3a41.port_a_first_bit_number = 9;
defparam ram_block3a41.port_a_last_address = 8191;
defparam ram_block3a41.port_a_logical_ram_depth = 16384;
defparam ram_block3a41.port_a_logical_ram_width = 32;
defparam ram_block3a41.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block3a41.port_b_address_clear = "none";
defparam ram_block3a41.port_b_address_clock = "clock1";
defparam ram_block3a41.port_b_address_width = 13;
defparam ram_block3a41.port_b_data_in_clock = "clock1";
defparam ram_block3a41.port_b_data_out_clear = "none";
defparam ram_block3a41.port_b_data_out_clock = "none";
defparam ram_block3a41.port_b_data_width = 1;
defparam ram_block3a41.port_b_first_address = 0;
defparam ram_block3a41.port_b_first_bit_number = 9;
defparam ram_block3a41.port_b_last_address = 8191;
defparam ram_block3a41.port_b_logical_ram_depth = 16384;
defparam ram_block3a41.port_b_logical_ram_width = 32;
defparam ram_block3a41.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block3a41.port_b_read_enable_clock = "clock1";
defparam ram_block3a41.port_b_write_enable_clock = "clock1";
defparam ram_block3a41.ram_block_type = "M9K";
defparam ram_block3a41.mem_init3 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a41.mem_init2 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a41.mem_init1 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a41.mem_init0 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
// synopsys translate_on

// Location: M9K_X37_Y38_N0
cycloneive_ram_block ram_block3a9(
	.portawe(\decode4|eq_node[0]~1_combout ),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(\decode5|eq_node[0]~1_combout ),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock1),
	.ena0(ramaddr),
	.ena1(!ram_rom_addr_reg_13),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({data_a[9]}),
	.portaaddr({address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain({data_b[9]}),
	.portbaddr({address_b[12],address_b[11],address_b[10],address_b[9],address_b[8],address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.devclrn(devclrn),
	.devpor(devpor),
	.portadataout(ram_block3a9_PORTADATAOUT_bus),
	.portbdataout(ram_block3a9_PORTBDATAOUT_bus));
// synopsys translate_off
defparam ram_block3a9.clk0_core_clock_enable = "ena0";
defparam ram_block3a9.clk1_core_clock_enable = "ena1";
defparam ram_block3a9.data_interleave_offset_in_bits = 1;
defparam ram_block3a9.data_interleave_width_in_bits = 1;
defparam ram_block3a9.init_file = "meminit.hex";
defparam ram_block3a9.init_file_layout = "port_a";
defparam ram_block3a9.logical_ram_name = "ram:RAM|altsyncram:altsyncram_component|altsyncram_99f1:auto_generated|altsyncram_fta2:altsyncram1|ALTSYNCRAM";
defparam ram_block3a9.mixed_port_feed_through_mode = "dont_care";
defparam ram_block3a9.operation_mode = "bidir_dual_port";
defparam ram_block3a9.port_a_address_clear = "none";
defparam ram_block3a9.port_a_address_width = 13;
defparam ram_block3a9.port_a_byte_enable_clock = "none";
defparam ram_block3a9.port_a_data_out_clear = "none";
defparam ram_block3a9.port_a_data_out_clock = "none";
defparam ram_block3a9.port_a_data_width = 1;
defparam ram_block3a9.port_a_first_address = 0;
defparam ram_block3a9.port_a_first_bit_number = 9;
defparam ram_block3a9.port_a_last_address = 8191;
defparam ram_block3a9.port_a_logical_ram_depth = 16384;
defparam ram_block3a9.port_a_logical_ram_width = 32;
defparam ram_block3a9.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block3a9.port_b_address_clear = "none";
defparam ram_block3a9.port_b_address_clock = "clock1";
defparam ram_block3a9.port_b_address_width = 13;
defparam ram_block3a9.port_b_data_in_clock = "clock1";
defparam ram_block3a9.port_b_data_out_clear = "none";
defparam ram_block3a9.port_b_data_out_clock = "none";
defparam ram_block3a9.port_b_data_width = 1;
defparam ram_block3a9.port_b_first_address = 0;
defparam ram_block3a9.port_b_first_bit_number = 9;
defparam ram_block3a9.port_b_last_address = 8191;
defparam ram_block3a9.port_b_logical_ram_depth = 16384;
defparam ram_block3a9.port_b_logical_ram_width = 32;
defparam ram_block3a9.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block3a9.port_b_read_enable_clock = "clock1";
defparam ram_block3a9.port_b_write_enable_clock = "clock1";
defparam ram_block3a9.ram_block_type = "M9K";
defparam ram_block3a9.mem_init3 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a9.mem_init2 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a9.mem_init1 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a9.mem_init0 = 2048'h0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000204210000220220080F;
// synopsys translate_on

// Location: M9K_X37_Y34_N0
cycloneive_ram_block ram_block3a42(
	.portawe(\decode4|eq_node[1]~0_combout ),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(\decode5|eq_node[1]~0_combout ),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock1),
	.ena0(!ramaddr),
	.ena1(ram_rom_addr_reg_13),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({data_a[10]}),
	.portaaddr({address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain({data_b[10]}),
	.portbaddr({address_b[12],address_b[11],address_b[10],address_b[9],address_b[8],address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.devclrn(devclrn),
	.devpor(devpor),
	.portadataout(ram_block3a42_PORTADATAOUT_bus),
	.portbdataout(ram_block3a42_PORTBDATAOUT_bus));
// synopsys translate_off
defparam ram_block3a42.clk0_core_clock_enable = "ena0";
defparam ram_block3a42.clk1_core_clock_enable = "ena1";
defparam ram_block3a42.data_interleave_offset_in_bits = 1;
defparam ram_block3a42.data_interleave_width_in_bits = 1;
defparam ram_block3a42.init_file = "meminit.hex";
defparam ram_block3a42.init_file_layout = "port_a";
defparam ram_block3a42.logical_ram_name = "ram:RAM|altsyncram:altsyncram_component|altsyncram_99f1:auto_generated|altsyncram_fta2:altsyncram1|ALTSYNCRAM";
defparam ram_block3a42.mixed_port_feed_through_mode = "dont_care";
defparam ram_block3a42.operation_mode = "bidir_dual_port";
defparam ram_block3a42.port_a_address_clear = "none";
defparam ram_block3a42.port_a_address_width = 13;
defparam ram_block3a42.port_a_byte_enable_clock = "none";
defparam ram_block3a42.port_a_data_out_clear = "none";
defparam ram_block3a42.port_a_data_out_clock = "none";
defparam ram_block3a42.port_a_data_width = 1;
defparam ram_block3a42.port_a_first_address = 0;
defparam ram_block3a42.port_a_first_bit_number = 10;
defparam ram_block3a42.port_a_last_address = 8191;
defparam ram_block3a42.port_a_logical_ram_depth = 16384;
defparam ram_block3a42.port_a_logical_ram_width = 32;
defparam ram_block3a42.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block3a42.port_b_address_clear = "none";
defparam ram_block3a42.port_b_address_clock = "clock1";
defparam ram_block3a42.port_b_address_width = 13;
defparam ram_block3a42.port_b_data_in_clock = "clock1";
defparam ram_block3a42.port_b_data_out_clear = "none";
defparam ram_block3a42.port_b_data_out_clock = "none";
defparam ram_block3a42.port_b_data_width = 1;
defparam ram_block3a42.port_b_first_address = 0;
defparam ram_block3a42.port_b_first_bit_number = 10;
defparam ram_block3a42.port_b_last_address = 8191;
defparam ram_block3a42.port_b_logical_ram_depth = 16384;
defparam ram_block3a42.port_b_logical_ram_width = 32;
defparam ram_block3a42.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block3a42.port_b_read_enable_clock = "clock1";
defparam ram_block3a42.port_b_write_enable_clock = "clock1";
defparam ram_block3a42.ram_block_type = "M9K";
defparam ram_block3a42.mem_init3 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a42.mem_init2 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a42.mem_init1 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a42.mem_init0 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
// synopsys translate_on

// Location: M9K_X37_Y32_N0
cycloneive_ram_block ram_block3a10(
	.portawe(\decode4|eq_node[0]~1_combout ),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(\decode5|eq_node[0]~1_combout ),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock1),
	.ena0(ramaddr),
	.ena1(!ram_rom_addr_reg_13),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({data_a[10]}),
	.portaaddr({address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain({data_b[10]}),
	.portbaddr({address_b[12],address_b[11],address_b[10],address_b[9],address_b[8],address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.devclrn(devclrn),
	.devpor(devpor),
	.portadataout(ram_block3a10_PORTADATAOUT_bus),
	.portbdataout(ram_block3a10_PORTBDATAOUT_bus));
// synopsys translate_off
defparam ram_block3a10.clk0_core_clock_enable = "ena0";
defparam ram_block3a10.clk1_core_clock_enable = "ena1";
defparam ram_block3a10.data_interleave_offset_in_bits = 1;
defparam ram_block3a10.data_interleave_width_in_bits = 1;
defparam ram_block3a10.init_file = "meminit.hex";
defparam ram_block3a10.init_file_layout = "port_a";
defparam ram_block3a10.logical_ram_name = "ram:RAM|altsyncram:altsyncram_component|altsyncram_99f1:auto_generated|altsyncram_fta2:altsyncram1|ALTSYNCRAM";
defparam ram_block3a10.mixed_port_feed_through_mode = "dont_care";
defparam ram_block3a10.operation_mode = "bidir_dual_port";
defparam ram_block3a10.port_a_address_clear = "none";
defparam ram_block3a10.port_a_address_width = 13;
defparam ram_block3a10.port_a_byte_enable_clock = "none";
defparam ram_block3a10.port_a_data_out_clear = "none";
defparam ram_block3a10.port_a_data_out_clock = "none";
defparam ram_block3a10.port_a_data_width = 1;
defparam ram_block3a10.port_a_first_address = 0;
defparam ram_block3a10.port_a_first_bit_number = 10;
defparam ram_block3a10.port_a_last_address = 8191;
defparam ram_block3a10.port_a_logical_ram_depth = 16384;
defparam ram_block3a10.port_a_logical_ram_width = 32;
defparam ram_block3a10.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block3a10.port_b_address_clear = "none";
defparam ram_block3a10.port_b_address_clock = "clock1";
defparam ram_block3a10.port_b_address_width = 13;
defparam ram_block3a10.port_b_data_in_clock = "clock1";
defparam ram_block3a10.port_b_data_out_clear = "none";
defparam ram_block3a10.port_b_data_out_clock = "none";
defparam ram_block3a10.port_b_data_width = 1;
defparam ram_block3a10.port_b_first_address = 0;
defparam ram_block3a10.port_b_first_bit_number = 10;
defparam ram_block3a10.port_b_last_address = 8191;
defparam ram_block3a10.port_b_logical_ram_depth = 16384;
defparam ram_block3a10.port_b_logical_ram_width = 32;
defparam ram_block3a10.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block3a10.port_b_read_enable_clock = "clock1";
defparam ram_block3a10.port_b_write_enable_clock = "clock1";
defparam ram_block3a10.ram_block_type = "M9K";
defparam ram_block3a10.mem_init3 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a10.mem_init2 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a10.mem_init1 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a10.mem_init0 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000002042100002202300003;
// synopsys translate_on

// Location: M9K_X64_Y29_N0
cycloneive_ram_block ram_block3a43(
	.portawe(\decode4|eq_node[1]~0_combout ),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(\decode5|eq_node[1]~0_combout ),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock1),
	.ena0(!ramaddr),
	.ena1(ram_rom_addr_reg_13),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({data_a[11]}),
	.portaaddr({address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain({data_b[11]}),
	.portbaddr({address_b[12],address_b[11],address_b[10],address_b[9],address_b[8],address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.devclrn(devclrn),
	.devpor(devpor),
	.portadataout(ram_block3a43_PORTADATAOUT_bus),
	.portbdataout(ram_block3a43_PORTBDATAOUT_bus));
// synopsys translate_off
defparam ram_block3a43.clk0_core_clock_enable = "ena0";
defparam ram_block3a43.clk1_core_clock_enable = "ena1";
defparam ram_block3a43.data_interleave_offset_in_bits = 1;
defparam ram_block3a43.data_interleave_width_in_bits = 1;
defparam ram_block3a43.init_file = "meminit.hex";
defparam ram_block3a43.init_file_layout = "port_a";
defparam ram_block3a43.logical_ram_name = "ram:RAM|altsyncram:altsyncram_component|altsyncram_99f1:auto_generated|altsyncram_fta2:altsyncram1|ALTSYNCRAM";
defparam ram_block3a43.mixed_port_feed_through_mode = "dont_care";
defparam ram_block3a43.operation_mode = "bidir_dual_port";
defparam ram_block3a43.port_a_address_clear = "none";
defparam ram_block3a43.port_a_address_width = 13;
defparam ram_block3a43.port_a_byte_enable_clock = "none";
defparam ram_block3a43.port_a_data_out_clear = "none";
defparam ram_block3a43.port_a_data_out_clock = "none";
defparam ram_block3a43.port_a_data_width = 1;
defparam ram_block3a43.port_a_first_address = 0;
defparam ram_block3a43.port_a_first_bit_number = 11;
defparam ram_block3a43.port_a_last_address = 8191;
defparam ram_block3a43.port_a_logical_ram_depth = 16384;
defparam ram_block3a43.port_a_logical_ram_width = 32;
defparam ram_block3a43.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block3a43.port_b_address_clear = "none";
defparam ram_block3a43.port_b_address_clock = "clock1";
defparam ram_block3a43.port_b_address_width = 13;
defparam ram_block3a43.port_b_data_in_clock = "clock1";
defparam ram_block3a43.port_b_data_out_clear = "none";
defparam ram_block3a43.port_b_data_out_clock = "none";
defparam ram_block3a43.port_b_data_width = 1;
defparam ram_block3a43.port_b_first_address = 0;
defparam ram_block3a43.port_b_first_bit_number = 11;
defparam ram_block3a43.port_b_last_address = 8191;
defparam ram_block3a43.port_b_logical_ram_depth = 16384;
defparam ram_block3a43.port_b_logical_ram_width = 32;
defparam ram_block3a43.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block3a43.port_b_read_enable_clock = "clock1";
defparam ram_block3a43.port_b_write_enable_clock = "clock1";
defparam ram_block3a43.ram_block_type = "M9K";
defparam ram_block3a43.mem_init3 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a43.mem_init2 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a43.mem_init1 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a43.mem_init0 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
// synopsys translate_on

// Location: M9K_X64_Y27_N0
cycloneive_ram_block ram_block3a11(
	.portawe(\decode4|eq_node[0]~1_combout ),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(\decode5|eq_node[0]~1_combout ),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock1),
	.ena0(ramaddr),
	.ena1(!ram_rom_addr_reg_13),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({data_a[11]}),
	.portaaddr({address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain({data_b[11]}),
	.portbaddr({address_b[12],address_b[11],address_b[10],address_b[9],address_b[8],address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.devclrn(devclrn),
	.devpor(devpor),
	.portadataout(ram_block3a11_PORTADATAOUT_bus),
	.portbdataout(ram_block3a11_PORTBDATAOUT_bus));
// synopsys translate_off
defparam ram_block3a11.clk0_core_clock_enable = "ena0";
defparam ram_block3a11.clk1_core_clock_enable = "ena1";
defparam ram_block3a11.data_interleave_offset_in_bits = 1;
defparam ram_block3a11.data_interleave_width_in_bits = 1;
defparam ram_block3a11.init_file = "meminit.hex";
defparam ram_block3a11.init_file_layout = "port_a";
defparam ram_block3a11.logical_ram_name = "ram:RAM|altsyncram:altsyncram_component|altsyncram_99f1:auto_generated|altsyncram_fta2:altsyncram1|ALTSYNCRAM";
defparam ram_block3a11.mixed_port_feed_through_mode = "dont_care";
defparam ram_block3a11.operation_mode = "bidir_dual_port";
defparam ram_block3a11.port_a_address_clear = "none";
defparam ram_block3a11.port_a_address_width = 13;
defparam ram_block3a11.port_a_byte_enable_clock = "none";
defparam ram_block3a11.port_a_data_out_clear = "none";
defparam ram_block3a11.port_a_data_out_clock = "none";
defparam ram_block3a11.port_a_data_width = 1;
defparam ram_block3a11.port_a_first_address = 0;
defparam ram_block3a11.port_a_first_bit_number = 11;
defparam ram_block3a11.port_a_last_address = 8191;
defparam ram_block3a11.port_a_logical_ram_depth = 16384;
defparam ram_block3a11.port_a_logical_ram_width = 32;
defparam ram_block3a11.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block3a11.port_b_address_clear = "none";
defparam ram_block3a11.port_b_address_clock = "clock1";
defparam ram_block3a11.port_b_address_width = 13;
defparam ram_block3a11.port_b_data_in_clock = "clock1";
defparam ram_block3a11.port_b_data_out_clear = "none";
defparam ram_block3a11.port_b_data_out_clock = "none";
defparam ram_block3a11.port_b_data_width = 1;
defparam ram_block3a11.port_b_first_address = 0;
defparam ram_block3a11.port_b_first_bit_number = 11;
defparam ram_block3a11.port_b_last_address = 8191;
defparam ram_block3a11.port_b_logical_ram_depth = 16384;
defparam ram_block3a11.port_b_logical_ram_width = 32;
defparam ram_block3a11.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block3a11.port_b_read_enable_clock = "clock1";
defparam ram_block3a11.port_b_write_enable_clock = "clock1";
defparam ram_block3a11.ram_block_type = "M9K";
defparam ram_block3a11.mem_init3 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a11.mem_init2 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a11.mem_init1 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a11.mem_init0 = 2048'h0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000204210800265A2A2233;
// synopsys translate_on

// Location: M9K_X51_Y35_N0
cycloneive_ram_block ram_block3a44(
	.portawe(\decode4|eq_node[1]~0_combout ),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(\decode5|eq_node[1]~0_combout ),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock1),
	.ena0(!ramaddr),
	.ena1(ram_rom_addr_reg_13),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({data_a[12]}),
	.portaaddr({address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain({data_b[12]}),
	.portbaddr({address_b[12],address_b[11],address_b[10],address_b[9],address_b[8],address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.devclrn(devclrn),
	.devpor(devpor),
	.portadataout(ram_block3a44_PORTADATAOUT_bus),
	.portbdataout(ram_block3a44_PORTBDATAOUT_bus));
// synopsys translate_off
defparam ram_block3a44.clk0_core_clock_enable = "ena0";
defparam ram_block3a44.clk1_core_clock_enable = "ena1";
defparam ram_block3a44.data_interleave_offset_in_bits = 1;
defparam ram_block3a44.data_interleave_width_in_bits = 1;
defparam ram_block3a44.init_file = "meminit.hex";
defparam ram_block3a44.init_file_layout = "port_a";
defparam ram_block3a44.logical_ram_name = "ram:RAM|altsyncram:altsyncram_component|altsyncram_99f1:auto_generated|altsyncram_fta2:altsyncram1|ALTSYNCRAM";
defparam ram_block3a44.mixed_port_feed_through_mode = "dont_care";
defparam ram_block3a44.operation_mode = "bidir_dual_port";
defparam ram_block3a44.port_a_address_clear = "none";
defparam ram_block3a44.port_a_address_width = 13;
defparam ram_block3a44.port_a_byte_enable_clock = "none";
defparam ram_block3a44.port_a_data_out_clear = "none";
defparam ram_block3a44.port_a_data_out_clock = "none";
defparam ram_block3a44.port_a_data_width = 1;
defparam ram_block3a44.port_a_first_address = 0;
defparam ram_block3a44.port_a_first_bit_number = 12;
defparam ram_block3a44.port_a_last_address = 8191;
defparam ram_block3a44.port_a_logical_ram_depth = 16384;
defparam ram_block3a44.port_a_logical_ram_width = 32;
defparam ram_block3a44.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block3a44.port_b_address_clear = "none";
defparam ram_block3a44.port_b_address_clock = "clock1";
defparam ram_block3a44.port_b_address_width = 13;
defparam ram_block3a44.port_b_data_in_clock = "clock1";
defparam ram_block3a44.port_b_data_out_clear = "none";
defparam ram_block3a44.port_b_data_out_clock = "none";
defparam ram_block3a44.port_b_data_width = 1;
defparam ram_block3a44.port_b_first_address = 0;
defparam ram_block3a44.port_b_first_bit_number = 12;
defparam ram_block3a44.port_b_last_address = 8191;
defparam ram_block3a44.port_b_logical_ram_depth = 16384;
defparam ram_block3a44.port_b_logical_ram_width = 32;
defparam ram_block3a44.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block3a44.port_b_read_enable_clock = "clock1";
defparam ram_block3a44.port_b_write_enable_clock = "clock1";
defparam ram_block3a44.ram_block_type = "M9K";
defparam ram_block3a44.mem_init3 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a44.mem_init2 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a44.mem_init1 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a44.mem_init0 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
// synopsys translate_on

// Location: M9K_X64_Y38_N0
cycloneive_ram_block ram_block3a12(
	.portawe(\decode4|eq_node[0]~1_combout ),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(\decode5|eq_node[0]~1_combout ),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock1),
	.ena0(ramaddr),
	.ena1(!ram_rom_addr_reg_13),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({data_a[12]}),
	.portaaddr({address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain({data_b[12]}),
	.portbaddr({address_b[12],address_b[11],address_b[10],address_b[9],address_b[8],address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.devclrn(devclrn),
	.devpor(devpor),
	.portadataout(ram_block3a12_PORTADATAOUT_bus),
	.portbdataout(ram_block3a12_PORTBDATAOUT_bus));
// synopsys translate_off
defparam ram_block3a12.clk0_core_clock_enable = "ena0";
defparam ram_block3a12.clk1_core_clock_enable = "ena1";
defparam ram_block3a12.data_interleave_offset_in_bits = 1;
defparam ram_block3a12.data_interleave_width_in_bits = 1;
defparam ram_block3a12.init_file = "meminit.hex";
defparam ram_block3a12.init_file_layout = "port_a";
defparam ram_block3a12.logical_ram_name = "ram:RAM|altsyncram:altsyncram_component|altsyncram_99f1:auto_generated|altsyncram_fta2:altsyncram1|ALTSYNCRAM";
defparam ram_block3a12.mixed_port_feed_through_mode = "dont_care";
defparam ram_block3a12.operation_mode = "bidir_dual_port";
defparam ram_block3a12.port_a_address_clear = "none";
defparam ram_block3a12.port_a_address_width = 13;
defparam ram_block3a12.port_a_byte_enable_clock = "none";
defparam ram_block3a12.port_a_data_out_clear = "none";
defparam ram_block3a12.port_a_data_out_clock = "none";
defparam ram_block3a12.port_a_data_width = 1;
defparam ram_block3a12.port_a_first_address = 0;
defparam ram_block3a12.port_a_first_bit_number = 12;
defparam ram_block3a12.port_a_last_address = 8191;
defparam ram_block3a12.port_a_logical_ram_depth = 16384;
defparam ram_block3a12.port_a_logical_ram_width = 32;
defparam ram_block3a12.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block3a12.port_b_address_clear = "none";
defparam ram_block3a12.port_b_address_clock = "clock1";
defparam ram_block3a12.port_b_address_width = 13;
defparam ram_block3a12.port_b_data_in_clock = "clock1";
defparam ram_block3a12.port_b_data_out_clear = "none";
defparam ram_block3a12.port_b_data_out_clock = "none";
defparam ram_block3a12.port_b_data_width = 1;
defparam ram_block3a12.port_b_first_address = 0;
defparam ram_block3a12.port_b_first_bit_number = 12;
defparam ram_block3a12.port_b_last_address = 8191;
defparam ram_block3a12.port_b_logical_ram_depth = 16384;
defparam ram_block3a12.port_b_logical_ram_width = 32;
defparam ram_block3a12.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block3a12.port_b_read_enable_clock = "clock1";
defparam ram_block3a12.port_b_write_enable_clock = "clock1";
defparam ram_block3a12.ram_block_type = "M9K";
defparam ram_block3a12.mem_init3 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a12.mem_init2 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a12.mem_init1 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a12.mem_init0 = 2048'h000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000020421000022022C2043;
// synopsys translate_on

// Location: M9K_X37_Y36_N0
cycloneive_ram_block ram_block3a45(
	.portawe(\decode4|eq_node[1]~0_combout ),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(\decode5|eq_node[1]~0_combout ),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock1),
	.ena0(!ramaddr),
	.ena1(ram_rom_addr_reg_13),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({data_a[13]}),
	.portaaddr({address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain({data_b[13]}),
	.portbaddr({address_b[12],address_b[11],address_b[10],address_b[9],address_b[8],address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.devclrn(devclrn),
	.devpor(devpor),
	.portadataout(ram_block3a45_PORTADATAOUT_bus),
	.portbdataout(ram_block3a45_PORTBDATAOUT_bus));
// synopsys translate_off
defparam ram_block3a45.clk0_core_clock_enable = "ena0";
defparam ram_block3a45.clk1_core_clock_enable = "ena1";
defparam ram_block3a45.data_interleave_offset_in_bits = 1;
defparam ram_block3a45.data_interleave_width_in_bits = 1;
defparam ram_block3a45.init_file = "meminit.hex";
defparam ram_block3a45.init_file_layout = "port_a";
defparam ram_block3a45.logical_ram_name = "ram:RAM|altsyncram:altsyncram_component|altsyncram_99f1:auto_generated|altsyncram_fta2:altsyncram1|ALTSYNCRAM";
defparam ram_block3a45.mixed_port_feed_through_mode = "dont_care";
defparam ram_block3a45.operation_mode = "bidir_dual_port";
defparam ram_block3a45.port_a_address_clear = "none";
defparam ram_block3a45.port_a_address_width = 13;
defparam ram_block3a45.port_a_byte_enable_clock = "none";
defparam ram_block3a45.port_a_data_out_clear = "none";
defparam ram_block3a45.port_a_data_out_clock = "none";
defparam ram_block3a45.port_a_data_width = 1;
defparam ram_block3a45.port_a_first_address = 0;
defparam ram_block3a45.port_a_first_bit_number = 13;
defparam ram_block3a45.port_a_last_address = 8191;
defparam ram_block3a45.port_a_logical_ram_depth = 16384;
defparam ram_block3a45.port_a_logical_ram_width = 32;
defparam ram_block3a45.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block3a45.port_b_address_clear = "none";
defparam ram_block3a45.port_b_address_clock = "clock1";
defparam ram_block3a45.port_b_address_width = 13;
defparam ram_block3a45.port_b_data_in_clock = "clock1";
defparam ram_block3a45.port_b_data_out_clear = "none";
defparam ram_block3a45.port_b_data_out_clock = "none";
defparam ram_block3a45.port_b_data_width = 1;
defparam ram_block3a45.port_b_first_address = 0;
defparam ram_block3a45.port_b_first_bit_number = 13;
defparam ram_block3a45.port_b_last_address = 8191;
defparam ram_block3a45.port_b_logical_ram_depth = 16384;
defparam ram_block3a45.port_b_logical_ram_width = 32;
defparam ram_block3a45.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block3a45.port_b_read_enable_clock = "clock1";
defparam ram_block3a45.port_b_write_enable_clock = "clock1";
defparam ram_block3a45.ram_block_type = "M9K";
defparam ram_block3a45.mem_init3 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a45.mem_init2 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a45.mem_init1 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a45.mem_init0 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
// synopsys translate_on

// Location: M9K_X37_Y33_N0
cycloneive_ram_block ram_block3a13(
	.portawe(\decode4|eq_node[0]~1_combout ),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(\decode5|eq_node[0]~1_combout ),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock1),
	.ena0(ramaddr),
	.ena1(!ram_rom_addr_reg_13),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({data_a[13]}),
	.portaaddr({address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain({data_b[13]}),
	.portbaddr({address_b[12],address_b[11],address_b[10],address_b[9],address_b[8],address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.devclrn(devclrn),
	.devpor(devpor),
	.portadataout(ram_block3a13_PORTADATAOUT_bus),
	.portbdataout(ram_block3a13_PORTBDATAOUT_bus));
// synopsys translate_off
defparam ram_block3a13.clk0_core_clock_enable = "ena0";
defparam ram_block3a13.clk1_core_clock_enable = "ena1";
defparam ram_block3a13.data_interleave_offset_in_bits = 1;
defparam ram_block3a13.data_interleave_width_in_bits = 1;
defparam ram_block3a13.init_file = "meminit.hex";
defparam ram_block3a13.init_file_layout = "port_a";
defparam ram_block3a13.logical_ram_name = "ram:RAM|altsyncram:altsyncram_component|altsyncram_99f1:auto_generated|altsyncram_fta2:altsyncram1|ALTSYNCRAM";
defparam ram_block3a13.mixed_port_feed_through_mode = "dont_care";
defparam ram_block3a13.operation_mode = "bidir_dual_port";
defparam ram_block3a13.port_a_address_clear = "none";
defparam ram_block3a13.port_a_address_width = 13;
defparam ram_block3a13.port_a_byte_enable_clock = "none";
defparam ram_block3a13.port_a_data_out_clear = "none";
defparam ram_block3a13.port_a_data_out_clock = "none";
defparam ram_block3a13.port_a_data_width = 1;
defparam ram_block3a13.port_a_first_address = 0;
defparam ram_block3a13.port_a_first_bit_number = 13;
defparam ram_block3a13.port_a_last_address = 8191;
defparam ram_block3a13.port_a_logical_ram_depth = 16384;
defparam ram_block3a13.port_a_logical_ram_width = 32;
defparam ram_block3a13.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block3a13.port_b_address_clear = "none";
defparam ram_block3a13.port_b_address_clock = "clock1";
defparam ram_block3a13.port_b_address_width = 13;
defparam ram_block3a13.port_b_data_in_clock = "clock1";
defparam ram_block3a13.port_b_data_out_clear = "none";
defparam ram_block3a13.port_b_data_out_clock = "none";
defparam ram_block3a13.port_b_data_width = 1;
defparam ram_block3a13.port_b_first_address = 0;
defparam ram_block3a13.port_b_first_bit_number = 13;
defparam ram_block3a13.port_b_last_address = 8191;
defparam ram_block3a13.port_b_logical_ram_depth = 16384;
defparam ram_block3a13.port_b_logical_ram_width = 32;
defparam ram_block3a13.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block3a13.port_b_read_enable_clock = "clock1";
defparam ram_block3a13.port_b_write_enable_clock = "clock1";
defparam ram_block3a13.ram_block_type = "M9K";
defparam ram_block3a13.mem_init3 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a13.mem_init2 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a13.mem_init1 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a13.mem_init0 = 2048'h000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000020421000022022F5213;
// synopsys translate_on

// Location: M9K_X51_Y34_N0
cycloneive_ram_block ram_block3a46(
	.portawe(\decode4|eq_node[1]~0_combout ),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(\decode5|eq_node[1]~0_combout ),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock1),
	.ena0(!ramaddr),
	.ena1(ram_rom_addr_reg_13),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({data_a[14]}),
	.portaaddr({address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain({data_b[14]}),
	.portbaddr({address_b[12],address_b[11],address_b[10],address_b[9],address_b[8],address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.devclrn(devclrn),
	.devpor(devpor),
	.portadataout(ram_block3a46_PORTADATAOUT_bus),
	.portbdataout(ram_block3a46_PORTBDATAOUT_bus));
// synopsys translate_off
defparam ram_block3a46.clk0_core_clock_enable = "ena0";
defparam ram_block3a46.clk1_core_clock_enable = "ena1";
defparam ram_block3a46.data_interleave_offset_in_bits = 1;
defparam ram_block3a46.data_interleave_width_in_bits = 1;
defparam ram_block3a46.init_file = "meminit.hex";
defparam ram_block3a46.init_file_layout = "port_a";
defparam ram_block3a46.logical_ram_name = "ram:RAM|altsyncram:altsyncram_component|altsyncram_99f1:auto_generated|altsyncram_fta2:altsyncram1|ALTSYNCRAM";
defparam ram_block3a46.mixed_port_feed_through_mode = "dont_care";
defparam ram_block3a46.operation_mode = "bidir_dual_port";
defparam ram_block3a46.port_a_address_clear = "none";
defparam ram_block3a46.port_a_address_width = 13;
defparam ram_block3a46.port_a_byte_enable_clock = "none";
defparam ram_block3a46.port_a_data_out_clear = "none";
defparam ram_block3a46.port_a_data_out_clock = "none";
defparam ram_block3a46.port_a_data_width = 1;
defparam ram_block3a46.port_a_first_address = 0;
defparam ram_block3a46.port_a_first_bit_number = 14;
defparam ram_block3a46.port_a_last_address = 8191;
defparam ram_block3a46.port_a_logical_ram_depth = 16384;
defparam ram_block3a46.port_a_logical_ram_width = 32;
defparam ram_block3a46.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block3a46.port_b_address_clear = "none";
defparam ram_block3a46.port_b_address_clock = "clock1";
defparam ram_block3a46.port_b_address_width = 13;
defparam ram_block3a46.port_b_data_in_clock = "clock1";
defparam ram_block3a46.port_b_data_out_clear = "none";
defparam ram_block3a46.port_b_data_out_clock = "none";
defparam ram_block3a46.port_b_data_width = 1;
defparam ram_block3a46.port_b_first_address = 0;
defparam ram_block3a46.port_b_first_bit_number = 14;
defparam ram_block3a46.port_b_last_address = 8191;
defparam ram_block3a46.port_b_logical_ram_depth = 16384;
defparam ram_block3a46.port_b_logical_ram_width = 32;
defparam ram_block3a46.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block3a46.port_b_read_enable_clock = "clock1";
defparam ram_block3a46.port_b_write_enable_clock = "clock1";
defparam ram_block3a46.ram_block_type = "M9K";
defparam ram_block3a46.mem_init3 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a46.mem_init2 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a46.mem_init1 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a46.mem_init0 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
// synopsys translate_on

// Location: M9K_X51_Y38_N0
cycloneive_ram_block ram_block3a14(
	.portawe(\decode4|eq_node[0]~1_combout ),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(\decode5|eq_node[0]~1_combout ),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock1),
	.ena0(ramaddr),
	.ena1(!ram_rom_addr_reg_13),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({data_a[14]}),
	.portaaddr({address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain({data_b[14]}),
	.portbaddr({address_b[12],address_b[11],address_b[10],address_b[9],address_b[8],address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.devclrn(devclrn),
	.devpor(devpor),
	.portadataout(ram_block3a14_PORTADATAOUT_bus),
	.portbdataout(ram_block3a14_PORTBDATAOUT_bus));
// synopsys translate_off
defparam ram_block3a14.clk0_core_clock_enable = "ena0";
defparam ram_block3a14.clk1_core_clock_enable = "ena1";
defparam ram_block3a14.data_interleave_offset_in_bits = 1;
defparam ram_block3a14.data_interleave_width_in_bits = 1;
defparam ram_block3a14.init_file = "meminit.hex";
defparam ram_block3a14.init_file_layout = "port_a";
defparam ram_block3a14.logical_ram_name = "ram:RAM|altsyncram:altsyncram_component|altsyncram_99f1:auto_generated|altsyncram_fta2:altsyncram1|ALTSYNCRAM";
defparam ram_block3a14.mixed_port_feed_through_mode = "dont_care";
defparam ram_block3a14.operation_mode = "bidir_dual_port";
defparam ram_block3a14.port_a_address_clear = "none";
defparam ram_block3a14.port_a_address_width = 13;
defparam ram_block3a14.port_a_byte_enable_clock = "none";
defparam ram_block3a14.port_a_data_out_clear = "none";
defparam ram_block3a14.port_a_data_out_clock = "none";
defparam ram_block3a14.port_a_data_width = 1;
defparam ram_block3a14.port_a_first_address = 0;
defparam ram_block3a14.port_a_first_bit_number = 14;
defparam ram_block3a14.port_a_last_address = 8191;
defparam ram_block3a14.port_a_logical_ram_depth = 16384;
defparam ram_block3a14.port_a_logical_ram_width = 32;
defparam ram_block3a14.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block3a14.port_b_address_clear = "none";
defparam ram_block3a14.port_b_address_clock = "clock1";
defparam ram_block3a14.port_b_address_width = 13;
defparam ram_block3a14.port_b_data_in_clock = "clock1";
defparam ram_block3a14.port_b_data_out_clear = "none";
defparam ram_block3a14.port_b_data_out_clock = "none";
defparam ram_block3a14.port_b_data_width = 1;
defparam ram_block3a14.port_b_first_address = 0;
defparam ram_block3a14.port_b_first_bit_number = 14;
defparam ram_block3a14.port_b_last_address = 8191;
defparam ram_block3a14.port_b_logical_ram_depth = 16384;
defparam ram_block3a14.port_b_logical_ram_width = 32;
defparam ram_block3a14.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block3a14.port_b_read_enable_clock = "clock1";
defparam ram_block3a14.port_b_write_enable_clock = "clock1";
defparam ram_block3a14.ram_block_type = "M9K";
defparam ram_block3a14.mem_init3 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a14.mem_init2 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a14.mem_init1 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a14.mem_init0 = 2048'h0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000204210000224A200503;
// synopsys translate_on

// Location: M9K_X37_Y37_N0
cycloneive_ram_block ram_block3a47(
	.portawe(\decode4|eq_node[1]~0_combout ),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(\decode5|eq_node[1]~0_combout ),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock1),
	.ena0(!ramaddr),
	.ena1(ram_rom_addr_reg_13),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({data_a[15]}),
	.portaaddr({address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain({data_b[15]}),
	.portbaddr({address_b[12],address_b[11],address_b[10],address_b[9],address_b[8],address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.devclrn(devclrn),
	.devpor(devpor),
	.portadataout(ram_block3a47_PORTADATAOUT_bus),
	.portbdataout(ram_block3a47_PORTBDATAOUT_bus));
// synopsys translate_off
defparam ram_block3a47.clk0_core_clock_enable = "ena0";
defparam ram_block3a47.clk1_core_clock_enable = "ena1";
defparam ram_block3a47.data_interleave_offset_in_bits = 1;
defparam ram_block3a47.data_interleave_width_in_bits = 1;
defparam ram_block3a47.init_file = "meminit.hex";
defparam ram_block3a47.init_file_layout = "port_a";
defparam ram_block3a47.logical_ram_name = "ram:RAM|altsyncram:altsyncram_component|altsyncram_99f1:auto_generated|altsyncram_fta2:altsyncram1|ALTSYNCRAM";
defparam ram_block3a47.mixed_port_feed_through_mode = "dont_care";
defparam ram_block3a47.operation_mode = "bidir_dual_port";
defparam ram_block3a47.port_a_address_clear = "none";
defparam ram_block3a47.port_a_address_width = 13;
defparam ram_block3a47.port_a_byte_enable_clock = "none";
defparam ram_block3a47.port_a_data_out_clear = "none";
defparam ram_block3a47.port_a_data_out_clock = "none";
defparam ram_block3a47.port_a_data_width = 1;
defparam ram_block3a47.port_a_first_address = 0;
defparam ram_block3a47.port_a_first_bit_number = 15;
defparam ram_block3a47.port_a_last_address = 8191;
defparam ram_block3a47.port_a_logical_ram_depth = 16384;
defparam ram_block3a47.port_a_logical_ram_width = 32;
defparam ram_block3a47.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block3a47.port_b_address_clear = "none";
defparam ram_block3a47.port_b_address_clock = "clock1";
defparam ram_block3a47.port_b_address_width = 13;
defparam ram_block3a47.port_b_data_in_clock = "clock1";
defparam ram_block3a47.port_b_data_out_clear = "none";
defparam ram_block3a47.port_b_data_out_clock = "none";
defparam ram_block3a47.port_b_data_width = 1;
defparam ram_block3a47.port_b_first_address = 0;
defparam ram_block3a47.port_b_first_bit_number = 15;
defparam ram_block3a47.port_b_last_address = 8191;
defparam ram_block3a47.port_b_logical_ram_depth = 16384;
defparam ram_block3a47.port_b_logical_ram_width = 32;
defparam ram_block3a47.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block3a47.port_b_read_enable_clock = "clock1";
defparam ram_block3a47.port_b_write_enable_clock = "clock1";
defparam ram_block3a47.ram_block_type = "M9K";
defparam ram_block3a47.mem_init3 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a47.mem_init2 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a47.mem_init1 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a47.mem_init0 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
// synopsys translate_on

// Location: M9K_X37_Y39_N0
cycloneive_ram_block ram_block3a15(
	.portawe(\decode4|eq_node[0]~1_combout ),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(\decode5|eq_node[0]~1_combout ),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock1),
	.ena0(ramaddr),
	.ena1(!ram_rom_addr_reg_13),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({data_a[15]}),
	.portaaddr({address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain({data_b[15]}),
	.portbaddr({address_b[12],address_b[11],address_b[10],address_b[9],address_b[8],address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.devclrn(devclrn),
	.devpor(devpor),
	.portadataout(ram_block3a15_PORTADATAOUT_bus),
	.portbdataout(ram_block3a15_PORTBDATAOUT_bus));
// synopsys translate_off
defparam ram_block3a15.clk0_core_clock_enable = "ena0";
defparam ram_block3a15.clk1_core_clock_enable = "ena1";
defparam ram_block3a15.data_interleave_offset_in_bits = 1;
defparam ram_block3a15.data_interleave_width_in_bits = 1;
defparam ram_block3a15.init_file = "meminit.hex";
defparam ram_block3a15.init_file_layout = "port_a";
defparam ram_block3a15.logical_ram_name = "ram:RAM|altsyncram:altsyncram_component|altsyncram_99f1:auto_generated|altsyncram_fta2:altsyncram1|ALTSYNCRAM";
defparam ram_block3a15.mixed_port_feed_through_mode = "dont_care";
defparam ram_block3a15.operation_mode = "bidir_dual_port";
defparam ram_block3a15.port_a_address_clear = "none";
defparam ram_block3a15.port_a_address_width = 13;
defparam ram_block3a15.port_a_byte_enable_clock = "none";
defparam ram_block3a15.port_a_data_out_clear = "none";
defparam ram_block3a15.port_a_data_out_clock = "none";
defparam ram_block3a15.port_a_data_width = 1;
defparam ram_block3a15.port_a_first_address = 0;
defparam ram_block3a15.port_a_first_bit_number = 15;
defparam ram_block3a15.port_a_last_address = 8191;
defparam ram_block3a15.port_a_logical_ram_depth = 16384;
defparam ram_block3a15.port_a_logical_ram_width = 32;
defparam ram_block3a15.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block3a15.port_b_address_clear = "none";
defparam ram_block3a15.port_b_address_clock = "clock1";
defparam ram_block3a15.port_b_address_width = 13;
defparam ram_block3a15.port_b_data_in_clock = "clock1";
defparam ram_block3a15.port_b_data_out_clear = "none";
defparam ram_block3a15.port_b_data_out_clock = "none";
defparam ram_block3a15.port_b_data_width = 1;
defparam ram_block3a15.port_b_first_address = 0;
defparam ram_block3a15.port_b_first_bit_number = 15;
defparam ram_block3a15.port_b_last_address = 8191;
defparam ram_block3a15.port_b_logical_ram_depth = 16384;
defparam ram_block3a15.port_b_logical_ram_width = 32;
defparam ram_block3a15.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block3a15.port_b_read_enable_clock = "clock1";
defparam ram_block3a15.port_b_write_enable_clock = "clock1";
defparam ram_block3a15.ram_block_type = "M9K";
defparam ram_block3a15.mem_init3 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a15.mem_init2 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a15.mem_init1 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a15.mem_init0 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000002042100002242206063;
// synopsys translate_on

// Location: M9K_X37_Y27_N0
cycloneive_ram_block ram_block3a48(
	.portawe(\decode4|eq_node[1]~0_combout ),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(\decode5|eq_node[1]~0_combout ),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock1),
	.ena0(!ramaddr),
	.ena1(ram_rom_addr_reg_13),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({data_a[16]}),
	.portaaddr({address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain({data_b[16]}),
	.portbaddr({address_b[12],address_b[11],address_b[10],address_b[9],address_b[8],address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.devclrn(devclrn),
	.devpor(devpor),
	.portadataout(ram_block3a48_PORTADATAOUT_bus),
	.portbdataout(ram_block3a48_PORTBDATAOUT_bus));
// synopsys translate_off
defparam ram_block3a48.clk0_core_clock_enable = "ena0";
defparam ram_block3a48.clk1_core_clock_enable = "ena1";
defparam ram_block3a48.data_interleave_offset_in_bits = 1;
defparam ram_block3a48.data_interleave_width_in_bits = 1;
defparam ram_block3a48.init_file = "meminit.hex";
defparam ram_block3a48.init_file_layout = "port_a";
defparam ram_block3a48.logical_ram_name = "ram:RAM|altsyncram:altsyncram_component|altsyncram_99f1:auto_generated|altsyncram_fta2:altsyncram1|ALTSYNCRAM";
defparam ram_block3a48.mixed_port_feed_through_mode = "dont_care";
defparam ram_block3a48.operation_mode = "bidir_dual_port";
defparam ram_block3a48.port_a_address_clear = "none";
defparam ram_block3a48.port_a_address_width = 13;
defparam ram_block3a48.port_a_byte_enable_clock = "none";
defparam ram_block3a48.port_a_data_out_clear = "none";
defparam ram_block3a48.port_a_data_out_clock = "none";
defparam ram_block3a48.port_a_data_width = 1;
defparam ram_block3a48.port_a_first_address = 0;
defparam ram_block3a48.port_a_first_bit_number = 16;
defparam ram_block3a48.port_a_last_address = 8191;
defparam ram_block3a48.port_a_logical_ram_depth = 16384;
defparam ram_block3a48.port_a_logical_ram_width = 32;
defparam ram_block3a48.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block3a48.port_b_address_clear = "none";
defparam ram_block3a48.port_b_address_clock = "clock1";
defparam ram_block3a48.port_b_address_width = 13;
defparam ram_block3a48.port_b_data_in_clock = "clock1";
defparam ram_block3a48.port_b_data_out_clear = "none";
defparam ram_block3a48.port_b_data_out_clock = "none";
defparam ram_block3a48.port_b_data_width = 1;
defparam ram_block3a48.port_b_first_address = 0;
defparam ram_block3a48.port_b_first_bit_number = 16;
defparam ram_block3a48.port_b_last_address = 8191;
defparam ram_block3a48.port_b_logical_ram_depth = 16384;
defparam ram_block3a48.port_b_logical_ram_width = 32;
defparam ram_block3a48.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block3a48.port_b_read_enable_clock = "clock1";
defparam ram_block3a48.port_b_write_enable_clock = "clock1";
defparam ram_block3a48.ram_block_type = "M9K";
defparam ram_block3a48.mem_init3 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a48.mem_init2 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a48.mem_init1 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a48.mem_init0 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
// synopsys translate_on

// Location: M9K_X37_Y31_N0
cycloneive_ram_block ram_block3a16(
	.portawe(\decode4|eq_node[0]~1_combout ),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(\decode5|eq_node[0]~1_combout ),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock1),
	.ena0(ramaddr),
	.ena1(!ram_rom_addr_reg_13),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({data_a[16]}),
	.portaaddr({address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain({data_b[16]}),
	.portbaddr({address_b[12],address_b[11],address_b[10],address_b[9],address_b[8],address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.devclrn(devclrn),
	.devpor(devpor),
	.portadataout(ram_block3a16_PORTADATAOUT_bus),
	.portbdataout(ram_block3a16_PORTBDATAOUT_bus));
// synopsys translate_off
defparam ram_block3a16.clk0_core_clock_enable = "ena0";
defparam ram_block3a16.clk1_core_clock_enable = "ena1";
defparam ram_block3a16.data_interleave_offset_in_bits = 1;
defparam ram_block3a16.data_interleave_width_in_bits = 1;
defparam ram_block3a16.init_file = "meminit.hex";
defparam ram_block3a16.init_file_layout = "port_a";
defparam ram_block3a16.logical_ram_name = "ram:RAM|altsyncram:altsyncram_component|altsyncram_99f1:auto_generated|altsyncram_fta2:altsyncram1|ALTSYNCRAM";
defparam ram_block3a16.mixed_port_feed_through_mode = "dont_care";
defparam ram_block3a16.operation_mode = "bidir_dual_port";
defparam ram_block3a16.port_a_address_clear = "none";
defparam ram_block3a16.port_a_address_width = 13;
defparam ram_block3a16.port_a_byte_enable_clock = "none";
defparam ram_block3a16.port_a_data_out_clear = "none";
defparam ram_block3a16.port_a_data_out_clock = "none";
defparam ram_block3a16.port_a_data_width = 1;
defparam ram_block3a16.port_a_first_address = 0;
defparam ram_block3a16.port_a_first_bit_number = 16;
defparam ram_block3a16.port_a_last_address = 8191;
defparam ram_block3a16.port_a_logical_ram_depth = 16384;
defparam ram_block3a16.port_a_logical_ram_width = 32;
defparam ram_block3a16.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block3a16.port_b_address_clear = "none";
defparam ram_block3a16.port_b_address_clock = "clock1";
defparam ram_block3a16.port_b_address_width = 13;
defparam ram_block3a16.port_b_data_in_clock = "clock1";
defparam ram_block3a16.port_b_data_out_clear = "none";
defparam ram_block3a16.port_b_data_out_clock = "none";
defparam ram_block3a16.port_b_data_width = 1;
defparam ram_block3a16.port_b_first_address = 0;
defparam ram_block3a16.port_b_first_bit_number = 16;
defparam ram_block3a16.port_b_last_address = 8191;
defparam ram_block3a16.port_b_logical_ram_depth = 16384;
defparam ram_block3a16.port_b_logical_ram_width = 32;
defparam ram_block3a16.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block3a16.port_b_read_enable_clock = "clock1";
defparam ram_block3a16.port_b_write_enable_clock = "clock1";
defparam ram_block3a16.ram_block_type = "M9K";
defparam ram_block3a16.mem_init3 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a16.mem_init2 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a16.mem_init1 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a16.mem_init0 = 2048'h0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000205A122003613254042;
// synopsys translate_on

// Location: M9K_X64_Y35_N0
cycloneive_ram_block ram_block3a49(
	.portawe(\decode4|eq_node[1]~0_combout ),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(\decode5|eq_node[1]~0_combout ),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock1),
	.ena0(!ramaddr),
	.ena1(ram_rom_addr_reg_13),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({data_a[17]}),
	.portaaddr({address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain({data_b[17]}),
	.portbaddr({address_b[12],address_b[11],address_b[10],address_b[9],address_b[8],address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.devclrn(devclrn),
	.devpor(devpor),
	.portadataout(ram_block3a49_PORTADATAOUT_bus),
	.portbdataout(ram_block3a49_PORTBDATAOUT_bus));
// synopsys translate_off
defparam ram_block3a49.clk0_core_clock_enable = "ena0";
defparam ram_block3a49.clk1_core_clock_enable = "ena1";
defparam ram_block3a49.data_interleave_offset_in_bits = 1;
defparam ram_block3a49.data_interleave_width_in_bits = 1;
defparam ram_block3a49.init_file = "meminit.hex";
defparam ram_block3a49.init_file_layout = "port_a";
defparam ram_block3a49.logical_ram_name = "ram:RAM|altsyncram:altsyncram_component|altsyncram_99f1:auto_generated|altsyncram_fta2:altsyncram1|ALTSYNCRAM";
defparam ram_block3a49.mixed_port_feed_through_mode = "dont_care";
defparam ram_block3a49.operation_mode = "bidir_dual_port";
defparam ram_block3a49.port_a_address_clear = "none";
defparam ram_block3a49.port_a_address_width = 13;
defparam ram_block3a49.port_a_byte_enable_clock = "none";
defparam ram_block3a49.port_a_data_out_clear = "none";
defparam ram_block3a49.port_a_data_out_clock = "none";
defparam ram_block3a49.port_a_data_width = 1;
defparam ram_block3a49.port_a_first_address = 0;
defparam ram_block3a49.port_a_first_bit_number = 17;
defparam ram_block3a49.port_a_last_address = 8191;
defparam ram_block3a49.port_a_logical_ram_depth = 16384;
defparam ram_block3a49.port_a_logical_ram_width = 32;
defparam ram_block3a49.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block3a49.port_b_address_clear = "none";
defparam ram_block3a49.port_b_address_clock = "clock1";
defparam ram_block3a49.port_b_address_width = 13;
defparam ram_block3a49.port_b_data_in_clock = "clock1";
defparam ram_block3a49.port_b_data_out_clear = "none";
defparam ram_block3a49.port_b_data_out_clock = "none";
defparam ram_block3a49.port_b_data_width = 1;
defparam ram_block3a49.port_b_first_address = 0;
defparam ram_block3a49.port_b_first_bit_number = 17;
defparam ram_block3a49.port_b_last_address = 8191;
defparam ram_block3a49.port_b_logical_ram_depth = 16384;
defparam ram_block3a49.port_b_logical_ram_width = 32;
defparam ram_block3a49.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block3a49.port_b_read_enable_clock = "clock1";
defparam ram_block3a49.port_b_write_enable_clock = "clock1";
defparam ram_block3a49.ram_block_type = "M9K";
defparam ram_block3a49.mem_init3 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a49.mem_init2 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a49.mem_init1 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a49.mem_init0 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
// synopsys translate_on

// Location: M9K_X64_Y39_N0
cycloneive_ram_block ram_block3a17(
	.portawe(\decode4|eq_node[0]~1_combout ),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(\decode5|eq_node[0]~1_combout ),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock1),
	.ena0(ramaddr),
	.ena1(!ram_rom_addr_reg_13),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({data_a[17]}),
	.portaaddr({address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain({data_b[17]}),
	.portbaddr({address_b[12],address_b[11],address_b[10],address_b[9],address_b[8],address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.devclrn(devclrn),
	.devpor(devpor),
	.portadataout(ram_block3a17_PORTADATAOUT_bus),
	.portbdataout(ram_block3a17_PORTBDATAOUT_bus));
// synopsys translate_off
defparam ram_block3a17.clk0_core_clock_enable = "ena0";
defparam ram_block3a17.clk1_core_clock_enable = "ena1";
defparam ram_block3a17.data_interleave_offset_in_bits = 1;
defparam ram_block3a17.data_interleave_width_in_bits = 1;
defparam ram_block3a17.init_file = "meminit.hex";
defparam ram_block3a17.init_file_layout = "port_a";
defparam ram_block3a17.logical_ram_name = "ram:RAM|altsyncram:altsyncram_component|altsyncram_99f1:auto_generated|altsyncram_fta2:altsyncram1|ALTSYNCRAM";
defparam ram_block3a17.mixed_port_feed_through_mode = "dont_care";
defparam ram_block3a17.operation_mode = "bidir_dual_port";
defparam ram_block3a17.port_a_address_clear = "none";
defparam ram_block3a17.port_a_address_width = 13;
defparam ram_block3a17.port_a_byte_enable_clock = "none";
defparam ram_block3a17.port_a_data_out_clear = "none";
defparam ram_block3a17.port_a_data_out_clock = "none";
defparam ram_block3a17.port_a_data_width = 1;
defparam ram_block3a17.port_a_first_address = 0;
defparam ram_block3a17.port_a_first_bit_number = 17;
defparam ram_block3a17.port_a_last_address = 8191;
defparam ram_block3a17.port_a_logical_ram_depth = 16384;
defparam ram_block3a17.port_a_logical_ram_width = 32;
defparam ram_block3a17.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block3a17.port_b_address_clear = "none";
defparam ram_block3a17.port_b_address_clock = "clock1";
defparam ram_block3a17.port_b_address_width = 13;
defparam ram_block3a17.port_b_data_in_clock = "clock1";
defparam ram_block3a17.port_b_data_out_clear = "none";
defparam ram_block3a17.port_b_data_out_clock = "none";
defparam ram_block3a17.port_b_data_width = 1;
defparam ram_block3a17.port_b_first_address = 0;
defparam ram_block3a17.port_b_first_bit_number = 17;
defparam ram_block3a17.port_b_last_address = 8191;
defparam ram_block3a17.port_b_logical_ram_depth = 16384;
defparam ram_block3a17.port_b_logical_ram_width = 32;
defparam ram_block3a17.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block3a17.port_b_read_enable_clock = "clock1";
defparam ram_block3a17.port_b_write_enable_clock = "clock1";
defparam ram_block3a17.ram_block_type = "M9K";
defparam ram_block3a17.mem_init3 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a17.mem_init2 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a17.mem_init1 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a17.mem_init0 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000006C0340C001602060001;
// synopsys translate_on

// Location: M9K_X51_Y24_N0
cycloneive_ram_block ram_block3a50(
	.portawe(\decode4|eq_node[1]~0_combout ),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(\decode5|eq_node[1]~0_combout ),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock1),
	.ena0(!ramaddr),
	.ena1(ram_rom_addr_reg_13),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({data_a[18]}),
	.portaaddr({address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain({data_b[18]}),
	.portbaddr({address_b[12],address_b[11],address_b[10],address_b[9],address_b[8],address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.devclrn(devclrn),
	.devpor(devpor),
	.portadataout(ram_block3a50_PORTADATAOUT_bus),
	.portbdataout(ram_block3a50_PORTBDATAOUT_bus));
// synopsys translate_off
defparam ram_block3a50.clk0_core_clock_enable = "ena0";
defparam ram_block3a50.clk1_core_clock_enable = "ena1";
defparam ram_block3a50.data_interleave_offset_in_bits = 1;
defparam ram_block3a50.data_interleave_width_in_bits = 1;
defparam ram_block3a50.init_file = "meminit.hex";
defparam ram_block3a50.init_file_layout = "port_a";
defparam ram_block3a50.logical_ram_name = "ram:RAM|altsyncram:altsyncram_component|altsyncram_99f1:auto_generated|altsyncram_fta2:altsyncram1|ALTSYNCRAM";
defparam ram_block3a50.mixed_port_feed_through_mode = "dont_care";
defparam ram_block3a50.operation_mode = "bidir_dual_port";
defparam ram_block3a50.port_a_address_clear = "none";
defparam ram_block3a50.port_a_address_width = 13;
defparam ram_block3a50.port_a_byte_enable_clock = "none";
defparam ram_block3a50.port_a_data_out_clear = "none";
defparam ram_block3a50.port_a_data_out_clock = "none";
defparam ram_block3a50.port_a_data_width = 1;
defparam ram_block3a50.port_a_first_address = 0;
defparam ram_block3a50.port_a_first_bit_number = 18;
defparam ram_block3a50.port_a_last_address = 8191;
defparam ram_block3a50.port_a_logical_ram_depth = 16384;
defparam ram_block3a50.port_a_logical_ram_width = 32;
defparam ram_block3a50.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block3a50.port_b_address_clear = "none";
defparam ram_block3a50.port_b_address_clock = "clock1";
defparam ram_block3a50.port_b_address_width = 13;
defparam ram_block3a50.port_b_data_in_clock = "clock1";
defparam ram_block3a50.port_b_data_out_clear = "none";
defparam ram_block3a50.port_b_data_out_clock = "none";
defparam ram_block3a50.port_b_data_width = 1;
defparam ram_block3a50.port_b_first_address = 0;
defparam ram_block3a50.port_b_first_bit_number = 18;
defparam ram_block3a50.port_b_last_address = 8191;
defparam ram_block3a50.port_b_logical_ram_depth = 16384;
defparam ram_block3a50.port_b_logical_ram_width = 32;
defparam ram_block3a50.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block3a50.port_b_read_enable_clock = "clock1";
defparam ram_block3a50.port_b_write_enable_clock = "clock1";
defparam ram_block3a50.ram_block_type = "M9K";
defparam ram_block3a50.mem_init3 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a50.mem_init2 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a50.mem_init1 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a50.mem_init0 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
// synopsys translate_on

// Location: M9K_X64_Y24_N0
cycloneive_ram_block ram_block3a18(
	.portawe(\decode4|eq_node[0]~1_combout ),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(\decode5|eq_node[0]~1_combout ),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock1),
	.ena0(ramaddr),
	.ena1(!ram_rom_addr_reg_13),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({data_a[18]}),
	.portaaddr({address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain({data_b[18]}),
	.portbaddr({address_b[12],address_b[11],address_b[10],address_b[9],address_b[8],address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.devclrn(devclrn),
	.devpor(devpor),
	.portadataout(ram_block3a18_PORTADATAOUT_bus),
	.portbdataout(ram_block3a18_PORTBDATAOUT_bus));
// synopsys translate_off
defparam ram_block3a18.clk0_core_clock_enable = "ena0";
defparam ram_block3a18.clk1_core_clock_enable = "ena1";
defparam ram_block3a18.data_interleave_offset_in_bits = 1;
defparam ram_block3a18.data_interleave_width_in_bits = 1;
defparam ram_block3a18.init_file = "meminit.hex";
defparam ram_block3a18.init_file_layout = "port_a";
defparam ram_block3a18.logical_ram_name = "ram:RAM|altsyncram:altsyncram_component|altsyncram_99f1:auto_generated|altsyncram_fta2:altsyncram1|ALTSYNCRAM";
defparam ram_block3a18.mixed_port_feed_through_mode = "dont_care";
defparam ram_block3a18.operation_mode = "bidir_dual_port";
defparam ram_block3a18.port_a_address_clear = "none";
defparam ram_block3a18.port_a_address_width = 13;
defparam ram_block3a18.port_a_byte_enable_clock = "none";
defparam ram_block3a18.port_a_data_out_clear = "none";
defparam ram_block3a18.port_a_data_out_clock = "none";
defparam ram_block3a18.port_a_data_width = 1;
defparam ram_block3a18.port_a_first_address = 0;
defparam ram_block3a18.port_a_first_bit_number = 18;
defparam ram_block3a18.port_a_last_address = 8191;
defparam ram_block3a18.port_a_logical_ram_depth = 16384;
defparam ram_block3a18.port_a_logical_ram_width = 32;
defparam ram_block3a18.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block3a18.port_b_address_clear = "none";
defparam ram_block3a18.port_b_address_clock = "clock1";
defparam ram_block3a18.port_b_address_width = 13;
defparam ram_block3a18.port_b_data_in_clock = "clock1";
defparam ram_block3a18.port_b_data_out_clear = "none";
defparam ram_block3a18.port_b_data_out_clock = "none";
defparam ram_block3a18.port_b_data_width = 1;
defparam ram_block3a18.port_b_first_address = 0;
defparam ram_block3a18.port_b_first_bit_number = 18;
defparam ram_block3a18.port_b_last_address = 8191;
defparam ram_block3a18.port_b_logical_ram_depth = 16384;
defparam ram_block3a18.port_b_logical_ram_width = 32;
defparam ram_block3a18.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block3a18.port_b_read_enable_clock = "clock1";
defparam ram_block3a18.port_b_write_enable_clock = "clock1";
defparam ram_block3a18.ram_block_type = "M9K";
defparam ram_block3a18.mem_init3 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a18.mem_init2 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a18.mem_init1 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a18.mem_init0 = 2048'h000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000060C3180001703286867;
// synopsys translate_on

// Location: M9K_X64_Y36_N0
cycloneive_ram_block ram_block3a51(
	.portawe(\decode4|eq_node[1]~0_combout ),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(\decode5|eq_node[1]~0_combout ),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock1),
	.ena0(!ramaddr),
	.ena1(ram_rom_addr_reg_13),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({data_a[19]}),
	.portaaddr({address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain({data_b[19]}),
	.portbaddr({address_b[12],address_b[11],address_b[10],address_b[9],address_b[8],address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.devclrn(devclrn),
	.devpor(devpor),
	.portadataout(ram_block3a51_PORTADATAOUT_bus),
	.portbdataout(ram_block3a51_PORTBDATAOUT_bus));
// synopsys translate_off
defparam ram_block3a51.clk0_core_clock_enable = "ena0";
defparam ram_block3a51.clk1_core_clock_enable = "ena1";
defparam ram_block3a51.data_interleave_offset_in_bits = 1;
defparam ram_block3a51.data_interleave_width_in_bits = 1;
defparam ram_block3a51.init_file = "meminit.hex";
defparam ram_block3a51.init_file_layout = "port_a";
defparam ram_block3a51.logical_ram_name = "ram:RAM|altsyncram:altsyncram_component|altsyncram_99f1:auto_generated|altsyncram_fta2:altsyncram1|ALTSYNCRAM";
defparam ram_block3a51.mixed_port_feed_through_mode = "dont_care";
defparam ram_block3a51.operation_mode = "bidir_dual_port";
defparam ram_block3a51.port_a_address_clear = "none";
defparam ram_block3a51.port_a_address_width = 13;
defparam ram_block3a51.port_a_byte_enable_clock = "none";
defparam ram_block3a51.port_a_data_out_clear = "none";
defparam ram_block3a51.port_a_data_out_clock = "none";
defparam ram_block3a51.port_a_data_width = 1;
defparam ram_block3a51.port_a_first_address = 0;
defparam ram_block3a51.port_a_first_bit_number = 19;
defparam ram_block3a51.port_a_last_address = 8191;
defparam ram_block3a51.port_a_logical_ram_depth = 16384;
defparam ram_block3a51.port_a_logical_ram_width = 32;
defparam ram_block3a51.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block3a51.port_b_address_clear = "none";
defparam ram_block3a51.port_b_address_clock = "clock1";
defparam ram_block3a51.port_b_address_width = 13;
defparam ram_block3a51.port_b_data_in_clock = "clock1";
defparam ram_block3a51.port_b_data_out_clear = "none";
defparam ram_block3a51.port_b_data_out_clock = "none";
defparam ram_block3a51.port_b_data_width = 1;
defparam ram_block3a51.port_b_first_address = 0;
defparam ram_block3a51.port_b_first_bit_number = 19;
defparam ram_block3a51.port_b_last_address = 8191;
defparam ram_block3a51.port_b_logical_ram_depth = 16384;
defparam ram_block3a51.port_b_logical_ram_width = 32;
defparam ram_block3a51.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block3a51.port_b_read_enable_clock = "clock1";
defparam ram_block3a51.port_b_write_enable_clock = "clock1";
defparam ram_block3a51.ram_block_type = "M9K";
defparam ram_block3a51.mem_init3 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a51.mem_init2 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a51.mem_init1 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a51.mem_init0 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
// synopsys translate_on

// Location: M9K_X64_Y37_N0
cycloneive_ram_block ram_block3a19(
	.portawe(\decode4|eq_node[0]~1_combout ),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(\decode5|eq_node[0]~1_combout ),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock1),
	.ena0(ramaddr),
	.ena1(!ram_rom_addr_reg_13),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({data_a[19]}),
	.portaaddr({address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain({data_b[19]}),
	.portbaddr({address_b[12],address_b[11],address_b[10],address_b[9],address_b[8],address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.devclrn(devclrn),
	.devpor(devpor),
	.portadataout(ram_block3a19_PORTADATAOUT_bus),
	.portbdataout(ram_block3a19_PORTBDATAOUT_bus));
// synopsys translate_off
defparam ram_block3a19.clk0_core_clock_enable = "ena0";
defparam ram_block3a19.clk1_core_clock_enable = "ena1";
defparam ram_block3a19.data_interleave_offset_in_bits = 1;
defparam ram_block3a19.data_interleave_width_in_bits = 1;
defparam ram_block3a19.init_file = "meminit.hex";
defparam ram_block3a19.init_file_layout = "port_a";
defparam ram_block3a19.logical_ram_name = "ram:RAM|altsyncram:altsyncram_component|altsyncram_99f1:auto_generated|altsyncram_fta2:altsyncram1|ALTSYNCRAM";
defparam ram_block3a19.mixed_port_feed_through_mode = "dont_care";
defparam ram_block3a19.operation_mode = "bidir_dual_port";
defparam ram_block3a19.port_a_address_clear = "none";
defparam ram_block3a19.port_a_address_width = 13;
defparam ram_block3a19.port_a_byte_enable_clock = "none";
defparam ram_block3a19.port_a_data_out_clear = "none";
defparam ram_block3a19.port_a_data_out_clock = "none";
defparam ram_block3a19.port_a_data_width = 1;
defparam ram_block3a19.port_a_first_address = 0;
defparam ram_block3a19.port_a_first_bit_number = 19;
defparam ram_block3a19.port_a_last_address = 8191;
defparam ram_block3a19.port_a_logical_ram_depth = 16384;
defparam ram_block3a19.port_a_logical_ram_width = 32;
defparam ram_block3a19.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block3a19.port_b_address_clear = "none";
defparam ram_block3a19.port_b_address_clock = "clock1";
defparam ram_block3a19.port_b_address_width = 13;
defparam ram_block3a19.port_b_data_in_clock = "clock1";
defparam ram_block3a19.port_b_data_out_clear = "none";
defparam ram_block3a19.port_b_data_out_clock = "none";
defparam ram_block3a19.port_b_data_width = 1;
defparam ram_block3a19.port_b_first_address = 0;
defparam ram_block3a19.port_b_first_bit_number = 19;
defparam ram_block3a19.port_b_last_address = 8191;
defparam ram_block3a19.port_b_logical_ram_depth = 16384;
defparam ram_block3a19.port_b_logical_ram_width = 32;
defparam ram_block3a19.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block3a19.port_b_read_enable_clock = "clock1";
defparam ram_block3a19.port_b_write_enable_clock = "clock1";
defparam ram_block3a19.ram_block_type = "M9K";
defparam ram_block3a19.mem_init3 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a19.mem_init2 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a19.mem_init1 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a19.mem_init0 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001C38C6E09B6D7701203;
// synopsys translate_on

// Location: M9K_X64_Y34_N0
cycloneive_ram_block ram_block3a52(
	.portawe(\decode4|eq_node[1]~0_combout ),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(\decode5|eq_node[1]~0_combout ),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock1),
	.ena0(!ramaddr),
	.ena1(ram_rom_addr_reg_13),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({data_a[20]}),
	.portaaddr({address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain({data_b[20]}),
	.portbaddr({address_b[12],address_b[11],address_b[10],address_b[9],address_b[8],address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.devclrn(devclrn),
	.devpor(devpor),
	.portadataout(ram_block3a52_PORTADATAOUT_bus),
	.portbdataout(ram_block3a52_PORTBDATAOUT_bus));
// synopsys translate_off
defparam ram_block3a52.clk0_core_clock_enable = "ena0";
defparam ram_block3a52.clk1_core_clock_enable = "ena1";
defparam ram_block3a52.data_interleave_offset_in_bits = 1;
defparam ram_block3a52.data_interleave_width_in_bits = 1;
defparam ram_block3a52.init_file = "meminit.hex";
defparam ram_block3a52.init_file_layout = "port_a";
defparam ram_block3a52.logical_ram_name = "ram:RAM|altsyncram:altsyncram_component|altsyncram_99f1:auto_generated|altsyncram_fta2:altsyncram1|ALTSYNCRAM";
defparam ram_block3a52.mixed_port_feed_through_mode = "dont_care";
defparam ram_block3a52.operation_mode = "bidir_dual_port";
defparam ram_block3a52.port_a_address_clear = "none";
defparam ram_block3a52.port_a_address_width = 13;
defparam ram_block3a52.port_a_byte_enable_clock = "none";
defparam ram_block3a52.port_a_data_out_clear = "none";
defparam ram_block3a52.port_a_data_out_clock = "none";
defparam ram_block3a52.port_a_data_width = 1;
defparam ram_block3a52.port_a_first_address = 0;
defparam ram_block3a52.port_a_first_bit_number = 20;
defparam ram_block3a52.port_a_last_address = 8191;
defparam ram_block3a52.port_a_logical_ram_depth = 16384;
defparam ram_block3a52.port_a_logical_ram_width = 32;
defparam ram_block3a52.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block3a52.port_b_address_clear = "none";
defparam ram_block3a52.port_b_address_clock = "clock1";
defparam ram_block3a52.port_b_address_width = 13;
defparam ram_block3a52.port_b_data_in_clock = "clock1";
defparam ram_block3a52.port_b_data_out_clear = "none";
defparam ram_block3a52.port_b_data_out_clock = "none";
defparam ram_block3a52.port_b_data_width = 1;
defparam ram_block3a52.port_b_first_address = 0;
defparam ram_block3a52.port_b_first_bit_number = 20;
defparam ram_block3a52.port_b_last_address = 8191;
defparam ram_block3a52.port_b_logical_ram_depth = 16384;
defparam ram_block3a52.port_b_logical_ram_width = 32;
defparam ram_block3a52.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block3a52.port_b_read_enable_clock = "clock1";
defparam ram_block3a52.port_b_write_enable_clock = "clock1";
defparam ram_block3a52.ram_block_type = "M9K";
defparam ram_block3a52.mem_init3 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a52.mem_init2 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a52.mem_init1 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a52.mem_init0 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
// synopsys translate_on

// Location: M9K_X64_Y33_N0
cycloneive_ram_block ram_block3a20(
	.portawe(\decode4|eq_node[0]~1_combout ),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(\decode5|eq_node[0]~1_combout ),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock1),
	.ena0(ramaddr),
	.ena1(!ram_rom_addr_reg_13),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({data_a[20]}),
	.portaaddr({address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain({data_b[20]}),
	.portbaddr({address_b[12],address_b[11],address_b[10],address_b[9],address_b[8],address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.devclrn(devclrn),
	.devpor(devpor),
	.portadataout(ram_block3a20_PORTADATAOUT_bus),
	.portbdataout(ram_block3a20_PORTBDATAOUT_bus));
// synopsys translate_off
defparam ram_block3a20.clk0_core_clock_enable = "ena0";
defparam ram_block3a20.clk1_core_clock_enable = "ena1";
defparam ram_block3a20.data_interleave_offset_in_bits = 1;
defparam ram_block3a20.data_interleave_width_in_bits = 1;
defparam ram_block3a20.init_file = "meminit.hex";
defparam ram_block3a20.init_file_layout = "port_a";
defparam ram_block3a20.logical_ram_name = "ram:RAM|altsyncram:altsyncram_component|altsyncram_99f1:auto_generated|altsyncram_fta2:altsyncram1|ALTSYNCRAM";
defparam ram_block3a20.mixed_port_feed_through_mode = "dont_care";
defparam ram_block3a20.operation_mode = "bidir_dual_port";
defparam ram_block3a20.port_a_address_clear = "none";
defparam ram_block3a20.port_a_address_width = 13;
defparam ram_block3a20.port_a_byte_enable_clock = "none";
defparam ram_block3a20.port_a_data_out_clear = "none";
defparam ram_block3a20.port_a_data_out_clock = "none";
defparam ram_block3a20.port_a_data_width = 1;
defparam ram_block3a20.port_a_first_address = 0;
defparam ram_block3a20.port_a_first_bit_number = 20;
defparam ram_block3a20.port_a_last_address = 8191;
defparam ram_block3a20.port_a_logical_ram_depth = 16384;
defparam ram_block3a20.port_a_logical_ram_width = 32;
defparam ram_block3a20.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block3a20.port_b_address_clear = "none";
defparam ram_block3a20.port_b_address_clock = "clock1";
defparam ram_block3a20.port_b_address_width = 13;
defparam ram_block3a20.port_b_data_in_clock = "clock1";
defparam ram_block3a20.port_b_data_out_clear = "none";
defparam ram_block3a20.port_b_data_out_clock = "none";
defparam ram_block3a20.port_b_data_width = 1;
defparam ram_block3a20.port_b_first_address = 0;
defparam ram_block3a20.port_b_first_bit_number = 20;
defparam ram_block3a20.port_b_last_address = 8191;
defparam ram_block3a20.port_b_logical_ram_depth = 16384;
defparam ram_block3a20.port_b_logical_ram_width = 32;
defparam ram_block3a20.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block3a20.port_b_read_enable_clock = "clock1";
defparam ram_block3a20.port_b_write_enable_clock = "clock1";
defparam ram_block3a20.ram_block_type = "M9K";
defparam ram_block3a20.mem_init3 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a20.mem_init2 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a20.mem_init1 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a20.mem_init0 = 2048'h0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000A0832F000B;
// synopsys translate_on

// Location: M9K_X78_Y32_N0
cycloneive_ram_block ram_block3a53(
	.portawe(\decode4|eq_node[1]~0_combout ),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(\decode5|eq_node[1]~0_combout ),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock1),
	.ena0(!ramaddr),
	.ena1(ram_rom_addr_reg_13),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({data_a[21]}),
	.portaaddr({address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain({data_b[21]}),
	.portbaddr({address_b[12],address_b[11],address_b[10],address_b[9],address_b[8],address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.devclrn(devclrn),
	.devpor(devpor),
	.portadataout(ram_block3a53_PORTADATAOUT_bus),
	.portbdataout(ram_block3a53_PORTBDATAOUT_bus));
// synopsys translate_off
defparam ram_block3a53.clk0_core_clock_enable = "ena0";
defparam ram_block3a53.clk1_core_clock_enable = "ena1";
defparam ram_block3a53.data_interleave_offset_in_bits = 1;
defparam ram_block3a53.data_interleave_width_in_bits = 1;
defparam ram_block3a53.init_file = "meminit.hex";
defparam ram_block3a53.init_file_layout = "port_a";
defparam ram_block3a53.logical_ram_name = "ram:RAM|altsyncram:altsyncram_component|altsyncram_99f1:auto_generated|altsyncram_fta2:altsyncram1|ALTSYNCRAM";
defparam ram_block3a53.mixed_port_feed_through_mode = "dont_care";
defparam ram_block3a53.operation_mode = "bidir_dual_port";
defparam ram_block3a53.port_a_address_clear = "none";
defparam ram_block3a53.port_a_address_width = 13;
defparam ram_block3a53.port_a_byte_enable_clock = "none";
defparam ram_block3a53.port_a_data_out_clear = "none";
defparam ram_block3a53.port_a_data_out_clock = "none";
defparam ram_block3a53.port_a_data_width = 1;
defparam ram_block3a53.port_a_first_address = 0;
defparam ram_block3a53.port_a_first_bit_number = 21;
defparam ram_block3a53.port_a_last_address = 8191;
defparam ram_block3a53.port_a_logical_ram_depth = 16384;
defparam ram_block3a53.port_a_logical_ram_width = 32;
defparam ram_block3a53.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block3a53.port_b_address_clear = "none";
defparam ram_block3a53.port_b_address_clock = "clock1";
defparam ram_block3a53.port_b_address_width = 13;
defparam ram_block3a53.port_b_data_in_clock = "clock1";
defparam ram_block3a53.port_b_data_out_clear = "none";
defparam ram_block3a53.port_b_data_out_clock = "none";
defparam ram_block3a53.port_b_data_width = 1;
defparam ram_block3a53.port_b_first_address = 0;
defparam ram_block3a53.port_b_first_bit_number = 21;
defparam ram_block3a53.port_b_last_address = 8191;
defparam ram_block3a53.port_b_logical_ram_depth = 16384;
defparam ram_block3a53.port_b_logical_ram_width = 32;
defparam ram_block3a53.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block3a53.port_b_read_enable_clock = "clock1";
defparam ram_block3a53.port_b_write_enable_clock = "clock1";
defparam ram_block3a53.ram_block_type = "M9K";
defparam ram_block3a53.mem_init3 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a53.mem_init2 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a53.mem_init1 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a53.mem_init0 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
// synopsys translate_on

// Location: M9K_X78_Y28_N0
cycloneive_ram_block ram_block3a21(
	.portawe(\decode4|eq_node[0]~1_combout ),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(\decode5|eq_node[0]~1_combout ),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock1),
	.ena0(ramaddr),
	.ena1(!ram_rom_addr_reg_13),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({data_a[21]}),
	.portaaddr({address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain({data_b[21]}),
	.portbaddr({address_b[12],address_b[11],address_b[10],address_b[9],address_b[8],address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.devclrn(devclrn),
	.devpor(devpor),
	.portadataout(ram_block3a21_PORTADATAOUT_bus),
	.portbdataout(ram_block3a21_PORTBDATAOUT_bus));
// synopsys translate_off
defparam ram_block3a21.clk0_core_clock_enable = "ena0";
defparam ram_block3a21.clk1_core_clock_enable = "ena1";
defparam ram_block3a21.data_interleave_offset_in_bits = 1;
defparam ram_block3a21.data_interleave_width_in_bits = 1;
defparam ram_block3a21.init_file = "meminit.hex";
defparam ram_block3a21.init_file_layout = "port_a";
defparam ram_block3a21.logical_ram_name = "ram:RAM|altsyncram:altsyncram_component|altsyncram_99f1:auto_generated|altsyncram_fta2:altsyncram1|ALTSYNCRAM";
defparam ram_block3a21.mixed_port_feed_through_mode = "dont_care";
defparam ram_block3a21.operation_mode = "bidir_dual_port";
defparam ram_block3a21.port_a_address_clear = "none";
defparam ram_block3a21.port_a_address_width = 13;
defparam ram_block3a21.port_a_byte_enable_clock = "none";
defparam ram_block3a21.port_a_data_out_clear = "none";
defparam ram_block3a21.port_a_data_out_clock = "none";
defparam ram_block3a21.port_a_data_width = 1;
defparam ram_block3a21.port_a_first_address = 0;
defparam ram_block3a21.port_a_first_bit_number = 21;
defparam ram_block3a21.port_a_last_address = 8191;
defparam ram_block3a21.port_a_logical_ram_depth = 16384;
defparam ram_block3a21.port_a_logical_ram_width = 32;
defparam ram_block3a21.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block3a21.port_b_address_clear = "none";
defparam ram_block3a21.port_b_address_clock = "clock1";
defparam ram_block3a21.port_b_address_width = 13;
defparam ram_block3a21.port_b_data_in_clock = "clock1";
defparam ram_block3a21.port_b_data_out_clear = "none";
defparam ram_block3a21.port_b_data_out_clock = "none";
defparam ram_block3a21.port_b_data_width = 1;
defparam ram_block3a21.port_b_first_address = 0;
defparam ram_block3a21.port_b_first_bit_number = 21;
defparam ram_block3a21.port_b_last_address = 8191;
defparam ram_block3a21.port_b_logical_ram_depth = 16384;
defparam ram_block3a21.port_b_logical_ram_width = 32;
defparam ram_block3a21.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block3a21.port_b_read_enable_clock = "clock1";
defparam ram_block3a21.port_b_write_enable_clock = "clock1";
defparam ram_block3a21.ram_block_type = "M9K";
defparam ram_block3a21.mem_init3 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a21.mem_init2 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a21.mem_init1 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a21.mem_init0 = 2048'h0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000002A142119BCBBAB600000;
// synopsys translate_on

// Location: M9K_X78_Y35_N0
cycloneive_ram_block ram_block3a54(
	.portawe(\decode4|eq_node[1]~0_combout ),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(\decode5|eq_node[1]~0_combout ),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock1),
	.ena0(!ramaddr),
	.ena1(ram_rom_addr_reg_13),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({data_a[22]}),
	.portaaddr({address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain({data_b[22]}),
	.portbaddr({address_b[12],address_b[11],address_b[10],address_b[9],address_b[8],address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.devclrn(devclrn),
	.devpor(devpor),
	.portadataout(ram_block3a54_PORTADATAOUT_bus),
	.portbdataout(ram_block3a54_PORTBDATAOUT_bus));
// synopsys translate_off
defparam ram_block3a54.clk0_core_clock_enable = "ena0";
defparam ram_block3a54.clk1_core_clock_enable = "ena1";
defparam ram_block3a54.data_interleave_offset_in_bits = 1;
defparam ram_block3a54.data_interleave_width_in_bits = 1;
defparam ram_block3a54.init_file = "meminit.hex";
defparam ram_block3a54.init_file_layout = "port_a";
defparam ram_block3a54.logical_ram_name = "ram:RAM|altsyncram:altsyncram_component|altsyncram_99f1:auto_generated|altsyncram_fta2:altsyncram1|ALTSYNCRAM";
defparam ram_block3a54.mixed_port_feed_through_mode = "dont_care";
defparam ram_block3a54.operation_mode = "bidir_dual_port";
defparam ram_block3a54.port_a_address_clear = "none";
defparam ram_block3a54.port_a_address_width = 13;
defparam ram_block3a54.port_a_byte_enable_clock = "none";
defparam ram_block3a54.port_a_data_out_clear = "none";
defparam ram_block3a54.port_a_data_out_clock = "none";
defparam ram_block3a54.port_a_data_width = 1;
defparam ram_block3a54.port_a_first_address = 0;
defparam ram_block3a54.port_a_first_bit_number = 22;
defparam ram_block3a54.port_a_last_address = 8191;
defparam ram_block3a54.port_a_logical_ram_depth = 16384;
defparam ram_block3a54.port_a_logical_ram_width = 32;
defparam ram_block3a54.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block3a54.port_b_address_clear = "none";
defparam ram_block3a54.port_b_address_clock = "clock1";
defparam ram_block3a54.port_b_address_width = 13;
defparam ram_block3a54.port_b_data_in_clock = "clock1";
defparam ram_block3a54.port_b_data_out_clear = "none";
defparam ram_block3a54.port_b_data_out_clock = "none";
defparam ram_block3a54.port_b_data_width = 1;
defparam ram_block3a54.port_b_first_address = 0;
defparam ram_block3a54.port_b_first_bit_number = 22;
defparam ram_block3a54.port_b_last_address = 8191;
defparam ram_block3a54.port_b_logical_ram_depth = 16384;
defparam ram_block3a54.port_b_logical_ram_width = 32;
defparam ram_block3a54.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block3a54.port_b_read_enable_clock = "clock1";
defparam ram_block3a54.port_b_write_enable_clock = "clock1";
defparam ram_block3a54.ram_block_type = "M9K";
defparam ram_block3a54.mem_init3 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a54.mem_init2 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a54.mem_init1 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a54.mem_init0 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
// synopsys translate_on

// Location: M9K_X78_Y36_N0
cycloneive_ram_block ram_block3a22(
	.portawe(\decode4|eq_node[0]~1_combout ),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(\decode5|eq_node[0]~1_combout ),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock1),
	.ena0(ramaddr),
	.ena1(!ram_rom_addr_reg_13),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({data_a[22]}),
	.portaaddr({address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain({data_b[22]}),
	.portbaddr({address_b[12],address_b[11],address_b[10],address_b[9],address_b[8],address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.devclrn(devclrn),
	.devpor(devpor),
	.portadataout(ram_block3a22_PORTADATAOUT_bus),
	.portbdataout(ram_block3a22_PORTBDATAOUT_bus));
// synopsys translate_off
defparam ram_block3a22.clk0_core_clock_enable = "ena0";
defparam ram_block3a22.clk1_core_clock_enable = "ena1";
defparam ram_block3a22.data_interleave_offset_in_bits = 1;
defparam ram_block3a22.data_interleave_width_in_bits = 1;
defparam ram_block3a22.init_file = "meminit.hex";
defparam ram_block3a22.init_file_layout = "port_a";
defparam ram_block3a22.logical_ram_name = "ram:RAM|altsyncram:altsyncram_component|altsyncram_99f1:auto_generated|altsyncram_fta2:altsyncram1|ALTSYNCRAM";
defparam ram_block3a22.mixed_port_feed_through_mode = "dont_care";
defparam ram_block3a22.operation_mode = "bidir_dual_port";
defparam ram_block3a22.port_a_address_clear = "none";
defparam ram_block3a22.port_a_address_width = 13;
defparam ram_block3a22.port_a_byte_enable_clock = "none";
defparam ram_block3a22.port_a_data_out_clear = "none";
defparam ram_block3a22.port_a_data_out_clock = "none";
defparam ram_block3a22.port_a_data_width = 1;
defparam ram_block3a22.port_a_first_address = 0;
defparam ram_block3a22.port_a_first_bit_number = 22;
defparam ram_block3a22.port_a_last_address = 8191;
defparam ram_block3a22.port_a_logical_ram_depth = 16384;
defparam ram_block3a22.port_a_logical_ram_width = 32;
defparam ram_block3a22.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block3a22.port_b_address_clear = "none";
defparam ram_block3a22.port_b_address_clock = "clock1";
defparam ram_block3a22.port_b_address_width = 13;
defparam ram_block3a22.port_b_data_in_clock = "clock1";
defparam ram_block3a22.port_b_data_out_clear = "none";
defparam ram_block3a22.port_b_data_out_clock = "none";
defparam ram_block3a22.port_b_data_width = 1;
defparam ram_block3a22.port_b_first_address = 0;
defparam ram_block3a22.port_b_first_bit_number = 22;
defparam ram_block3a22.port_b_last_address = 8191;
defparam ram_block3a22.port_b_logical_ram_depth = 16384;
defparam ram_block3a22.port_b_logical_ram_width = 32;
defparam ram_block3a22.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block3a22.port_b_read_enable_clock = "clock1";
defparam ram_block3a22.port_b_write_enable_clock = "clock1";
defparam ram_block3a22.ram_block_type = "M9K";
defparam ram_block3a22.mem_init3 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a22.mem_init2 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a22.mem_init1 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a22.mem_init0 = 2048'h0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000002E403004A40002000000;
// synopsys translate_on

// Location: M9K_X64_Y23_N0
cycloneive_ram_block ram_block3a55(
	.portawe(\decode4|eq_node[1]~0_combout ),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(\decode5|eq_node[1]~0_combout ),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock1),
	.ena0(!ramaddr),
	.ena1(ram_rom_addr_reg_13),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({data_a[23]}),
	.portaaddr({address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain({data_b[23]}),
	.portbaddr({address_b[12],address_b[11],address_b[10],address_b[9],address_b[8],address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.devclrn(devclrn),
	.devpor(devpor),
	.portadataout(ram_block3a55_PORTADATAOUT_bus),
	.portbdataout(ram_block3a55_PORTBDATAOUT_bus));
// synopsys translate_off
defparam ram_block3a55.clk0_core_clock_enable = "ena0";
defparam ram_block3a55.clk1_core_clock_enable = "ena1";
defparam ram_block3a55.data_interleave_offset_in_bits = 1;
defparam ram_block3a55.data_interleave_width_in_bits = 1;
defparam ram_block3a55.init_file = "meminit.hex";
defparam ram_block3a55.init_file_layout = "port_a";
defparam ram_block3a55.logical_ram_name = "ram:RAM|altsyncram:altsyncram_component|altsyncram_99f1:auto_generated|altsyncram_fta2:altsyncram1|ALTSYNCRAM";
defparam ram_block3a55.mixed_port_feed_through_mode = "dont_care";
defparam ram_block3a55.operation_mode = "bidir_dual_port";
defparam ram_block3a55.port_a_address_clear = "none";
defparam ram_block3a55.port_a_address_width = 13;
defparam ram_block3a55.port_a_byte_enable_clock = "none";
defparam ram_block3a55.port_a_data_out_clear = "none";
defparam ram_block3a55.port_a_data_out_clock = "none";
defparam ram_block3a55.port_a_data_width = 1;
defparam ram_block3a55.port_a_first_address = 0;
defparam ram_block3a55.port_a_first_bit_number = 23;
defparam ram_block3a55.port_a_last_address = 8191;
defparam ram_block3a55.port_a_logical_ram_depth = 16384;
defparam ram_block3a55.port_a_logical_ram_width = 32;
defparam ram_block3a55.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block3a55.port_b_address_clear = "none";
defparam ram_block3a55.port_b_address_clock = "clock1";
defparam ram_block3a55.port_b_address_width = 13;
defparam ram_block3a55.port_b_data_in_clock = "clock1";
defparam ram_block3a55.port_b_data_out_clear = "none";
defparam ram_block3a55.port_b_data_out_clock = "none";
defparam ram_block3a55.port_b_data_width = 1;
defparam ram_block3a55.port_b_first_address = 0;
defparam ram_block3a55.port_b_first_bit_number = 23;
defparam ram_block3a55.port_b_last_address = 8191;
defparam ram_block3a55.port_b_logical_ram_depth = 16384;
defparam ram_block3a55.port_b_logical_ram_width = 32;
defparam ram_block3a55.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block3a55.port_b_read_enable_clock = "clock1";
defparam ram_block3a55.port_b_write_enable_clock = "clock1";
defparam ram_block3a55.ram_block_type = "M9K";
defparam ram_block3a55.mem_init3 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a55.mem_init2 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a55.mem_init1 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a55.mem_init0 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
// synopsys translate_on

// Location: M9K_X64_Y28_N0
cycloneive_ram_block ram_block3a23(
	.portawe(\decode4|eq_node[0]~1_combout ),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(\decode5|eq_node[0]~1_combout ),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock1),
	.ena0(ramaddr),
	.ena1(!ram_rom_addr_reg_13),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({data_a[23]}),
	.portaaddr({address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain({data_b[23]}),
	.portbaddr({address_b[12],address_b[11],address_b[10],address_b[9],address_b[8],address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.devclrn(devclrn),
	.devpor(devpor),
	.portadataout(ram_block3a23_PORTADATAOUT_bus),
	.portbdataout(ram_block3a23_PORTBDATAOUT_bus));
// synopsys translate_off
defparam ram_block3a23.clk0_core_clock_enable = "ena0";
defparam ram_block3a23.clk1_core_clock_enable = "ena1";
defparam ram_block3a23.data_interleave_offset_in_bits = 1;
defparam ram_block3a23.data_interleave_width_in_bits = 1;
defparam ram_block3a23.init_file = "meminit.hex";
defparam ram_block3a23.init_file_layout = "port_a";
defparam ram_block3a23.logical_ram_name = "ram:RAM|altsyncram:altsyncram_component|altsyncram_99f1:auto_generated|altsyncram_fta2:altsyncram1|ALTSYNCRAM";
defparam ram_block3a23.mixed_port_feed_through_mode = "dont_care";
defparam ram_block3a23.operation_mode = "bidir_dual_port";
defparam ram_block3a23.port_a_address_clear = "none";
defparam ram_block3a23.port_a_address_width = 13;
defparam ram_block3a23.port_a_byte_enable_clock = "none";
defparam ram_block3a23.port_a_data_out_clear = "none";
defparam ram_block3a23.port_a_data_out_clock = "none";
defparam ram_block3a23.port_a_data_width = 1;
defparam ram_block3a23.port_a_first_address = 0;
defparam ram_block3a23.port_a_first_bit_number = 23;
defparam ram_block3a23.port_a_last_address = 8191;
defparam ram_block3a23.port_a_logical_ram_depth = 16384;
defparam ram_block3a23.port_a_logical_ram_width = 32;
defparam ram_block3a23.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block3a23.port_b_address_clear = "none";
defparam ram_block3a23.port_b_address_clock = "clock1";
defparam ram_block3a23.port_b_address_width = 13;
defparam ram_block3a23.port_b_data_in_clock = "clock1";
defparam ram_block3a23.port_b_data_out_clear = "none";
defparam ram_block3a23.port_b_data_out_clock = "none";
defparam ram_block3a23.port_b_data_width = 1;
defparam ram_block3a23.port_b_first_address = 0;
defparam ram_block3a23.port_b_first_bit_number = 23;
defparam ram_block3a23.port_b_last_address = 8191;
defparam ram_block3a23.port_b_logical_ram_depth = 16384;
defparam ram_block3a23.port_b_logical_ram_width = 32;
defparam ram_block3a23.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block3a23.port_b_read_enable_clock = "clock1";
defparam ram_block3a23.port_b_write_enable_clock = "clock1";
defparam ram_block3a23.ram_block_type = "M9K";
defparam ram_block3a23.mem_init3 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a23.mem_init2 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a23.mem_init1 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a23.mem_init0 = 2048'h0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000002E5CB187BC004B601000;
// synopsys translate_on

// Location: M9K_X64_Y31_N0
cycloneive_ram_block ram_block3a56(
	.portawe(\decode4|eq_node[1]~0_combout ),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(\decode5|eq_node[1]~0_combout ),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock1),
	.ena0(!ramaddr),
	.ena1(ram_rom_addr_reg_13),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({data_a[24]}),
	.portaaddr({address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain({data_b[24]}),
	.portbaddr({address_b[12],address_b[11],address_b[10],address_b[9],address_b[8],address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.devclrn(devclrn),
	.devpor(devpor),
	.portadataout(ram_block3a56_PORTADATAOUT_bus),
	.portbdataout(ram_block3a56_PORTBDATAOUT_bus));
// synopsys translate_off
defparam ram_block3a56.clk0_core_clock_enable = "ena0";
defparam ram_block3a56.clk1_core_clock_enable = "ena1";
defparam ram_block3a56.data_interleave_offset_in_bits = 1;
defparam ram_block3a56.data_interleave_width_in_bits = 1;
defparam ram_block3a56.init_file = "meminit.hex";
defparam ram_block3a56.init_file_layout = "port_a";
defparam ram_block3a56.logical_ram_name = "ram:RAM|altsyncram:altsyncram_component|altsyncram_99f1:auto_generated|altsyncram_fta2:altsyncram1|ALTSYNCRAM";
defparam ram_block3a56.mixed_port_feed_through_mode = "dont_care";
defparam ram_block3a56.operation_mode = "bidir_dual_port";
defparam ram_block3a56.port_a_address_clear = "none";
defparam ram_block3a56.port_a_address_width = 13;
defparam ram_block3a56.port_a_byte_enable_clock = "none";
defparam ram_block3a56.port_a_data_out_clear = "none";
defparam ram_block3a56.port_a_data_out_clock = "none";
defparam ram_block3a56.port_a_data_width = 1;
defparam ram_block3a56.port_a_first_address = 0;
defparam ram_block3a56.port_a_first_bit_number = 24;
defparam ram_block3a56.port_a_last_address = 8191;
defparam ram_block3a56.port_a_logical_ram_depth = 16384;
defparam ram_block3a56.port_a_logical_ram_width = 32;
defparam ram_block3a56.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block3a56.port_b_address_clear = "none";
defparam ram_block3a56.port_b_address_clock = "clock1";
defparam ram_block3a56.port_b_address_width = 13;
defparam ram_block3a56.port_b_data_in_clock = "clock1";
defparam ram_block3a56.port_b_data_out_clear = "none";
defparam ram_block3a56.port_b_data_out_clock = "none";
defparam ram_block3a56.port_b_data_width = 1;
defparam ram_block3a56.port_b_first_address = 0;
defparam ram_block3a56.port_b_first_bit_number = 24;
defparam ram_block3a56.port_b_last_address = 8191;
defparam ram_block3a56.port_b_logical_ram_depth = 16384;
defparam ram_block3a56.port_b_logical_ram_width = 32;
defparam ram_block3a56.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block3a56.port_b_read_enable_clock = "clock1";
defparam ram_block3a56.port_b_write_enable_clock = "clock1";
defparam ram_block3a56.ram_block_type = "M9K";
defparam ram_block3a56.mem_init3 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a56.mem_init2 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a56.mem_init1 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a56.mem_init0 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
// synopsys translate_on

// Location: M9K_X64_Y32_N0
cycloneive_ram_block ram_block3a24(
	.portawe(\decode4|eq_node[0]~1_combout ),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(\decode5|eq_node[0]~1_combout ),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock1),
	.ena0(ramaddr),
	.ena1(!ram_rom_addr_reg_13),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({data_a[24]}),
	.portaaddr({address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain({data_b[24]}),
	.portbaddr({address_b[12],address_b[11],address_b[10],address_b[9],address_b[8],address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.devclrn(devclrn),
	.devpor(devpor),
	.portadataout(ram_block3a24_PORTADATAOUT_bus),
	.portbdataout(ram_block3a24_PORTBDATAOUT_bus));
// synopsys translate_off
defparam ram_block3a24.clk0_core_clock_enable = "ena0";
defparam ram_block3a24.clk1_core_clock_enable = "ena1";
defparam ram_block3a24.data_interleave_offset_in_bits = 1;
defparam ram_block3a24.data_interleave_width_in_bits = 1;
defparam ram_block3a24.init_file = "meminit.hex";
defparam ram_block3a24.init_file_layout = "port_a";
defparam ram_block3a24.logical_ram_name = "ram:RAM|altsyncram:altsyncram_component|altsyncram_99f1:auto_generated|altsyncram_fta2:altsyncram1|ALTSYNCRAM";
defparam ram_block3a24.mixed_port_feed_through_mode = "dont_care";
defparam ram_block3a24.operation_mode = "bidir_dual_port";
defparam ram_block3a24.port_a_address_clear = "none";
defparam ram_block3a24.port_a_address_width = 13;
defparam ram_block3a24.port_a_byte_enable_clock = "none";
defparam ram_block3a24.port_a_data_out_clear = "none";
defparam ram_block3a24.port_a_data_out_clock = "none";
defparam ram_block3a24.port_a_data_width = 1;
defparam ram_block3a24.port_a_first_address = 0;
defparam ram_block3a24.port_a_first_bit_number = 24;
defparam ram_block3a24.port_a_last_address = 8191;
defparam ram_block3a24.port_a_logical_ram_depth = 16384;
defparam ram_block3a24.port_a_logical_ram_width = 32;
defparam ram_block3a24.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block3a24.port_b_address_clear = "none";
defparam ram_block3a24.port_b_address_clock = "clock1";
defparam ram_block3a24.port_b_address_width = 13;
defparam ram_block3a24.port_b_data_in_clock = "clock1";
defparam ram_block3a24.port_b_data_out_clear = "none";
defparam ram_block3a24.port_b_data_out_clock = "none";
defparam ram_block3a24.port_b_data_width = 1;
defparam ram_block3a24.port_b_first_address = 0;
defparam ram_block3a24.port_b_first_bit_number = 24;
defparam ram_block3a24.port_b_last_address = 8191;
defparam ram_block3a24.port_b_logical_ram_depth = 16384;
defparam ram_block3a24.port_b_logical_ram_width = 32;
defparam ram_block3a24.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block3a24.port_b_read_enable_clock = "clock1";
defparam ram_block3a24.port_b_write_enable_clock = "clock1";
defparam ram_block3a24.ram_block_type = "M9K";
defparam ram_block3a24.mem_init3 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a24.mem_init2 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a24.mem_init1 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a24.mem_init0 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000021830C680DB793600400;
// synopsys translate_on

// Location: M9K_X78_Y34_N0
cycloneive_ram_block ram_block3a57(
	.portawe(\decode4|eq_node[1]~0_combout ),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(\decode5|eq_node[1]~0_combout ),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock1),
	.ena0(!ramaddr),
	.ena1(ram_rom_addr_reg_13),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({data_a[25]}),
	.portaaddr({address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain({data_b[25]}),
	.portbaddr({address_b[12],address_b[11],address_b[10],address_b[9],address_b[8],address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.devclrn(devclrn),
	.devpor(devpor),
	.portadataout(ram_block3a57_PORTADATAOUT_bus),
	.portbdataout(ram_block3a57_PORTBDATAOUT_bus));
// synopsys translate_off
defparam ram_block3a57.clk0_core_clock_enable = "ena0";
defparam ram_block3a57.clk1_core_clock_enable = "ena1";
defparam ram_block3a57.data_interleave_offset_in_bits = 1;
defparam ram_block3a57.data_interleave_width_in_bits = 1;
defparam ram_block3a57.init_file = "meminit.hex";
defparam ram_block3a57.init_file_layout = "port_a";
defparam ram_block3a57.logical_ram_name = "ram:RAM|altsyncram:altsyncram_component|altsyncram_99f1:auto_generated|altsyncram_fta2:altsyncram1|ALTSYNCRAM";
defparam ram_block3a57.mixed_port_feed_through_mode = "dont_care";
defparam ram_block3a57.operation_mode = "bidir_dual_port";
defparam ram_block3a57.port_a_address_clear = "none";
defparam ram_block3a57.port_a_address_width = 13;
defparam ram_block3a57.port_a_byte_enable_clock = "none";
defparam ram_block3a57.port_a_data_out_clear = "none";
defparam ram_block3a57.port_a_data_out_clock = "none";
defparam ram_block3a57.port_a_data_width = 1;
defparam ram_block3a57.port_a_first_address = 0;
defparam ram_block3a57.port_a_first_bit_number = 25;
defparam ram_block3a57.port_a_last_address = 8191;
defparam ram_block3a57.port_a_logical_ram_depth = 16384;
defparam ram_block3a57.port_a_logical_ram_width = 32;
defparam ram_block3a57.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block3a57.port_b_address_clear = "none";
defparam ram_block3a57.port_b_address_clock = "clock1";
defparam ram_block3a57.port_b_address_width = 13;
defparam ram_block3a57.port_b_data_in_clock = "clock1";
defparam ram_block3a57.port_b_data_out_clear = "none";
defparam ram_block3a57.port_b_data_out_clock = "none";
defparam ram_block3a57.port_b_data_width = 1;
defparam ram_block3a57.port_b_first_address = 0;
defparam ram_block3a57.port_b_first_bit_number = 25;
defparam ram_block3a57.port_b_last_address = 8191;
defparam ram_block3a57.port_b_logical_ram_depth = 16384;
defparam ram_block3a57.port_b_logical_ram_width = 32;
defparam ram_block3a57.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block3a57.port_b_read_enable_clock = "clock1";
defparam ram_block3a57.port_b_write_enable_clock = "clock1";
defparam ram_block3a57.ram_block_type = "M9K";
defparam ram_block3a57.mem_init3 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a57.mem_init2 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a57.mem_init1 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a57.mem_init0 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
// synopsys translate_on

// Location: M9K_X78_Y33_N0
cycloneive_ram_block ram_block3a25(
	.portawe(\decode4|eq_node[0]~1_combout ),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(\decode5|eq_node[0]~1_combout ),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock1),
	.ena0(ramaddr),
	.ena1(!ram_rom_addr_reg_13),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({data_a[25]}),
	.portaaddr({address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain({data_b[25]}),
	.portbaddr({address_b[12],address_b[11],address_b[10],address_b[9],address_b[8],address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.devclrn(devclrn),
	.devpor(devpor),
	.portadataout(ram_block3a25_PORTADATAOUT_bus),
	.portbdataout(ram_block3a25_PORTBDATAOUT_bus));
// synopsys translate_off
defparam ram_block3a25.clk0_core_clock_enable = "ena0";
defparam ram_block3a25.clk1_core_clock_enable = "ena1";
defparam ram_block3a25.data_interleave_offset_in_bits = 1;
defparam ram_block3a25.data_interleave_width_in_bits = 1;
defparam ram_block3a25.init_file = "meminit.hex";
defparam ram_block3a25.init_file_layout = "port_a";
defparam ram_block3a25.logical_ram_name = "ram:RAM|altsyncram:altsyncram_component|altsyncram_99f1:auto_generated|altsyncram_fta2:altsyncram1|ALTSYNCRAM";
defparam ram_block3a25.mixed_port_feed_through_mode = "dont_care";
defparam ram_block3a25.operation_mode = "bidir_dual_port";
defparam ram_block3a25.port_a_address_clear = "none";
defparam ram_block3a25.port_a_address_width = 13;
defparam ram_block3a25.port_a_byte_enable_clock = "none";
defparam ram_block3a25.port_a_data_out_clear = "none";
defparam ram_block3a25.port_a_data_out_clock = "none";
defparam ram_block3a25.port_a_data_width = 1;
defparam ram_block3a25.port_a_first_address = 0;
defparam ram_block3a25.port_a_first_bit_number = 25;
defparam ram_block3a25.port_a_last_address = 8191;
defparam ram_block3a25.port_a_logical_ram_depth = 16384;
defparam ram_block3a25.port_a_logical_ram_width = 32;
defparam ram_block3a25.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block3a25.port_b_address_clear = "none";
defparam ram_block3a25.port_b_address_clock = "clock1";
defparam ram_block3a25.port_b_address_width = 13;
defparam ram_block3a25.port_b_data_in_clock = "clock1";
defparam ram_block3a25.port_b_data_out_clear = "none";
defparam ram_block3a25.port_b_data_out_clock = "none";
defparam ram_block3a25.port_b_data_width = 1;
defparam ram_block3a25.port_b_first_address = 0;
defparam ram_block3a25.port_b_first_bit_number = 25;
defparam ram_block3a25.port_b_last_address = 8191;
defparam ram_block3a25.port_b_logical_ram_depth = 16384;
defparam ram_block3a25.port_b_logical_ram_width = 32;
defparam ram_block3a25.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block3a25.port_b_read_enable_clock = "clock1";
defparam ram_block3a25.port_b_write_enable_clock = "clock1";
defparam ram_block3a25.ram_block_type = "M9K";
defparam ram_block3a25.mem_init3 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a25.mem_init2 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a25.mem_init1 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a25.mem_init0 = 2048'h000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000200000000CB783600310;
// synopsys translate_on

// Location: M9K_X78_Y26_N0
cycloneive_ram_block ram_block3a58(
	.portawe(\decode4|eq_node[1]~0_combout ),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(\decode5|eq_node[1]~0_combout ),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock1),
	.ena0(!ramaddr),
	.ena1(ram_rom_addr_reg_13),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({data_a[26]}),
	.portaaddr({address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain({data_b[26]}),
	.portbaddr({address_b[12],address_b[11],address_b[10],address_b[9],address_b[8],address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.devclrn(devclrn),
	.devpor(devpor),
	.portadataout(ram_block3a58_PORTADATAOUT_bus),
	.portbdataout(ram_block3a58_PORTBDATAOUT_bus));
// synopsys translate_off
defparam ram_block3a58.clk0_core_clock_enable = "ena0";
defparam ram_block3a58.clk1_core_clock_enable = "ena1";
defparam ram_block3a58.data_interleave_offset_in_bits = 1;
defparam ram_block3a58.data_interleave_width_in_bits = 1;
defparam ram_block3a58.init_file = "meminit.hex";
defparam ram_block3a58.init_file_layout = "port_a";
defparam ram_block3a58.logical_ram_name = "ram:RAM|altsyncram:altsyncram_component|altsyncram_99f1:auto_generated|altsyncram_fta2:altsyncram1|ALTSYNCRAM";
defparam ram_block3a58.mixed_port_feed_through_mode = "dont_care";
defparam ram_block3a58.operation_mode = "bidir_dual_port";
defparam ram_block3a58.port_a_address_clear = "none";
defparam ram_block3a58.port_a_address_width = 13;
defparam ram_block3a58.port_a_byte_enable_clock = "none";
defparam ram_block3a58.port_a_data_out_clear = "none";
defparam ram_block3a58.port_a_data_out_clock = "none";
defparam ram_block3a58.port_a_data_width = 1;
defparam ram_block3a58.port_a_first_address = 0;
defparam ram_block3a58.port_a_first_bit_number = 26;
defparam ram_block3a58.port_a_last_address = 8191;
defparam ram_block3a58.port_a_logical_ram_depth = 16384;
defparam ram_block3a58.port_a_logical_ram_width = 32;
defparam ram_block3a58.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block3a58.port_b_address_clear = "none";
defparam ram_block3a58.port_b_address_clock = "clock1";
defparam ram_block3a58.port_b_address_width = 13;
defparam ram_block3a58.port_b_data_in_clock = "clock1";
defparam ram_block3a58.port_b_data_out_clear = "none";
defparam ram_block3a58.port_b_data_out_clock = "none";
defparam ram_block3a58.port_b_data_width = 1;
defparam ram_block3a58.port_b_first_address = 0;
defparam ram_block3a58.port_b_first_bit_number = 26;
defparam ram_block3a58.port_b_last_address = 8191;
defparam ram_block3a58.port_b_logical_ram_depth = 16384;
defparam ram_block3a58.port_b_logical_ram_width = 32;
defparam ram_block3a58.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block3a58.port_b_read_enable_clock = "clock1";
defparam ram_block3a58.port_b_write_enable_clock = "clock1";
defparam ram_block3a58.ram_block_type = "M9K";
defparam ram_block3a58.mem_init3 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a58.mem_init2 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a58.mem_init1 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a58.mem_init0 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
// synopsys translate_on

// Location: M9K_X78_Y25_N0
cycloneive_ram_block ram_block3a26(
	.portawe(\decode4|eq_node[0]~1_combout ),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(\decode5|eq_node[0]~1_combout ),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock1),
	.ena0(ramaddr),
	.ena1(!ram_rom_addr_reg_13),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({data_a[26]}),
	.portaaddr({address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain({data_b[26]}),
	.portbaddr({address_b[12],address_b[11],address_b[10],address_b[9],address_b[8],address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.devclrn(devclrn),
	.devpor(devpor),
	.portadataout(ram_block3a26_PORTADATAOUT_bus),
	.portbdataout(ram_block3a26_PORTBDATAOUT_bus));
// synopsys translate_off
defparam ram_block3a26.clk0_core_clock_enable = "ena0";
defparam ram_block3a26.clk1_core_clock_enable = "ena1";
defparam ram_block3a26.data_interleave_offset_in_bits = 1;
defparam ram_block3a26.data_interleave_width_in_bits = 1;
defparam ram_block3a26.init_file = "meminit.hex";
defparam ram_block3a26.init_file_layout = "port_a";
defparam ram_block3a26.logical_ram_name = "ram:RAM|altsyncram:altsyncram_component|altsyncram_99f1:auto_generated|altsyncram_fta2:altsyncram1|ALTSYNCRAM";
defparam ram_block3a26.mixed_port_feed_through_mode = "dont_care";
defparam ram_block3a26.operation_mode = "bidir_dual_port";
defparam ram_block3a26.port_a_address_clear = "none";
defparam ram_block3a26.port_a_address_width = 13;
defparam ram_block3a26.port_a_byte_enable_clock = "none";
defparam ram_block3a26.port_a_data_out_clear = "none";
defparam ram_block3a26.port_a_data_out_clock = "none";
defparam ram_block3a26.port_a_data_width = 1;
defparam ram_block3a26.port_a_first_address = 0;
defparam ram_block3a26.port_a_first_bit_number = 26;
defparam ram_block3a26.port_a_last_address = 8191;
defparam ram_block3a26.port_a_logical_ram_depth = 16384;
defparam ram_block3a26.port_a_logical_ram_width = 32;
defparam ram_block3a26.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block3a26.port_b_address_clear = "none";
defparam ram_block3a26.port_b_address_clock = "clock1";
defparam ram_block3a26.port_b_address_width = 13;
defparam ram_block3a26.port_b_data_in_clock = "clock1";
defparam ram_block3a26.port_b_data_out_clear = "none";
defparam ram_block3a26.port_b_data_out_clock = "none";
defparam ram_block3a26.port_b_data_width = 1;
defparam ram_block3a26.port_b_first_address = 0;
defparam ram_block3a26.port_b_first_bit_number = 26;
defparam ram_block3a26.port_b_last_address = 8191;
defparam ram_block3a26.port_b_logical_ram_depth = 16384;
defparam ram_block3a26.port_b_logical_ram_width = 32;
defparam ram_block3a26.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block3a26.port_b_read_enable_clock = "clock1";
defparam ram_block3a26.port_b_write_enable_clock = "clock1";
defparam ram_block3a26.ram_block_type = "M9K";
defparam ram_block3a26.mem_init3 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a26.mem_init2 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a26.mem_init1 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a26.mem_init0 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000007CFBDE639B287F0888F;
// synopsys translate_on

// Location: M9K_X78_Y31_N0
cycloneive_ram_block ram_block3a59(
	.portawe(\decode4|eq_node[1]~0_combout ),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(\decode5|eq_node[1]~0_combout ),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock1),
	.ena0(!ramaddr),
	.ena1(ram_rom_addr_reg_13),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({data_a[27]}),
	.portaaddr({address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain({data_b[27]}),
	.portbaddr({address_b[12],address_b[11],address_b[10],address_b[9],address_b[8],address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.devclrn(devclrn),
	.devpor(devpor),
	.portadataout(ram_block3a59_PORTADATAOUT_bus),
	.portbdataout(ram_block3a59_PORTBDATAOUT_bus));
// synopsys translate_off
defparam ram_block3a59.clk0_core_clock_enable = "ena0";
defparam ram_block3a59.clk1_core_clock_enable = "ena1";
defparam ram_block3a59.data_interleave_offset_in_bits = 1;
defparam ram_block3a59.data_interleave_width_in_bits = 1;
defparam ram_block3a59.init_file = "meminit.hex";
defparam ram_block3a59.init_file_layout = "port_a";
defparam ram_block3a59.logical_ram_name = "ram:RAM|altsyncram:altsyncram_component|altsyncram_99f1:auto_generated|altsyncram_fta2:altsyncram1|ALTSYNCRAM";
defparam ram_block3a59.mixed_port_feed_through_mode = "dont_care";
defparam ram_block3a59.operation_mode = "bidir_dual_port";
defparam ram_block3a59.port_a_address_clear = "none";
defparam ram_block3a59.port_a_address_width = 13;
defparam ram_block3a59.port_a_byte_enable_clock = "none";
defparam ram_block3a59.port_a_data_out_clear = "none";
defparam ram_block3a59.port_a_data_out_clock = "none";
defparam ram_block3a59.port_a_data_width = 1;
defparam ram_block3a59.port_a_first_address = 0;
defparam ram_block3a59.port_a_first_bit_number = 27;
defparam ram_block3a59.port_a_last_address = 8191;
defparam ram_block3a59.port_a_logical_ram_depth = 16384;
defparam ram_block3a59.port_a_logical_ram_width = 32;
defparam ram_block3a59.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block3a59.port_b_address_clear = "none";
defparam ram_block3a59.port_b_address_clock = "clock1";
defparam ram_block3a59.port_b_address_width = 13;
defparam ram_block3a59.port_b_data_in_clock = "clock1";
defparam ram_block3a59.port_b_data_out_clear = "none";
defparam ram_block3a59.port_b_data_out_clock = "none";
defparam ram_block3a59.port_b_data_width = 1;
defparam ram_block3a59.port_b_first_address = 0;
defparam ram_block3a59.port_b_first_bit_number = 27;
defparam ram_block3a59.port_b_last_address = 8191;
defparam ram_block3a59.port_b_logical_ram_depth = 16384;
defparam ram_block3a59.port_b_logical_ram_width = 32;
defparam ram_block3a59.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block3a59.port_b_read_enable_clock = "clock1";
defparam ram_block3a59.port_b_write_enable_clock = "clock1";
defparam ram_block3a59.ram_block_type = "M9K";
defparam ram_block3a59.mem_init3 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a59.mem_init2 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a59.mem_init1 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a59.mem_init0 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
// synopsys translate_on

// Location: M9K_X78_Y27_N0
cycloneive_ram_block ram_block3a27(
	.portawe(\decode4|eq_node[0]~1_combout ),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(\decode5|eq_node[0]~1_combout ),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock1),
	.ena0(ramaddr),
	.ena1(!ram_rom_addr_reg_13),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({data_a[27]}),
	.portaaddr({address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain({data_b[27]}),
	.portbaddr({address_b[12],address_b[11],address_b[10],address_b[9],address_b[8],address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.devclrn(devclrn),
	.devpor(devpor),
	.portadataout(ram_block3a27_PORTADATAOUT_bus),
	.portbdataout(ram_block3a27_PORTBDATAOUT_bus));
// synopsys translate_off
defparam ram_block3a27.clk0_core_clock_enable = "ena0";
defparam ram_block3a27.clk1_core_clock_enable = "ena1";
defparam ram_block3a27.data_interleave_offset_in_bits = 1;
defparam ram_block3a27.data_interleave_width_in_bits = 1;
defparam ram_block3a27.init_file = "meminit.hex";
defparam ram_block3a27.init_file_layout = "port_a";
defparam ram_block3a27.logical_ram_name = "ram:RAM|altsyncram:altsyncram_component|altsyncram_99f1:auto_generated|altsyncram_fta2:altsyncram1|ALTSYNCRAM";
defparam ram_block3a27.mixed_port_feed_through_mode = "dont_care";
defparam ram_block3a27.operation_mode = "bidir_dual_port";
defparam ram_block3a27.port_a_address_clear = "none";
defparam ram_block3a27.port_a_address_width = 13;
defparam ram_block3a27.port_a_byte_enable_clock = "none";
defparam ram_block3a27.port_a_data_out_clear = "none";
defparam ram_block3a27.port_a_data_out_clock = "none";
defparam ram_block3a27.port_a_data_width = 1;
defparam ram_block3a27.port_a_first_address = 0;
defparam ram_block3a27.port_a_first_bit_number = 27;
defparam ram_block3a27.port_a_last_address = 8191;
defparam ram_block3a27.port_a_logical_ram_depth = 16384;
defparam ram_block3a27.port_a_logical_ram_width = 32;
defparam ram_block3a27.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block3a27.port_b_address_clear = "none";
defparam ram_block3a27.port_b_address_clock = "clock1";
defparam ram_block3a27.port_b_address_width = 13;
defparam ram_block3a27.port_b_data_in_clock = "clock1";
defparam ram_block3a27.port_b_data_out_clear = "none";
defparam ram_block3a27.port_b_data_out_clock = "none";
defparam ram_block3a27.port_b_data_width = 1;
defparam ram_block3a27.port_b_first_address = 0;
defparam ram_block3a27.port_b_first_bit_number = 27;
defparam ram_block3a27.port_b_last_address = 8191;
defparam ram_block3a27.port_b_logical_ram_depth = 16384;
defparam ram_block3a27.port_b_logical_ram_width = 32;
defparam ram_block3a27.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block3a27.port_b_read_enable_clock = "clock1";
defparam ram_block3a27.port_b_write_enable_clock = "clock1";
defparam ram_block3a27.ram_block_type = "M9K";
defparam ram_block3a27.mem_init3 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a27.mem_init2 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a27.mem_init1 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a27.mem_init0 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010E1C6264AD282C08088;
// synopsys translate_on

// Location: M9K_X78_Y30_N0
cycloneive_ram_block ram_block3a60(
	.portawe(\decode4|eq_node[1]~0_combout ),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(\decode5|eq_node[1]~0_combout ),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock1),
	.ena0(!ramaddr),
	.ena1(ram_rom_addr_reg_13),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({data_a[28]}),
	.portaaddr({address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain({data_b[28]}),
	.portbaddr({address_b[12],address_b[11],address_b[10],address_b[9],address_b[8],address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.devclrn(devclrn),
	.devpor(devpor),
	.portadataout(ram_block3a60_PORTADATAOUT_bus),
	.portbdataout(ram_block3a60_PORTBDATAOUT_bus));
// synopsys translate_off
defparam ram_block3a60.clk0_core_clock_enable = "ena0";
defparam ram_block3a60.clk1_core_clock_enable = "ena1";
defparam ram_block3a60.data_interleave_offset_in_bits = 1;
defparam ram_block3a60.data_interleave_width_in_bits = 1;
defparam ram_block3a60.init_file = "meminit.hex";
defparam ram_block3a60.init_file_layout = "port_a";
defparam ram_block3a60.logical_ram_name = "ram:RAM|altsyncram:altsyncram_component|altsyncram_99f1:auto_generated|altsyncram_fta2:altsyncram1|ALTSYNCRAM";
defparam ram_block3a60.mixed_port_feed_through_mode = "dont_care";
defparam ram_block3a60.operation_mode = "bidir_dual_port";
defparam ram_block3a60.port_a_address_clear = "none";
defparam ram_block3a60.port_a_address_width = 13;
defparam ram_block3a60.port_a_byte_enable_clock = "none";
defparam ram_block3a60.port_a_data_out_clear = "none";
defparam ram_block3a60.port_a_data_out_clock = "none";
defparam ram_block3a60.port_a_data_width = 1;
defparam ram_block3a60.port_a_first_address = 0;
defparam ram_block3a60.port_a_first_bit_number = 28;
defparam ram_block3a60.port_a_last_address = 8191;
defparam ram_block3a60.port_a_logical_ram_depth = 16384;
defparam ram_block3a60.port_a_logical_ram_width = 32;
defparam ram_block3a60.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block3a60.port_b_address_clear = "none";
defparam ram_block3a60.port_b_address_clock = "clock1";
defparam ram_block3a60.port_b_address_width = 13;
defparam ram_block3a60.port_b_data_in_clock = "clock1";
defparam ram_block3a60.port_b_data_out_clear = "none";
defparam ram_block3a60.port_b_data_out_clock = "none";
defparam ram_block3a60.port_b_data_width = 1;
defparam ram_block3a60.port_b_first_address = 0;
defparam ram_block3a60.port_b_first_bit_number = 28;
defparam ram_block3a60.port_b_last_address = 8191;
defparam ram_block3a60.port_b_logical_ram_depth = 16384;
defparam ram_block3a60.port_b_logical_ram_width = 32;
defparam ram_block3a60.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block3a60.port_b_read_enable_clock = "clock1";
defparam ram_block3a60.port_b_write_enable_clock = "clock1";
defparam ram_block3a60.ram_block_type = "M9K";
defparam ram_block3a60.mem_init3 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a60.mem_init2 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a60.mem_init1 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a60.mem_init0 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
// synopsys translate_on

// Location: M9K_X78_Y29_N0
cycloneive_ram_block ram_block3a28(
	.portawe(\decode4|eq_node[0]~1_combout ),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(\decode5|eq_node[0]~1_combout ),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock1),
	.ena0(ramaddr),
	.ena1(!ram_rom_addr_reg_13),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({data_a[28]}),
	.portaaddr({address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain({data_b[28]}),
	.portbaddr({address_b[12],address_b[11],address_b[10],address_b[9],address_b[8],address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.devclrn(devclrn),
	.devpor(devpor),
	.portadataout(ram_block3a28_PORTADATAOUT_bus),
	.portbdataout(ram_block3a28_PORTBDATAOUT_bus));
// synopsys translate_off
defparam ram_block3a28.clk0_core_clock_enable = "ena0";
defparam ram_block3a28.clk1_core_clock_enable = "ena1";
defparam ram_block3a28.data_interleave_offset_in_bits = 1;
defparam ram_block3a28.data_interleave_width_in_bits = 1;
defparam ram_block3a28.init_file = "meminit.hex";
defparam ram_block3a28.init_file_layout = "port_a";
defparam ram_block3a28.logical_ram_name = "ram:RAM|altsyncram:altsyncram_component|altsyncram_99f1:auto_generated|altsyncram_fta2:altsyncram1|ALTSYNCRAM";
defparam ram_block3a28.mixed_port_feed_through_mode = "dont_care";
defparam ram_block3a28.operation_mode = "bidir_dual_port";
defparam ram_block3a28.port_a_address_clear = "none";
defparam ram_block3a28.port_a_address_width = 13;
defparam ram_block3a28.port_a_byte_enable_clock = "none";
defparam ram_block3a28.port_a_data_out_clear = "none";
defparam ram_block3a28.port_a_data_out_clock = "none";
defparam ram_block3a28.port_a_data_width = 1;
defparam ram_block3a28.port_a_first_address = 0;
defparam ram_block3a28.port_a_first_bit_number = 28;
defparam ram_block3a28.port_a_last_address = 8191;
defparam ram_block3a28.port_a_logical_ram_depth = 16384;
defparam ram_block3a28.port_a_logical_ram_width = 32;
defparam ram_block3a28.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block3a28.port_b_address_clear = "none";
defparam ram_block3a28.port_b_address_clock = "clock1";
defparam ram_block3a28.port_b_address_width = 13;
defparam ram_block3a28.port_b_data_in_clock = "clock1";
defparam ram_block3a28.port_b_data_out_clear = "none";
defparam ram_block3a28.port_b_data_out_clock = "none";
defparam ram_block3a28.port_b_data_width = 1;
defparam ram_block3a28.port_b_first_address = 0;
defparam ram_block3a28.port_b_first_bit_number = 28;
defparam ram_block3a28.port_b_last_address = 8191;
defparam ram_block3a28.port_b_logical_ram_depth = 16384;
defparam ram_block3a28.port_b_logical_ram_width = 32;
defparam ram_block3a28.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block3a28.port_b_read_enable_clock = "clock1";
defparam ram_block3a28.port_b_write_enable_clock = "clock1";
defparam ram_block3a28.ram_block_type = "M9K";
defparam ram_block3a28.mem_init3 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a28.mem_init2 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a28.mem_init1 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a28.mem_init0 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000008100011B00926100807;
// synopsys translate_on

// Location: M9K_X78_Y37_N0
cycloneive_ram_block ram_block3a61(
	.portawe(\decode4|eq_node[1]~0_combout ),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(\decode5|eq_node[1]~0_combout ),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock1),
	.ena0(!ramaddr),
	.ena1(ram_rom_addr_reg_13),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({data_a[29]}),
	.portaaddr({address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain({data_b[29]}),
	.portbaddr({address_b[12],address_b[11],address_b[10],address_b[9],address_b[8],address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.devclrn(devclrn),
	.devpor(devpor),
	.portadataout(ram_block3a61_PORTADATAOUT_bus),
	.portbdataout(ram_block3a61_PORTBDATAOUT_bus));
// synopsys translate_off
defparam ram_block3a61.clk0_core_clock_enable = "ena0";
defparam ram_block3a61.clk1_core_clock_enable = "ena1";
defparam ram_block3a61.data_interleave_offset_in_bits = 1;
defparam ram_block3a61.data_interleave_width_in_bits = 1;
defparam ram_block3a61.init_file = "meminit.hex";
defparam ram_block3a61.init_file_layout = "port_a";
defparam ram_block3a61.logical_ram_name = "ram:RAM|altsyncram:altsyncram_component|altsyncram_99f1:auto_generated|altsyncram_fta2:altsyncram1|ALTSYNCRAM";
defparam ram_block3a61.mixed_port_feed_through_mode = "dont_care";
defparam ram_block3a61.operation_mode = "bidir_dual_port";
defparam ram_block3a61.port_a_address_clear = "none";
defparam ram_block3a61.port_a_address_width = 13;
defparam ram_block3a61.port_a_byte_enable_clock = "none";
defparam ram_block3a61.port_a_data_out_clear = "none";
defparam ram_block3a61.port_a_data_out_clock = "none";
defparam ram_block3a61.port_a_data_width = 1;
defparam ram_block3a61.port_a_first_address = 0;
defparam ram_block3a61.port_a_first_bit_number = 29;
defparam ram_block3a61.port_a_last_address = 8191;
defparam ram_block3a61.port_a_logical_ram_depth = 16384;
defparam ram_block3a61.port_a_logical_ram_width = 32;
defparam ram_block3a61.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block3a61.port_b_address_clear = "none";
defparam ram_block3a61.port_b_address_clock = "clock1";
defparam ram_block3a61.port_b_address_width = 13;
defparam ram_block3a61.port_b_data_in_clock = "clock1";
defparam ram_block3a61.port_b_data_out_clear = "none";
defparam ram_block3a61.port_b_data_out_clock = "none";
defparam ram_block3a61.port_b_data_width = 1;
defparam ram_block3a61.port_b_first_address = 0;
defparam ram_block3a61.port_b_first_bit_number = 29;
defparam ram_block3a61.port_b_last_address = 8191;
defparam ram_block3a61.port_b_logical_ram_depth = 16384;
defparam ram_block3a61.port_b_logical_ram_width = 32;
defparam ram_block3a61.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block3a61.port_b_read_enable_clock = "clock1";
defparam ram_block3a61.port_b_write_enable_clock = "clock1";
defparam ram_block3a61.ram_block_type = "M9K";
defparam ram_block3a61.mem_init3 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a61.mem_init2 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a61.mem_init1 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a61.mem_init0 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
// synopsys translate_on

// Location: M9K_X78_Y38_N0
cycloneive_ram_block ram_block3a29(
	.portawe(\decode4|eq_node[0]~1_combout ),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(\decode5|eq_node[0]~1_combout ),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock1),
	.ena0(ramaddr),
	.ena1(!ram_rom_addr_reg_13),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({data_a[29]}),
	.portaaddr({address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain({data_b[29]}),
	.portbaddr({address_b[12],address_b[11],address_b[10],address_b[9],address_b[8],address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.devclrn(devclrn),
	.devpor(devpor),
	.portadataout(ram_block3a29_PORTADATAOUT_bus),
	.portbdataout(ram_block3a29_PORTBDATAOUT_bus));
// synopsys translate_off
defparam ram_block3a29.clk0_core_clock_enable = "ena0";
defparam ram_block3a29.clk1_core_clock_enable = "ena1";
defparam ram_block3a29.data_interleave_offset_in_bits = 1;
defparam ram_block3a29.data_interleave_width_in_bits = 1;
defparam ram_block3a29.init_file = "meminit.hex";
defparam ram_block3a29.init_file_layout = "port_a";
defparam ram_block3a29.logical_ram_name = "ram:RAM|altsyncram:altsyncram_component|altsyncram_99f1:auto_generated|altsyncram_fta2:altsyncram1|ALTSYNCRAM";
defparam ram_block3a29.mixed_port_feed_through_mode = "dont_care";
defparam ram_block3a29.operation_mode = "bidir_dual_port";
defparam ram_block3a29.port_a_address_clear = "none";
defparam ram_block3a29.port_a_address_width = 13;
defparam ram_block3a29.port_a_byte_enable_clock = "none";
defparam ram_block3a29.port_a_data_out_clear = "none";
defparam ram_block3a29.port_a_data_out_clock = "none";
defparam ram_block3a29.port_a_data_width = 1;
defparam ram_block3a29.port_a_first_address = 0;
defparam ram_block3a29.port_a_first_bit_number = 29;
defparam ram_block3a29.port_a_last_address = 8191;
defparam ram_block3a29.port_a_logical_ram_depth = 16384;
defparam ram_block3a29.port_a_logical_ram_width = 32;
defparam ram_block3a29.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block3a29.port_b_address_clear = "none";
defparam ram_block3a29.port_b_address_clock = "clock1";
defparam ram_block3a29.port_b_address_width = 13;
defparam ram_block3a29.port_b_data_in_clock = "clock1";
defparam ram_block3a29.port_b_data_out_clear = "none";
defparam ram_block3a29.port_b_data_out_clock = "none";
defparam ram_block3a29.port_b_data_width = 1;
defparam ram_block3a29.port_b_first_address = 0;
defparam ram_block3a29.port_b_first_bit_number = 29;
defparam ram_block3a29.port_b_last_address = 8191;
defparam ram_block3a29.port_b_logical_ram_depth = 16384;
defparam ram_block3a29.port_b_logical_ram_width = 32;
defparam ram_block3a29.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block3a29.port_b_read_enable_clock = "clock1";
defparam ram_block3a29.port_b_write_enable_clock = "clock1";
defparam ram_block3a29.ram_block_type = "M9K";
defparam ram_block3a29.mem_init3 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a29.mem_init2 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a29.mem_init1 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a29.mem_init0 = 2048'h000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000078F3DE001B007700807;
// synopsys translate_on

// Location: M9K_X37_Y30_N0
cycloneive_ram_block ram_block3a62(
	.portawe(\decode4|eq_node[1]~0_combout ),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(\decode5|eq_node[1]~0_combout ),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock1),
	.ena0(!ramaddr),
	.ena1(ram_rom_addr_reg_13),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({data_a[30]}),
	.portaaddr({address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain({data_b[30]}),
	.portbaddr({address_b[12],address_b[11],address_b[10],address_b[9],address_b[8],address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.devclrn(devclrn),
	.devpor(devpor),
	.portadataout(ram_block3a62_PORTADATAOUT_bus),
	.portbdataout(ram_block3a62_PORTBDATAOUT_bus));
// synopsys translate_off
defparam ram_block3a62.clk0_core_clock_enable = "ena0";
defparam ram_block3a62.clk1_core_clock_enable = "ena1";
defparam ram_block3a62.data_interleave_offset_in_bits = 1;
defparam ram_block3a62.data_interleave_width_in_bits = 1;
defparam ram_block3a62.init_file = "meminit.hex";
defparam ram_block3a62.init_file_layout = "port_a";
defparam ram_block3a62.logical_ram_name = "ram:RAM|altsyncram:altsyncram_component|altsyncram_99f1:auto_generated|altsyncram_fta2:altsyncram1|ALTSYNCRAM";
defparam ram_block3a62.mixed_port_feed_through_mode = "dont_care";
defparam ram_block3a62.operation_mode = "bidir_dual_port";
defparam ram_block3a62.port_a_address_clear = "none";
defparam ram_block3a62.port_a_address_width = 13;
defparam ram_block3a62.port_a_byte_enable_clock = "none";
defparam ram_block3a62.port_a_data_out_clear = "none";
defparam ram_block3a62.port_a_data_out_clock = "none";
defparam ram_block3a62.port_a_data_width = 1;
defparam ram_block3a62.port_a_first_address = 0;
defparam ram_block3a62.port_a_first_bit_number = 30;
defparam ram_block3a62.port_a_last_address = 8191;
defparam ram_block3a62.port_a_logical_ram_depth = 16384;
defparam ram_block3a62.port_a_logical_ram_width = 32;
defparam ram_block3a62.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block3a62.port_b_address_clear = "none";
defparam ram_block3a62.port_b_address_clock = "clock1";
defparam ram_block3a62.port_b_address_width = 13;
defparam ram_block3a62.port_b_data_in_clock = "clock1";
defparam ram_block3a62.port_b_data_out_clear = "none";
defparam ram_block3a62.port_b_data_out_clock = "none";
defparam ram_block3a62.port_b_data_width = 1;
defparam ram_block3a62.port_b_first_address = 0;
defparam ram_block3a62.port_b_first_bit_number = 30;
defparam ram_block3a62.port_b_last_address = 8191;
defparam ram_block3a62.port_b_logical_ram_depth = 16384;
defparam ram_block3a62.port_b_logical_ram_width = 32;
defparam ram_block3a62.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block3a62.port_b_read_enable_clock = "clock1";
defparam ram_block3a62.port_b_write_enable_clock = "clock1";
defparam ram_block3a62.ram_block_type = "M9K";
defparam ram_block3a62.mem_init3 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a62.mem_init2 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a62.mem_init1 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a62.mem_init0 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
// synopsys translate_on

// Location: M9K_X64_Y30_N0
cycloneive_ram_block ram_block3a30(
	.portawe(\decode4|eq_node[0]~1_combout ),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(\decode5|eq_node[0]~1_combout ),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock1),
	.ena0(ramaddr),
	.ena1(!ram_rom_addr_reg_13),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({data_a[30]}),
	.portaaddr({address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain({data_b[30]}),
	.portbaddr({address_b[12],address_b[11],address_b[10],address_b[9],address_b[8],address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.devclrn(devclrn),
	.devpor(devpor),
	.portadataout(ram_block3a30_PORTADATAOUT_bus),
	.portbdataout(ram_block3a30_PORTBDATAOUT_bus));
// synopsys translate_off
defparam ram_block3a30.clk0_core_clock_enable = "ena0";
defparam ram_block3a30.clk1_core_clock_enable = "ena1";
defparam ram_block3a30.data_interleave_offset_in_bits = 1;
defparam ram_block3a30.data_interleave_width_in_bits = 1;
defparam ram_block3a30.init_file = "meminit.hex";
defparam ram_block3a30.init_file_layout = "port_a";
defparam ram_block3a30.logical_ram_name = "ram:RAM|altsyncram:altsyncram_component|altsyncram_99f1:auto_generated|altsyncram_fta2:altsyncram1|ALTSYNCRAM";
defparam ram_block3a30.mixed_port_feed_through_mode = "dont_care";
defparam ram_block3a30.operation_mode = "bidir_dual_port";
defparam ram_block3a30.port_a_address_clear = "none";
defparam ram_block3a30.port_a_address_width = 13;
defparam ram_block3a30.port_a_byte_enable_clock = "none";
defparam ram_block3a30.port_a_data_out_clear = "none";
defparam ram_block3a30.port_a_data_out_clock = "none";
defparam ram_block3a30.port_a_data_width = 1;
defparam ram_block3a30.port_a_first_address = 0;
defparam ram_block3a30.port_a_first_bit_number = 30;
defparam ram_block3a30.port_a_last_address = 8191;
defparam ram_block3a30.port_a_logical_ram_depth = 16384;
defparam ram_block3a30.port_a_logical_ram_width = 32;
defparam ram_block3a30.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block3a30.port_b_address_clear = "none";
defparam ram_block3a30.port_b_address_clock = "clock1";
defparam ram_block3a30.port_b_address_width = 13;
defparam ram_block3a30.port_b_data_in_clock = "clock1";
defparam ram_block3a30.port_b_data_out_clear = "none";
defparam ram_block3a30.port_b_data_out_clock = "none";
defparam ram_block3a30.port_b_data_width = 1;
defparam ram_block3a30.port_b_first_address = 0;
defparam ram_block3a30.port_b_first_bit_number = 30;
defparam ram_block3a30.port_b_last_address = 8191;
defparam ram_block3a30.port_b_logical_ram_depth = 16384;
defparam ram_block3a30.port_b_logical_ram_width = 32;
defparam ram_block3a30.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block3a30.port_b_read_enable_clock = "clock1";
defparam ram_block3a30.port_b_write_enable_clock = "clock1";
defparam ram_block3a30.ram_block_type = "M9K";
defparam ram_block3a30.mem_init3 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a30.mem_init2 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a30.mem_init1 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a30.mem_init0 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000002000000;
// synopsys translate_on

// Location: M9K_X51_Y26_N0
cycloneive_ram_block ram_block3a63(
	.portawe(\decode4|eq_node[1]~0_combout ),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(\decode5|eq_node[1]~0_combout ),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock1),
	.ena0(!ramaddr),
	.ena1(ram_rom_addr_reg_13),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({data_a[31]}),
	.portaaddr({address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain({data_b[31]}),
	.portbaddr({address_b[12],address_b[11],address_b[10],address_b[9],address_b[8],address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.devclrn(devclrn),
	.devpor(devpor),
	.portadataout(ram_block3a63_PORTADATAOUT_bus),
	.portbdataout(ram_block3a63_PORTBDATAOUT_bus));
// synopsys translate_off
defparam ram_block3a63.clk0_core_clock_enable = "ena0";
defparam ram_block3a63.clk1_core_clock_enable = "ena1";
defparam ram_block3a63.data_interleave_offset_in_bits = 1;
defparam ram_block3a63.data_interleave_width_in_bits = 1;
defparam ram_block3a63.init_file = "meminit.hex";
defparam ram_block3a63.init_file_layout = "port_a";
defparam ram_block3a63.logical_ram_name = "ram:RAM|altsyncram:altsyncram_component|altsyncram_99f1:auto_generated|altsyncram_fta2:altsyncram1|ALTSYNCRAM";
defparam ram_block3a63.mixed_port_feed_through_mode = "dont_care";
defparam ram_block3a63.operation_mode = "bidir_dual_port";
defparam ram_block3a63.port_a_address_clear = "none";
defparam ram_block3a63.port_a_address_width = 13;
defparam ram_block3a63.port_a_byte_enable_clock = "none";
defparam ram_block3a63.port_a_data_out_clear = "none";
defparam ram_block3a63.port_a_data_out_clock = "none";
defparam ram_block3a63.port_a_data_width = 1;
defparam ram_block3a63.port_a_first_address = 0;
defparam ram_block3a63.port_a_first_bit_number = 31;
defparam ram_block3a63.port_a_last_address = 8191;
defparam ram_block3a63.port_a_logical_ram_depth = 16384;
defparam ram_block3a63.port_a_logical_ram_width = 32;
defparam ram_block3a63.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block3a63.port_b_address_clear = "none";
defparam ram_block3a63.port_b_address_clock = "clock1";
defparam ram_block3a63.port_b_address_width = 13;
defparam ram_block3a63.port_b_data_in_clock = "clock1";
defparam ram_block3a63.port_b_data_out_clear = "none";
defparam ram_block3a63.port_b_data_out_clock = "none";
defparam ram_block3a63.port_b_data_width = 1;
defparam ram_block3a63.port_b_first_address = 0;
defparam ram_block3a63.port_b_first_bit_number = 31;
defparam ram_block3a63.port_b_last_address = 8191;
defparam ram_block3a63.port_b_logical_ram_depth = 16384;
defparam ram_block3a63.port_b_logical_ram_width = 32;
defparam ram_block3a63.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block3a63.port_b_read_enable_clock = "clock1";
defparam ram_block3a63.port_b_write_enable_clock = "clock1";
defparam ram_block3a63.ram_block_type = "M9K";
defparam ram_block3a63.mem_init3 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a63.mem_init2 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a63.mem_init1 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a63.mem_init0 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
// synopsys translate_on

// Location: M9K_X64_Y26_N0
cycloneive_ram_block ram_block3a31(
	.portawe(\decode4|eq_node[0]~1_combout ),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(\decode5|eq_node[0]~1_combout ),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock1),
	.ena0(ramaddr),
	.ena1(!ram_rom_addr_reg_13),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({data_a[31]}),
	.portaaddr({address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain({data_b[31]}),
	.portbaddr({address_b[12],address_b[11],address_b[10],address_b[9],address_b[8],address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.devclrn(devclrn),
	.devpor(devpor),
	.portadataout(ram_block3a31_PORTADATAOUT_bus),
	.portbdataout(ram_block3a31_PORTBDATAOUT_bus));
// synopsys translate_off
defparam ram_block3a31.clk0_core_clock_enable = "ena0";
defparam ram_block3a31.clk1_core_clock_enable = "ena1";
defparam ram_block3a31.data_interleave_offset_in_bits = 1;
defparam ram_block3a31.data_interleave_width_in_bits = 1;
defparam ram_block3a31.init_file = "meminit.hex";
defparam ram_block3a31.init_file_layout = "port_a";
defparam ram_block3a31.logical_ram_name = "ram:RAM|altsyncram:altsyncram_component|altsyncram_99f1:auto_generated|altsyncram_fta2:altsyncram1|ALTSYNCRAM";
defparam ram_block3a31.mixed_port_feed_through_mode = "dont_care";
defparam ram_block3a31.operation_mode = "bidir_dual_port";
defparam ram_block3a31.port_a_address_clear = "none";
defparam ram_block3a31.port_a_address_width = 13;
defparam ram_block3a31.port_a_byte_enable_clock = "none";
defparam ram_block3a31.port_a_data_out_clear = "none";
defparam ram_block3a31.port_a_data_out_clock = "none";
defparam ram_block3a31.port_a_data_width = 1;
defparam ram_block3a31.port_a_first_address = 0;
defparam ram_block3a31.port_a_first_bit_number = 31;
defparam ram_block3a31.port_a_last_address = 8191;
defparam ram_block3a31.port_a_logical_ram_depth = 16384;
defparam ram_block3a31.port_a_logical_ram_width = 32;
defparam ram_block3a31.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block3a31.port_b_address_clear = "none";
defparam ram_block3a31.port_b_address_clock = "clock1";
defparam ram_block3a31.port_b_address_width = 13;
defparam ram_block3a31.port_b_data_in_clock = "clock1";
defparam ram_block3a31.port_b_data_out_clear = "none";
defparam ram_block3a31.port_b_data_out_clock = "none";
defparam ram_block3a31.port_b_data_width = 1;
defparam ram_block3a31.port_b_first_address = 0;
defparam ram_block3a31.port_b_first_bit_number = 31;
defparam ram_block3a31.port_b_last_address = 8191;
defparam ram_block3a31.port_b_logical_ram_depth = 16384;
defparam ram_block3a31.port_b_logical_ram_width = 32;
defparam ram_block3a31.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block3a31.port_b_read_enable_clock = "clock1";
defparam ram_block3a31.port_b_write_enable_clock = "clock1";
defparam ram_block3a31.ram_block_type = "M9K";
defparam ram_block3a31.mem_init3 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a31.mem_init2 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a31.mem_init1 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a31.mem_init0 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000C18426089282400008;
// synopsys translate_on

// Location: FF_X54_Y34_N21
dffeas \address_reg_a[0] (
	.clk(clock0),
	.d(address_a[13]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(address_reg_a_0),
	.prn(vcc));
// synopsys translate_off
defparam \address_reg_a[0] .is_wysiwyg = "true";
defparam \address_reg_a[0] .power_up = "low";
// synopsys translate_on

// Location: FF_X50_Y29_N7
dffeas \address_reg_b[0] (
	.clk(clock1),
	.d(\address_reg_b[0]~feeder_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(address_reg_b_0),
	.prn(vcc));
// synopsys translate_off
defparam \address_reg_b[0] .is_wysiwyg = "true";
defparam \address_reg_b[0] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X50_Y29_N6
cycloneive_lcell_comb \address_reg_b[0]~feeder (
// Equation(s):
// \address_reg_b[0]~feeder_combout  = ram_rom_addr_reg_13

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(ram_rom_addr_reg_13),
	.cin(gnd),
	.combout(\address_reg_b[0]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \address_reg_b[0]~feeder .lut_mask = 16'hFF00;
defparam \address_reg_b[0]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

endmodule

module decode_jsa (
	ramaddr,
	ramWEN,
	always1,
	eq_node_1,
	eq_node_0,
	devpor,
	devclrn,
	devoe);
input 	ramaddr;
input 	ramWEN;
input 	always1;
output 	eq_node_1;
output 	eq_node_0;

// Design Ports Information

input 	devpor;
input 	devclrn;
input 	devoe;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
assign unknown = 1'bx;



// Location: LCCOMB_X54_Y34_N8
cycloneive_lcell_comb \eq_node[1]~0 (
// Equation(s):
// eq_node_1 = (!\ramWEN~0_combout  & (!\ramaddr~27_combout  & always1))

	.dataa(ramWEN),
	.datab(gnd),
	.datac(ramaddr),
	.datad(always1),
	.cin(gnd),
	.combout(eq_node_1),
	.cout());
// synopsys translate_off
defparam \eq_node[1]~0 .lut_mask = 16'h0500;
defparam \eq_node[1]~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y34_N22
cycloneive_lcell_comb \eq_node[0]~1 (
// Equation(s):
// eq_node_0 = (!\ramWEN~0_combout  & (\ramaddr~27_combout  & always1))

	.dataa(ramWEN),
	.datab(gnd),
	.datac(ramaddr),
	.datad(always1),
	.cin(gnd),
	.combout(eq_node_0),
	.cout());
// synopsys translate_off
defparam \eq_node[0]~1 .lut_mask = 16'h5000;
defparam \eq_node[0]~1 .sum_lutc_input = "datac";
// synopsys translate_on

endmodule

module decode_jsa_1 (
	ram_rom_addr_reg_13,
	sdr,
	eq_node_1,
	eq_node_0,
	irf_reg_2_1,
	state_5,
	devpor,
	devclrn,
	devoe);
input 	ram_rom_addr_reg_13;
input 	sdr;
output 	eq_node_1;
output 	eq_node_0;
input 	irf_reg_2_1;
input 	state_5;

// Design Ports Information

input 	devpor;
input 	devclrn;
input 	devoe;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
assign unknown = 1'bx;



// Location: LCCOMB_X46_Y34_N28
cycloneive_lcell_comb \eq_node[1]~0 (
// Equation(s):
// eq_node_1 = (sdr & (\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irf_reg[1][2]~q  & (ram_rom_addr_reg_13 & \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [5])))

	.dataa(sdr),
	.datab(irf_reg_2_1),
	.datac(ram_rom_addr_reg_13),
	.datad(state_5),
	.cin(gnd),
	.combout(eq_node_1),
	.cout());
// synopsys translate_off
defparam \eq_node[1]~0 .lut_mask = 16'h8000;
defparam \eq_node[1]~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X46_Y34_N10
cycloneive_lcell_comb \eq_node[0]~1 (
// Equation(s):
// eq_node_0 = (sdr & (\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irf_reg[1][2]~q  & (!ram_rom_addr_reg_13 & \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [5])))

	.dataa(sdr),
	.datab(irf_reg_2_1),
	.datac(ram_rom_addr_reg_13),
	.datad(state_5),
	.cin(gnd),
	.combout(eq_node_0),
	.cout());
// synopsys translate_off
defparam \eq_node[0]~1 .lut_mask = 16'h0800;
defparam \eq_node[0]~1 .sum_lutc_input = "datac";
// synopsys translate_on

endmodule

module sld_mod_ram_rom (
	ram_block3a32,
	ram_block3a0,
	ram_block3a33,
	ram_block3a1,
	ram_block3a34,
	ram_block3a2,
	ram_block3a35,
	ram_block3a3,
	ram_block3a36,
	ram_block3a4,
	ram_block3a37,
	ram_block3a5,
	ram_block3a38,
	ram_block3a6,
	ram_block3a39,
	ram_block3a7,
	ram_block3a40,
	ram_block3a8,
	ram_block3a41,
	ram_block3a9,
	ram_block3a42,
	ram_block3a10,
	ram_block3a43,
	ram_block3a11,
	ram_block3a44,
	ram_block3a12,
	ram_block3a45,
	ram_block3a13,
	ram_block3a46,
	ram_block3a14,
	ram_block3a47,
	ram_block3a15,
	ram_block3a48,
	ram_block3a16,
	ram_block3a49,
	ram_block3a17,
	ram_block3a50,
	ram_block3a18,
	ram_block3a51,
	ram_block3a19,
	ram_block3a52,
	ram_block3a20,
	ram_block3a53,
	ram_block3a21,
	ram_block3a54,
	ram_block3a22,
	ram_block3a55,
	ram_block3a23,
	ram_block3a56,
	ram_block3a24,
	ram_block3a57,
	ram_block3a25,
	ram_block3a58,
	ram_block3a26,
	ram_block3a59,
	ram_block3a27,
	ram_block3a60,
	ram_block3a28,
	ram_block3a61,
	ram_block3a29,
	ram_block3a62,
	ram_block3a30,
	ram_block3a63,
	ram_block3a31,
	is_in_use_reg1,
	ram_rom_data_reg_0,
	ram_rom_addr_reg_13,
	ram_rom_addr_reg_0,
	ram_rom_addr_reg_1,
	ram_rom_addr_reg_2,
	ram_rom_addr_reg_3,
	ram_rom_addr_reg_4,
	ram_rom_addr_reg_5,
	ram_rom_addr_reg_6,
	ram_rom_addr_reg_7,
	ram_rom_addr_reg_8,
	ram_rom_addr_reg_9,
	ram_rom_addr_reg_10,
	ram_rom_addr_reg_11,
	ram_rom_addr_reg_12,
	ram_rom_data_reg_1,
	ram_rom_data_reg_2,
	ram_rom_data_reg_3,
	ram_rom_data_reg_4,
	ram_rom_data_reg_5,
	ram_rom_data_reg_6,
	ram_rom_data_reg_7,
	ram_rom_data_reg_8,
	ram_rom_data_reg_9,
	ram_rom_data_reg_10,
	ram_rom_data_reg_11,
	ram_rom_data_reg_12,
	ram_rom_data_reg_13,
	ram_rom_data_reg_14,
	ram_rom_data_reg_15,
	ram_rom_data_reg_16,
	ram_rom_data_reg_17,
	ram_rom_data_reg_18,
	ram_rom_data_reg_19,
	ram_rom_data_reg_20,
	ram_rom_data_reg_21,
	ram_rom_data_reg_22,
	ram_rom_data_reg_23,
	ram_rom_data_reg_24,
	ram_rom_data_reg_25,
	ram_rom_data_reg_26,
	ram_rom_data_reg_27,
	ram_rom_data_reg_28,
	ram_rom_data_reg_29,
	ram_rom_data_reg_30,
	ram_rom_data_reg_31,
	ir_loaded_address_reg_0,
	ir_loaded_address_reg_1,
	ir_loaded_address_reg_2,
	ir_loaded_address_reg_3,
	tdo,
	sdr,
	address_reg_b_0,
	altera_internal_jtag,
	state_4,
	ir_in,
	irf_reg_1_1,
	irf_reg_2_1,
	irf_reg_4_1,
	node_ena_1,
	clr,
	virtual_ir_scan_reg,
	state_3,
	state_5,
	state_8,
	raw_tck,
	devpor,
	devclrn,
	devoe);
input 	ram_block3a32;
input 	ram_block3a0;
input 	ram_block3a33;
input 	ram_block3a1;
input 	ram_block3a34;
input 	ram_block3a2;
input 	ram_block3a35;
input 	ram_block3a3;
input 	ram_block3a36;
input 	ram_block3a4;
input 	ram_block3a37;
input 	ram_block3a5;
input 	ram_block3a38;
input 	ram_block3a6;
input 	ram_block3a39;
input 	ram_block3a7;
input 	ram_block3a40;
input 	ram_block3a8;
input 	ram_block3a41;
input 	ram_block3a9;
input 	ram_block3a42;
input 	ram_block3a10;
input 	ram_block3a43;
input 	ram_block3a11;
input 	ram_block3a44;
input 	ram_block3a12;
input 	ram_block3a45;
input 	ram_block3a13;
input 	ram_block3a46;
input 	ram_block3a14;
input 	ram_block3a47;
input 	ram_block3a15;
input 	ram_block3a48;
input 	ram_block3a16;
input 	ram_block3a49;
input 	ram_block3a17;
input 	ram_block3a50;
input 	ram_block3a18;
input 	ram_block3a51;
input 	ram_block3a19;
input 	ram_block3a52;
input 	ram_block3a20;
input 	ram_block3a53;
input 	ram_block3a21;
input 	ram_block3a54;
input 	ram_block3a22;
input 	ram_block3a55;
input 	ram_block3a23;
input 	ram_block3a56;
input 	ram_block3a24;
input 	ram_block3a57;
input 	ram_block3a25;
input 	ram_block3a58;
input 	ram_block3a26;
input 	ram_block3a59;
input 	ram_block3a27;
input 	ram_block3a60;
input 	ram_block3a28;
input 	ram_block3a61;
input 	ram_block3a29;
input 	ram_block3a62;
input 	ram_block3a30;
input 	ram_block3a63;
input 	ram_block3a31;
output 	is_in_use_reg1;
output 	ram_rom_data_reg_0;
output 	ram_rom_addr_reg_13;
output 	ram_rom_addr_reg_0;
output 	ram_rom_addr_reg_1;
output 	ram_rom_addr_reg_2;
output 	ram_rom_addr_reg_3;
output 	ram_rom_addr_reg_4;
output 	ram_rom_addr_reg_5;
output 	ram_rom_addr_reg_6;
output 	ram_rom_addr_reg_7;
output 	ram_rom_addr_reg_8;
output 	ram_rom_addr_reg_9;
output 	ram_rom_addr_reg_10;
output 	ram_rom_addr_reg_11;
output 	ram_rom_addr_reg_12;
output 	ram_rom_data_reg_1;
output 	ram_rom_data_reg_2;
output 	ram_rom_data_reg_3;
output 	ram_rom_data_reg_4;
output 	ram_rom_data_reg_5;
output 	ram_rom_data_reg_6;
output 	ram_rom_data_reg_7;
output 	ram_rom_data_reg_8;
output 	ram_rom_data_reg_9;
output 	ram_rom_data_reg_10;
output 	ram_rom_data_reg_11;
output 	ram_rom_data_reg_12;
output 	ram_rom_data_reg_13;
output 	ram_rom_data_reg_14;
output 	ram_rom_data_reg_15;
output 	ram_rom_data_reg_16;
output 	ram_rom_data_reg_17;
output 	ram_rom_data_reg_18;
output 	ram_rom_data_reg_19;
output 	ram_rom_data_reg_20;
output 	ram_rom_data_reg_21;
output 	ram_rom_data_reg_22;
output 	ram_rom_data_reg_23;
output 	ram_rom_data_reg_24;
output 	ram_rom_data_reg_25;
output 	ram_rom_data_reg_26;
output 	ram_rom_data_reg_27;
output 	ram_rom_data_reg_28;
output 	ram_rom_data_reg_29;
output 	ram_rom_data_reg_30;
output 	ram_rom_data_reg_31;
output 	ir_loaded_address_reg_0;
output 	ir_loaded_address_reg_1;
output 	ir_loaded_address_reg_2;
output 	ir_loaded_address_reg_3;
output 	tdo;
output 	sdr;
input 	address_reg_b_0;
input 	altera_internal_jtag;
input 	state_4;
input 	[4:0] ir_in;
input 	irf_reg_1_1;
input 	irf_reg_2_1;
input 	irf_reg_4_1;
input 	node_ena_1;
input 	clr;
input 	virtual_ir_scan_reg;
input 	state_3;
input 	state_5;
input 	state_8;
input 	raw_tck;

// Design Ports Information

input 	devpor;
input 	devclrn;
input 	devoe;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
assign unknown = 1'bx;

wire \Add1~0_combout ;
wire \Add1~3 ;
wire \Add1~5 ;
wire \Add1~4_combout ;
wire \Add1~7 ;
wire \Add1~6_combout ;
wire \Add1~9 ;
wire \Add1~8_combout ;
wire \Add1~10_combout ;
wire \ram_rom_data_shift_cntr_reg[3]~8_combout ;
wire \is_in_use_reg~0_combout ;
wire \ram_rom_data_reg[0]~0_combout ;
wire \Add1~1 ;
wire \Add1~2_combout ;
wire \ram_rom_data_shift_cntr_reg[5]~4_combout ;
wire \ram_rom_data_shift_cntr_reg[5]~12_combout ;
wire \ram_rom_data_shift_cntr_reg[2]~9_combout ;
wire \ram_rom_data_shift_cntr_reg[5]~10_combout ;
wire \ram_rom_data_shift_cntr_reg[4]~7_combout ;
wire \Equal1~0_combout ;
wire \ram_rom_data_shift_cntr_reg[5]~11_combout ;
wire \ram_rom_data_shift_cntr_reg[0]~6_combout ;
wire \Equal1~1_combout ;
wire \ram_rom_data_shift_cntr_reg[1]~5_combout ;
wire \process_0~2_combout ;
wire \ram_rom_data_reg[12]~32_combout ;
wire \ram_rom_addr_reg[0]~15 ;
wire \ram_rom_addr_reg[1]~17 ;
wire \ram_rom_addr_reg[2]~19 ;
wire \ram_rom_addr_reg[3]~21 ;
wire \ram_rom_addr_reg[4]~23 ;
wire \ram_rom_addr_reg[5]~25 ;
wire \ram_rom_addr_reg[6]~27 ;
wire \ram_rom_addr_reg[7]~29 ;
wire \ram_rom_addr_reg[8]~31 ;
wire \ram_rom_addr_reg[9]~33 ;
wire \ram_rom_addr_reg[10]~35 ;
wire \ram_rom_addr_reg[11]~37 ;
wire \ram_rom_addr_reg[12]~39 ;
wire \ram_rom_addr_reg[13]~40_combout ;
wire \process_0~3_combout ;
wire \ram_rom_addr_reg[5]~42_combout ;
wire \ram_rom_addr_reg[5]~43_combout ;
wire \ram_rom_addr_reg[0]~14_combout ;
wire \ram_rom_addr_reg[1]~16_combout ;
wire \ram_rom_addr_reg[2]~18_combout ;
wire \ram_rom_addr_reg[3]~20_combout ;
wire \ram_rom_addr_reg[4]~22_combout ;
wire \ram_rom_addr_reg[5]~24_combout ;
wire \ram_rom_addr_reg[6]~26_combout ;
wire \ram_rom_addr_reg[7]~28_combout ;
wire \ram_rom_addr_reg[8]~30_combout ;
wire \ram_rom_addr_reg[9]~32_combout ;
wire \ram_rom_addr_reg[10]~34_combout ;
wire \ram_rom_addr_reg[11]~36_combout ;
wire \ram_rom_addr_reg[12]~38_combout ;
wire \ram_rom_data_reg[1]~1_combout ;
wire \ram_rom_data_reg[2]~2_combout ;
wire \ram_rom_data_reg[3]~3_combout ;
wire \ram_rom_data_reg[4]~4_combout ;
wire \ram_rom_data_reg[5]~5_combout ;
wire \ram_rom_data_reg[6]~6_combout ;
wire \ram_rom_data_reg[7]~7_combout ;
wire \ram_rom_data_reg[8]~8_combout ;
wire \ram_rom_data_reg[9]~9_combout ;
wire \ram_rom_data_reg[10]~10_combout ;
wire \ram_rom_data_reg[11]~11_combout ;
wire \ram_rom_data_reg[12]~12_combout ;
wire \ram_rom_data_reg[13]~13_combout ;
wire \ram_rom_data_reg[14]~14_combout ;
wire \ram_rom_data_reg[15]~15_combout ;
wire \ram_rom_data_reg[16]~16_combout ;
wire \ram_rom_data_reg[17]~17_combout ;
wire \ram_rom_data_reg[18]~18_combout ;
wire \ram_rom_data_reg[19]~19_combout ;
wire \ram_rom_data_reg[20]~20_combout ;
wire \ram_rom_data_reg[21]~21_combout ;
wire \ram_rom_data_reg[22]~22_combout ;
wire \ram_rom_data_reg[23]~23_combout ;
wire \ram_rom_data_reg[24]~24_combout ;
wire \ram_rom_data_reg[25]~25_combout ;
wire \ram_rom_data_reg[26]~26_combout ;
wire \ram_rom_data_reg[27]~27_combout ;
wire \ram_rom_data_reg[28]~28_combout ;
wire \ram_rom_data_reg[29]~29_combout ;
wire \ram_rom_data_reg[30]~30_combout ;
wire \ram_rom_data_reg[31]~31_combout ;
wire \ir_loaded_address_reg[0]~feeder_combout ;
wire \process_0~0_combout ;
wire \process_0~1_combout ;
wire \ir_loaded_address_reg[1]~feeder_combout ;
wire \ir_loaded_address_reg[2]~feeder_combout ;
wire \ir_loaded_address_reg[3]~feeder_combout ;
wire \bypass_reg_out~0_combout ;
wire \bypass_reg_out~q ;
wire \tdo~0_combout ;
wire [5:0] ram_rom_data_shift_cntr_reg;
wire [3:0] \ram_rom_logic_gen:name_gen:info_rom_sr|WORD_SR ;


sld_rom_sr \ram_rom_logic_gen:name_gen:info_rom_sr (
	.WORD_SR_0(\ram_rom_logic_gen:name_gen:info_rom_sr|WORD_SR [0]),
	.sdr(sdr),
	.altera_internal_jtag(altera_internal_jtag),
	.state_4(state_4),
	.virtual_ir_scan_reg(virtual_ir_scan_reg),
	.state_3(state_3),
	.state_8(state_8),
	.TCK(raw_tck),
	.devpor(devpor),
	.devclrn(devclrn),
	.devoe(devoe));

// Location: LCCOMB_X47_Y34_N12
cycloneive_lcell_comb \Add1~0 (
	.dataa(ram_rom_data_shift_cntr_reg[0]),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(gnd),
	.combout(\Add1~0_combout ),
	.cout(\Add1~1 ));
// synopsys translate_off
defparam \Add1~0 .lut_mask = 16'h55AA;
defparam \Add1~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X47_Y34_N14
cycloneive_lcell_comb \Add1~2 (
	.dataa(gnd),
	.datab(ram_rom_data_shift_cntr_reg[1]),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add1~1 ),
	.combout(\Add1~2_combout ),
	.cout(\Add1~3 ));
// synopsys translate_off
defparam \Add1~2 .lut_mask = 16'h3C3F;
defparam \Add1~2 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X47_Y34_N16
cycloneive_lcell_comb \Add1~4 (
	.dataa(gnd),
	.datab(ram_rom_data_shift_cntr_reg[2]),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add1~3 ),
	.combout(\Add1~4_combout ),
	.cout(\Add1~5 ));
// synopsys translate_off
defparam \Add1~4 .lut_mask = 16'hC30C;
defparam \Add1~4 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X47_Y34_N18
cycloneive_lcell_comb \Add1~6 (
	.dataa(ram_rom_data_shift_cntr_reg[3]),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add1~5 ),
	.combout(\Add1~6_combout ),
	.cout(\Add1~7 ));
// synopsys translate_off
defparam \Add1~6 .lut_mask = 16'h5A5F;
defparam \Add1~6 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X47_Y34_N20
cycloneive_lcell_comb \Add1~8 (
	.dataa(gnd),
	.datab(ram_rom_data_shift_cntr_reg[4]),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add1~7 ),
	.combout(\Add1~8_combout ),
	.cout(\Add1~9 ));
// synopsys translate_off
defparam \Add1~8 .lut_mask = 16'hC30C;
defparam \Add1~8 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X47_Y34_N22
cycloneive_lcell_comb \Add1~10 (
	.dataa(ram_rom_data_shift_cntr_reg[5]),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.cin(\Add1~9 ),
	.combout(\Add1~10_combout ),
	.cout());
// synopsys translate_off
defparam \Add1~10 .lut_mask = 16'h5A5A;
defparam \Add1~10 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: FF_X47_Y34_N11
dffeas \ram_rom_data_shift_cntr_reg[3] (
	.clk(raw_tck),
	.d(\ram_rom_data_shift_cntr_reg[3]~8_combout ),
	.asdata(vcc),
	.clrn(!ir_in[3]),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(ram_rom_data_shift_cntr_reg[3]),
	.prn(vcc));
// synopsys translate_off
defparam \ram_rom_data_shift_cntr_reg[3] .is_wysiwyg = "true";
defparam \ram_rom_data_shift_cntr_reg[3] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X47_Y34_N10
cycloneive_lcell_comb \ram_rom_data_shift_cntr_reg[3]~8 (
	.dataa(\Add1~6_combout ),
	.datab(\ram_rom_data_shift_cntr_reg[5]~11_combout ),
	.datac(ram_rom_data_shift_cntr_reg[3]),
	.datad(\ram_rom_data_shift_cntr_reg[5]~12_combout ),
	.cin(gnd),
	.combout(\ram_rom_data_shift_cntr_reg[3]~8_combout ),
	.cout());
// synopsys translate_off
defparam \ram_rom_data_shift_cntr_reg[3]~8 .lut_mask = 16'hC0EA;
defparam \ram_rom_data_shift_cntr_reg[3]~8 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X46_Y34_N9
dffeas is_in_use_reg(
	.clk(raw_tck),
	.d(\is_in_use_reg~0_combout ),
	.asdata(vcc),
	.clrn(!clr),
	.aload(gnd),
	.sclr(gnd),
	.sload(ir_in[0]),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(is_in_use_reg1),
	.prn(vcc));
// synopsys translate_off
defparam is_in_use_reg.is_wysiwyg = "true";
defparam is_in_use_reg.power_up = "low";
// synopsys translate_on

// Location: FF_X50_Y29_N17
dffeas \ram_rom_data_reg[0] (
	.clk(raw_tck),
	.d(\ram_rom_data_reg[0]~0_combout ),
	.asdata(ram_rom_data_reg_1),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(\process_0~2_combout ),
	.ena(\ram_rom_data_reg[12]~32_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(ram_rom_data_reg_0),
	.prn(vcc));
// synopsys translate_off
defparam \ram_rom_data_reg[0] .is_wysiwyg = "true";
defparam \ram_rom_data_reg[0] .power_up = "low";
// synopsys translate_on

// Location: FF_X46_Y35_N29
dffeas \ram_rom_addr_reg[13] (
	.clk(raw_tck),
	.d(\ram_rom_addr_reg[13]~40_combout ),
	.asdata(altera_internal_jtag),
	.clrn(!ir_in[0]),
	.aload(gnd),
	.sclr(gnd),
	.sload(\process_0~3_combout ),
	.ena(\ram_rom_addr_reg[5]~43_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(ram_rom_addr_reg_13),
	.prn(vcc));
// synopsys translate_off
defparam \ram_rom_addr_reg[13] .is_wysiwyg = "true";
defparam \ram_rom_addr_reg[13] .power_up = "low";
// synopsys translate_on

// Location: FF_X46_Y35_N3
dffeas \ram_rom_addr_reg[0] (
	.clk(raw_tck),
	.d(\ram_rom_addr_reg[0]~14_combout ),
	.asdata(ram_rom_addr_reg_1),
	.clrn(!ir_in[0]),
	.aload(gnd),
	.sclr(gnd),
	.sload(\process_0~3_combout ),
	.ena(\ram_rom_addr_reg[5]~43_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(ram_rom_addr_reg_0),
	.prn(vcc));
// synopsys translate_off
defparam \ram_rom_addr_reg[0] .is_wysiwyg = "true";
defparam \ram_rom_addr_reg[0] .power_up = "low";
// synopsys translate_on

// Location: FF_X46_Y35_N5
dffeas \ram_rom_addr_reg[1] (
	.clk(raw_tck),
	.d(\ram_rom_addr_reg[1]~16_combout ),
	.asdata(ram_rom_addr_reg_2),
	.clrn(!ir_in[0]),
	.aload(gnd),
	.sclr(gnd),
	.sload(\process_0~3_combout ),
	.ena(\ram_rom_addr_reg[5]~43_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(ram_rom_addr_reg_1),
	.prn(vcc));
// synopsys translate_off
defparam \ram_rom_addr_reg[1] .is_wysiwyg = "true";
defparam \ram_rom_addr_reg[1] .power_up = "low";
// synopsys translate_on

// Location: FF_X46_Y35_N7
dffeas \ram_rom_addr_reg[2] (
	.clk(raw_tck),
	.d(\ram_rom_addr_reg[2]~18_combout ),
	.asdata(ram_rom_addr_reg_3),
	.clrn(!ir_in[0]),
	.aload(gnd),
	.sclr(gnd),
	.sload(\process_0~3_combout ),
	.ena(\ram_rom_addr_reg[5]~43_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(ram_rom_addr_reg_2),
	.prn(vcc));
// synopsys translate_off
defparam \ram_rom_addr_reg[2] .is_wysiwyg = "true";
defparam \ram_rom_addr_reg[2] .power_up = "low";
// synopsys translate_on

// Location: FF_X46_Y35_N9
dffeas \ram_rom_addr_reg[3] (
	.clk(raw_tck),
	.d(\ram_rom_addr_reg[3]~20_combout ),
	.asdata(ram_rom_addr_reg_4),
	.clrn(!ir_in[0]),
	.aload(gnd),
	.sclr(gnd),
	.sload(\process_0~3_combout ),
	.ena(\ram_rom_addr_reg[5]~43_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(ram_rom_addr_reg_3),
	.prn(vcc));
// synopsys translate_off
defparam \ram_rom_addr_reg[3] .is_wysiwyg = "true";
defparam \ram_rom_addr_reg[3] .power_up = "low";
// synopsys translate_on

// Location: FF_X46_Y35_N11
dffeas \ram_rom_addr_reg[4] (
	.clk(raw_tck),
	.d(\ram_rom_addr_reg[4]~22_combout ),
	.asdata(ram_rom_addr_reg_5),
	.clrn(!ir_in[0]),
	.aload(gnd),
	.sclr(gnd),
	.sload(\process_0~3_combout ),
	.ena(\ram_rom_addr_reg[5]~43_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(ram_rom_addr_reg_4),
	.prn(vcc));
// synopsys translate_off
defparam \ram_rom_addr_reg[4] .is_wysiwyg = "true";
defparam \ram_rom_addr_reg[4] .power_up = "low";
// synopsys translate_on

// Location: FF_X46_Y35_N13
dffeas \ram_rom_addr_reg[5] (
	.clk(raw_tck),
	.d(\ram_rom_addr_reg[5]~24_combout ),
	.asdata(ram_rom_addr_reg_6),
	.clrn(!ir_in[0]),
	.aload(gnd),
	.sclr(gnd),
	.sload(\process_0~3_combout ),
	.ena(\ram_rom_addr_reg[5]~43_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(ram_rom_addr_reg_5),
	.prn(vcc));
// synopsys translate_off
defparam \ram_rom_addr_reg[5] .is_wysiwyg = "true";
defparam \ram_rom_addr_reg[5] .power_up = "low";
// synopsys translate_on

// Location: FF_X46_Y35_N15
dffeas \ram_rom_addr_reg[6] (
	.clk(raw_tck),
	.d(\ram_rom_addr_reg[6]~26_combout ),
	.asdata(ram_rom_addr_reg_7),
	.clrn(!ir_in[0]),
	.aload(gnd),
	.sclr(gnd),
	.sload(\process_0~3_combout ),
	.ena(\ram_rom_addr_reg[5]~43_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(ram_rom_addr_reg_6),
	.prn(vcc));
// synopsys translate_off
defparam \ram_rom_addr_reg[6] .is_wysiwyg = "true";
defparam \ram_rom_addr_reg[6] .power_up = "low";
// synopsys translate_on

// Location: FF_X46_Y35_N17
dffeas \ram_rom_addr_reg[7] (
	.clk(raw_tck),
	.d(\ram_rom_addr_reg[7]~28_combout ),
	.asdata(ram_rom_addr_reg_8),
	.clrn(!ir_in[0]),
	.aload(gnd),
	.sclr(gnd),
	.sload(\process_0~3_combout ),
	.ena(\ram_rom_addr_reg[5]~43_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(ram_rom_addr_reg_7),
	.prn(vcc));
// synopsys translate_off
defparam \ram_rom_addr_reg[7] .is_wysiwyg = "true";
defparam \ram_rom_addr_reg[7] .power_up = "low";
// synopsys translate_on

// Location: FF_X46_Y35_N19
dffeas \ram_rom_addr_reg[8] (
	.clk(raw_tck),
	.d(\ram_rom_addr_reg[8]~30_combout ),
	.asdata(ram_rom_addr_reg_9),
	.clrn(!ir_in[0]),
	.aload(gnd),
	.sclr(gnd),
	.sload(\process_0~3_combout ),
	.ena(\ram_rom_addr_reg[5]~43_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(ram_rom_addr_reg_8),
	.prn(vcc));
// synopsys translate_off
defparam \ram_rom_addr_reg[8] .is_wysiwyg = "true";
defparam \ram_rom_addr_reg[8] .power_up = "low";
// synopsys translate_on

// Location: FF_X46_Y35_N21
dffeas \ram_rom_addr_reg[9] (
	.clk(raw_tck),
	.d(\ram_rom_addr_reg[9]~32_combout ),
	.asdata(ram_rom_addr_reg_10),
	.clrn(!ir_in[0]),
	.aload(gnd),
	.sclr(gnd),
	.sload(\process_0~3_combout ),
	.ena(\ram_rom_addr_reg[5]~43_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(ram_rom_addr_reg_9),
	.prn(vcc));
// synopsys translate_off
defparam \ram_rom_addr_reg[9] .is_wysiwyg = "true";
defparam \ram_rom_addr_reg[9] .power_up = "low";
// synopsys translate_on

// Location: FF_X46_Y35_N23
dffeas \ram_rom_addr_reg[10] (
	.clk(raw_tck),
	.d(\ram_rom_addr_reg[10]~34_combout ),
	.asdata(ram_rom_addr_reg_11),
	.clrn(!ir_in[0]),
	.aload(gnd),
	.sclr(gnd),
	.sload(\process_0~3_combout ),
	.ena(\ram_rom_addr_reg[5]~43_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(ram_rom_addr_reg_10),
	.prn(vcc));
// synopsys translate_off
defparam \ram_rom_addr_reg[10] .is_wysiwyg = "true";
defparam \ram_rom_addr_reg[10] .power_up = "low";
// synopsys translate_on

// Location: FF_X46_Y35_N25
dffeas \ram_rom_addr_reg[11] (
	.clk(raw_tck),
	.d(\ram_rom_addr_reg[11]~36_combout ),
	.asdata(ram_rom_addr_reg_12),
	.clrn(!ir_in[0]),
	.aload(gnd),
	.sclr(gnd),
	.sload(\process_0~3_combout ),
	.ena(\ram_rom_addr_reg[5]~43_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(ram_rom_addr_reg_11),
	.prn(vcc));
// synopsys translate_off
defparam \ram_rom_addr_reg[11] .is_wysiwyg = "true";
defparam \ram_rom_addr_reg[11] .power_up = "low";
// synopsys translate_on

// Location: FF_X46_Y35_N27
dffeas \ram_rom_addr_reg[12] (
	.clk(raw_tck),
	.d(\ram_rom_addr_reg[12]~38_combout ),
	.asdata(ram_rom_addr_reg_13),
	.clrn(!ir_in[0]),
	.aload(gnd),
	.sclr(gnd),
	.sload(\process_0~3_combout ),
	.ena(\ram_rom_addr_reg[5]~43_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(ram_rom_addr_reg_12),
	.prn(vcc));
// synopsys translate_off
defparam \ram_rom_addr_reg[12] .is_wysiwyg = "true";
defparam \ram_rom_addr_reg[12] .power_up = "low";
// synopsys translate_on

// Location: FF_X50_Y29_N19
dffeas \ram_rom_data_reg[1] (
	.clk(raw_tck),
	.d(\ram_rom_data_reg[1]~1_combout ),
	.asdata(ram_rom_data_reg_2),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(\process_0~2_combout ),
	.ena(\ram_rom_data_reg[12]~32_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(ram_rom_data_reg_1),
	.prn(vcc));
// synopsys translate_off
defparam \ram_rom_data_reg[1] .is_wysiwyg = "true";
defparam \ram_rom_data_reg[1] .power_up = "low";
// synopsys translate_on

// Location: FF_X50_Y29_N13
dffeas \ram_rom_data_reg[2] (
	.clk(raw_tck),
	.d(\ram_rom_data_reg[2]~2_combout ),
	.asdata(ram_rom_data_reg_3),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(\process_0~2_combout ),
	.ena(\ram_rom_data_reg[12]~32_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(ram_rom_data_reg_2),
	.prn(vcc));
// synopsys translate_off
defparam \ram_rom_data_reg[2] .is_wysiwyg = "true";
defparam \ram_rom_data_reg[2] .power_up = "low";
// synopsys translate_on

// Location: FF_X50_Y29_N31
dffeas \ram_rom_data_reg[3] (
	.clk(raw_tck),
	.d(\ram_rom_data_reg[3]~3_combout ),
	.asdata(ram_rom_data_reg_4),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(\process_0~2_combout ),
	.ena(\ram_rom_data_reg[12]~32_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(ram_rom_data_reg_3),
	.prn(vcc));
// synopsys translate_off
defparam \ram_rom_data_reg[3] .is_wysiwyg = "true";
defparam \ram_rom_data_reg[3] .power_up = "low";
// synopsys translate_on

// Location: FF_X50_Y29_N1
dffeas \ram_rom_data_reg[4] (
	.clk(raw_tck),
	.d(\ram_rom_data_reg[4]~4_combout ),
	.asdata(ram_rom_data_reg_5),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(\process_0~2_combout ),
	.ena(\ram_rom_data_reg[12]~32_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(ram_rom_data_reg_4),
	.prn(vcc));
// synopsys translate_off
defparam \ram_rom_data_reg[4] .is_wysiwyg = "true";
defparam \ram_rom_data_reg[4] .power_up = "low";
// synopsys translate_on

// Location: FF_X50_Y29_N15
dffeas \ram_rom_data_reg[5] (
	.clk(raw_tck),
	.d(\ram_rom_data_reg[5]~5_combout ),
	.asdata(ram_rom_data_reg_6),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(\process_0~2_combout ),
	.ena(\ram_rom_data_reg[12]~32_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(ram_rom_data_reg_5),
	.prn(vcc));
// synopsys translate_off
defparam \ram_rom_data_reg[5] .is_wysiwyg = "true";
defparam \ram_rom_data_reg[5] .power_up = "low";
// synopsys translate_on

// Location: FF_X50_Y29_N9
dffeas \ram_rom_data_reg[6] (
	.clk(raw_tck),
	.d(\ram_rom_data_reg[6]~6_combout ),
	.asdata(ram_rom_data_reg_7),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(\process_0~2_combout ),
	.ena(\ram_rom_data_reg[12]~32_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(ram_rom_data_reg_6),
	.prn(vcc));
// synopsys translate_off
defparam \ram_rom_data_reg[6] .is_wysiwyg = "true";
defparam \ram_rom_data_reg[6] .power_up = "low";
// synopsys translate_on

// Location: FF_X50_Y29_N23
dffeas \ram_rom_data_reg[7] (
	.clk(raw_tck),
	.d(\ram_rom_data_reg[7]~7_combout ),
	.asdata(ram_rom_data_reg_8),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(\process_0~2_combout ),
	.ena(\ram_rom_data_reg[12]~32_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(ram_rom_data_reg_7),
	.prn(vcc));
// synopsys translate_off
defparam \ram_rom_data_reg[7] .is_wysiwyg = "true";
defparam \ram_rom_data_reg[7] .power_up = "low";
// synopsys translate_on

// Location: FF_X50_Y29_N29
dffeas \ram_rom_data_reg[8] (
	.clk(raw_tck),
	.d(\ram_rom_data_reg[8]~8_combout ),
	.asdata(ram_rom_data_reg_9),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(\process_0~2_combout ),
	.ena(\ram_rom_data_reg[12]~32_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(ram_rom_data_reg_8),
	.prn(vcc));
// synopsys translate_off
defparam \ram_rom_data_reg[8] .is_wysiwyg = "true";
defparam \ram_rom_data_reg[8] .power_up = "low";
// synopsys translate_on

// Location: FF_X48_Y35_N13
dffeas \ram_rom_data_reg[9] (
	.clk(raw_tck),
	.d(\ram_rom_data_reg[9]~9_combout ),
	.asdata(ram_rom_data_reg_10),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(\process_0~2_combout ),
	.ena(\ram_rom_data_reg[12]~32_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(ram_rom_data_reg_9),
	.prn(vcc));
// synopsys translate_off
defparam \ram_rom_data_reg[9] .is_wysiwyg = "true";
defparam \ram_rom_data_reg[9] .power_up = "low";
// synopsys translate_on

// Location: FF_X48_Y35_N31
dffeas \ram_rom_data_reg[10] (
	.clk(raw_tck),
	.d(\ram_rom_data_reg[10]~10_combout ),
	.asdata(ram_rom_data_reg_11),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(\process_0~2_combout ),
	.ena(\ram_rom_data_reg[12]~32_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(ram_rom_data_reg_10),
	.prn(vcc));
// synopsys translate_off
defparam \ram_rom_data_reg[10] .is_wysiwyg = "true";
defparam \ram_rom_data_reg[10] .power_up = "low";
// synopsys translate_on

// Location: FF_X48_Y35_N9
dffeas \ram_rom_data_reg[11] (
	.clk(raw_tck),
	.d(\ram_rom_data_reg[11]~11_combout ),
	.asdata(ram_rom_data_reg_12),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(\process_0~2_combout ),
	.ena(\ram_rom_data_reg[12]~32_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(ram_rom_data_reg_11),
	.prn(vcc));
// synopsys translate_off
defparam \ram_rom_data_reg[11] .is_wysiwyg = "true";
defparam \ram_rom_data_reg[11] .power_up = "low";
// synopsys translate_on

// Location: FF_X48_Y35_N27
dffeas \ram_rom_data_reg[12] (
	.clk(raw_tck),
	.d(\ram_rom_data_reg[12]~12_combout ),
	.asdata(ram_rom_data_reg_13),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(\process_0~2_combout ),
	.ena(\ram_rom_data_reg[12]~32_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(ram_rom_data_reg_12),
	.prn(vcc));
// synopsys translate_off
defparam \ram_rom_data_reg[12] .is_wysiwyg = "true";
defparam \ram_rom_data_reg[12] .power_up = "low";
// synopsys translate_on

// Location: FF_X48_Y35_N17
dffeas \ram_rom_data_reg[13] (
	.clk(raw_tck),
	.d(\ram_rom_data_reg[13]~13_combout ),
	.asdata(ram_rom_data_reg_14),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(\process_0~2_combout ),
	.ena(\ram_rom_data_reg[12]~32_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(ram_rom_data_reg_13),
	.prn(vcc));
// synopsys translate_off
defparam \ram_rom_data_reg[13] .is_wysiwyg = "true";
defparam \ram_rom_data_reg[13] .power_up = "low";
// synopsys translate_on

// Location: FF_X48_Y35_N19
dffeas \ram_rom_data_reg[14] (
	.clk(raw_tck),
	.d(\ram_rom_data_reg[14]~14_combout ),
	.asdata(ram_rom_data_reg_15),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(\process_0~2_combout ),
	.ena(\ram_rom_data_reg[12]~32_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(ram_rom_data_reg_14),
	.prn(vcc));
// synopsys translate_off
defparam \ram_rom_data_reg[14] .is_wysiwyg = "true";
defparam \ram_rom_data_reg[14] .power_up = "low";
// synopsys translate_on

// Location: FF_X48_Y35_N29
dffeas \ram_rom_data_reg[15] (
	.clk(raw_tck),
	.d(\ram_rom_data_reg[15]~15_combout ),
	.asdata(ram_rom_data_reg_16),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(\process_0~2_combout ),
	.ena(\ram_rom_data_reg[12]~32_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(ram_rom_data_reg_15),
	.prn(vcc));
// synopsys translate_off
defparam \ram_rom_data_reg[15] .is_wysiwyg = "true";
defparam \ram_rom_data_reg[15] .power_up = "low";
// synopsys translate_on

// Location: FF_X48_Y35_N15
dffeas \ram_rom_data_reg[16] (
	.clk(raw_tck),
	.d(\ram_rom_data_reg[16]~16_combout ),
	.asdata(ram_rom_data_reg_17),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(\process_0~2_combout ),
	.ena(\ram_rom_data_reg[12]~32_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(ram_rom_data_reg_16),
	.prn(vcc));
// synopsys translate_off
defparam \ram_rom_data_reg[16] .is_wysiwyg = "true";
defparam \ram_rom_data_reg[16] .power_up = "low";
// synopsys translate_on

// Location: FF_X48_Y35_N21
dffeas \ram_rom_data_reg[17] (
	.clk(raw_tck),
	.d(\ram_rom_data_reg[17]~17_combout ),
	.asdata(ram_rom_data_reg_18),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(\process_0~2_combout ),
	.ena(\ram_rom_data_reg[12]~32_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(ram_rom_data_reg_17),
	.prn(vcc));
// synopsys translate_off
defparam \ram_rom_data_reg[17] .is_wysiwyg = "true";
defparam \ram_rom_data_reg[17] .power_up = "low";
// synopsys translate_on

// Location: FF_X63_Y29_N25
dffeas \ram_rom_data_reg[18] (
	.clk(raw_tck),
	.d(\ram_rom_data_reg[18]~18_combout ),
	.asdata(ram_rom_data_reg_19),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(\process_0~2_combout ),
	.ena(\ram_rom_data_reg[12]~32_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(ram_rom_data_reg_18),
	.prn(vcc));
// synopsys translate_off
defparam \ram_rom_data_reg[18] .is_wysiwyg = "true";
defparam \ram_rom_data_reg[18] .power_up = "low";
// synopsys translate_on

// Location: FF_X63_Y29_N31
dffeas \ram_rom_data_reg[19] (
	.clk(raw_tck),
	.d(\ram_rom_data_reg[19]~19_combout ),
	.asdata(ram_rom_data_reg_20),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(\process_0~2_combout ),
	.ena(\ram_rom_data_reg[12]~32_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(ram_rom_data_reg_19),
	.prn(vcc));
// synopsys translate_off
defparam \ram_rom_data_reg[19] .is_wysiwyg = "true";
defparam \ram_rom_data_reg[19] .power_up = "low";
// synopsys translate_on

// Location: FF_X74_Y31_N29
dffeas \ram_rom_data_reg[20] (
	.clk(raw_tck),
	.d(\ram_rom_data_reg[20]~20_combout ),
	.asdata(ram_rom_data_reg_21),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(\process_0~2_combout ),
	.ena(\ram_rom_data_reg[12]~32_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(ram_rom_data_reg_20),
	.prn(vcc));
// synopsys translate_off
defparam \ram_rom_data_reg[20] .is_wysiwyg = "true";
defparam \ram_rom_data_reg[20] .power_up = "low";
// synopsys translate_on

// Location: FF_X74_Y31_N27
dffeas \ram_rom_data_reg[21] (
	.clk(raw_tck),
	.d(\ram_rom_data_reg[21]~21_combout ),
	.asdata(ram_rom_data_reg_22),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(\process_0~2_combout ),
	.ena(\ram_rom_data_reg[12]~32_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(ram_rom_data_reg_21),
	.prn(vcc));
// synopsys translate_off
defparam \ram_rom_data_reg[21] .is_wysiwyg = "true";
defparam \ram_rom_data_reg[21] .power_up = "low";
// synopsys translate_on

// Location: FF_X74_Y31_N25
dffeas \ram_rom_data_reg[22] (
	.clk(raw_tck),
	.d(\ram_rom_data_reg[22]~22_combout ),
	.asdata(ram_rom_data_reg_23),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(\process_0~2_combout ),
	.ena(\ram_rom_data_reg[12]~32_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(ram_rom_data_reg_22),
	.prn(vcc));
// synopsys translate_off
defparam \ram_rom_data_reg[22] .is_wysiwyg = "true";
defparam \ram_rom_data_reg[22] .power_up = "low";
// synopsys translate_on

// Location: FF_X74_Y31_N15
dffeas \ram_rom_data_reg[23] (
	.clk(raw_tck),
	.d(\ram_rom_data_reg[23]~23_combout ),
	.asdata(ram_rom_data_reg_24),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(\process_0~2_combout ),
	.ena(\ram_rom_data_reg[12]~32_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(ram_rom_data_reg_23),
	.prn(vcc));
// synopsys translate_off
defparam \ram_rom_data_reg[23] .is_wysiwyg = "true";
defparam \ram_rom_data_reg[23] .power_up = "low";
// synopsys translate_on

// Location: FF_X74_Y31_N1
dffeas \ram_rom_data_reg[24] (
	.clk(raw_tck),
	.d(\ram_rom_data_reg[24]~24_combout ),
	.asdata(ram_rom_data_reg_25),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(\process_0~2_combout ),
	.ena(\ram_rom_data_reg[12]~32_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(ram_rom_data_reg_24),
	.prn(vcc));
// synopsys translate_off
defparam \ram_rom_data_reg[24] .is_wysiwyg = "true";
defparam \ram_rom_data_reg[24] .power_up = "low";
// synopsys translate_on

// Location: FF_X74_Y31_N31
dffeas \ram_rom_data_reg[25] (
	.clk(raw_tck),
	.d(\ram_rom_data_reg[25]~25_combout ),
	.asdata(ram_rom_data_reg_26),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(\process_0~2_combout ),
	.ena(\ram_rom_data_reg[12]~32_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(ram_rom_data_reg_25),
	.prn(vcc));
// synopsys translate_off
defparam \ram_rom_data_reg[25] .is_wysiwyg = "true";
defparam \ram_rom_data_reg[25] .power_up = "low";
// synopsys translate_on

// Location: FF_X74_Y31_N21
dffeas \ram_rom_data_reg[26] (
	.clk(raw_tck),
	.d(\ram_rom_data_reg[26]~26_combout ),
	.asdata(ram_rom_data_reg_27),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(\process_0~2_combout ),
	.ena(\ram_rom_data_reg[12]~32_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(ram_rom_data_reg_26),
	.prn(vcc));
// synopsys translate_off
defparam \ram_rom_data_reg[26] .is_wysiwyg = "true";
defparam \ram_rom_data_reg[26] .power_up = "low";
// synopsys translate_on

// Location: FF_X74_Y31_N11
dffeas \ram_rom_data_reg[27] (
	.clk(raw_tck),
	.d(\ram_rom_data_reg[27]~27_combout ),
	.asdata(ram_rom_data_reg_28),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(\process_0~2_combout ),
	.ena(\ram_rom_data_reg[12]~32_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(ram_rom_data_reg_27),
	.prn(vcc));
// synopsys translate_off
defparam \ram_rom_data_reg[27] .is_wysiwyg = "true";
defparam \ram_rom_data_reg[27] .power_up = "low";
// synopsys translate_on

// Location: FF_X74_Y31_N9
dffeas \ram_rom_data_reg[28] (
	.clk(raw_tck),
	.d(\ram_rom_data_reg[28]~28_combout ),
	.asdata(ram_rom_data_reg_29),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(\process_0~2_combout ),
	.ena(\ram_rom_data_reg[12]~32_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(ram_rom_data_reg_28),
	.prn(vcc));
// synopsys translate_off
defparam \ram_rom_data_reg[28] .is_wysiwyg = "true";
defparam \ram_rom_data_reg[28] .power_up = "low";
// synopsys translate_on

// Location: FF_X74_Y31_N19
dffeas \ram_rom_data_reg[29] (
	.clk(raw_tck),
	.d(\ram_rom_data_reg[29]~29_combout ),
	.asdata(ram_rom_data_reg_30),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(\process_0~2_combout ),
	.ena(\ram_rom_data_reg[12]~32_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(ram_rom_data_reg_29),
	.prn(vcc));
// synopsys translate_off
defparam \ram_rom_data_reg[29] .is_wysiwyg = "true";
defparam \ram_rom_data_reg[29] .power_up = "low";
// synopsys translate_on

// Location: FF_X50_Y29_N27
dffeas \ram_rom_data_reg[30] (
	.clk(raw_tck),
	.d(\ram_rom_data_reg[30]~30_combout ),
	.asdata(ram_rom_data_reg_31),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(\process_0~2_combout ),
	.ena(\ram_rom_data_reg[12]~32_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(ram_rom_data_reg_30),
	.prn(vcc));
// synopsys translate_off
defparam \ram_rom_data_reg[30] .is_wysiwyg = "true";
defparam \ram_rom_data_reg[30] .power_up = "low";
// synopsys translate_on

// Location: FF_X50_Y29_N25
dffeas \ram_rom_data_reg[31] (
	.clk(raw_tck),
	.d(\ram_rom_data_reg[31]~31_combout ),
	.asdata(altera_internal_jtag),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(\process_0~2_combout ),
	.ena(\ram_rom_data_reg[12]~32_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(ram_rom_data_reg_31),
	.prn(vcc));
// synopsys translate_off
defparam \ram_rom_data_reg[31] .is_wysiwyg = "true";
defparam \ram_rom_data_reg[31] .power_up = "low";
// synopsys translate_on

// Location: FF_X46_Y34_N31
dffeas \ir_loaded_address_reg[0] (
	.clk(raw_tck),
	.d(\ir_loaded_address_reg[0]~feeder_combout ),
	.asdata(vcc),
	.clrn(!\process_0~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\process_0~1_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(ir_loaded_address_reg_0),
	.prn(vcc));
// synopsys translate_off
defparam \ir_loaded_address_reg[0] .is_wysiwyg = "true";
defparam \ir_loaded_address_reg[0] .power_up = "low";
// synopsys translate_on

// Location: FF_X46_Y31_N1
dffeas \ir_loaded_address_reg[1] (
	.clk(raw_tck),
	.d(\ir_loaded_address_reg[1]~feeder_combout ),
	.asdata(vcc),
	.clrn(!\process_0~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\process_0~1_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(ir_loaded_address_reg_1),
	.prn(vcc));
// synopsys translate_off
defparam \ir_loaded_address_reg[1] .is_wysiwyg = "true";
defparam \ir_loaded_address_reg[1] .power_up = "low";
// synopsys translate_on

// Location: FF_X46_Y31_N11
dffeas \ir_loaded_address_reg[2] (
	.clk(raw_tck),
	.d(\ir_loaded_address_reg[2]~feeder_combout ),
	.asdata(vcc),
	.clrn(!\process_0~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\process_0~1_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(ir_loaded_address_reg_2),
	.prn(vcc));
// synopsys translate_off
defparam \ir_loaded_address_reg[2] .is_wysiwyg = "true";
defparam \ir_loaded_address_reg[2] .power_up = "low";
// synopsys translate_on

// Location: FF_X46_Y31_N5
dffeas \ir_loaded_address_reg[3] (
	.clk(raw_tck),
	.d(\ir_loaded_address_reg[3]~feeder_combout ),
	.asdata(vcc),
	.clrn(!\process_0~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\process_0~1_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(ir_loaded_address_reg_3),
	.prn(vcc));
// synopsys translate_off
defparam \ir_loaded_address_reg[3] .is_wysiwyg = "true";
defparam \ir_loaded_address_reg[3] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X46_Y34_N20
cycloneive_lcell_comb \tdo~1 (
	.dataa(\ram_rom_logic_gen:name_gen:info_rom_sr|WORD_SR [0]),
	.datab(gnd),
	.datac(ir_in[0]),
	.datad(\tdo~0_combout ),
	.cin(gnd),
	.combout(tdo),
	.cout());
// synopsys translate_off
defparam \tdo~1 .lut_mask = 16'hAFA0;
defparam \tdo~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X46_Y34_N6
cycloneive_lcell_comb \sdr~0 (
	.dataa(gnd),
	.datab(gnd),
	.datac(virtual_ir_scan_reg),
	.datad(node_ena_1),
	.cin(gnd),
	.combout(sdr),
	.cout());
// synopsys translate_off
defparam \sdr~0 .lut_mask = 16'h0F00;
defparam \sdr~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X46_Y34_N8
cycloneive_lcell_comb \is_in_use_reg~0 (
	.dataa(gnd),
	.datab(gnd),
	.datac(is_in_use_reg1),
	.datad(irf_reg_4_1),
	.cin(gnd),
	.combout(\is_in_use_reg~0_combout ),
	.cout());
// synopsys translate_off
defparam \is_in_use_reg~0 .lut_mask = 16'h00F0;
defparam \is_in_use_reg~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X50_Y29_N16
cycloneive_lcell_comb \ram_rom_data_reg[0]~0 (
	.dataa(address_reg_b_0),
	.datab(ram_block3a0),
	.datac(gnd),
	.datad(ram_block3a32),
	.cin(gnd),
	.combout(\ram_rom_data_reg[0]~0_combout ),
	.cout());
// synopsys translate_off
defparam \ram_rom_data_reg[0]~0 .lut_mask = 16'hEE44;
defparam \ram_rom_data_reg[0]~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X46_Y34_N26
cycloneive_lcell_comb \ram_rom_data_shift_cntr_reg[5]~4 (
	.dataa(sdr),
	.datab(state_4),
	.datac(irf_reg_1_1),
	.datad(irf_reg_2_1),
	.cin(gnd),
	.combout(\ram_rom_data_shift_cntr_reg[5]~4_combout ),
	.cout());
// synopsys translate_off
defparam \ram_rom_data_shift_cntr_reg[5]~4 .lut_mask = 16'h8880;
defparam \ram_rom_data_shift_cntr_reg[5]~4 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X47_Y34_N2
cycloneive_lcell_comb \ram_rom_data_shift_cntr_reg[5]~12 (
	.dataa(ram_rom_data_shift_cntr_reg[0]),
	.datab(ram_rom_data_shift_cntr_reg[1]),
	.datac(\ram_rom_data_shift_cntr_reg[5]~4_combout ),
	.datad(\Equal1~0_combout ),
	.cin(gnd),
	.combout(\ram_rom_data_shift_cntr_reg[5]~12_combout ),
	.cout());
// synopsys translate_off
defparam \ram_rom_data_shift_cntr_reg[5]~12 .lut_mask = 16'h8F0F;
defparam \ram_rom_data_shift_cntr_reg[5]~12 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X47_Y34_N8
cycloneive_lcell_comb \ram_rom_data_shift_cntr_reg[2]~9 (
	.dataa(\Add1~4_combout ),
	.datab(\ram_rom_data_shift_cntr_reg[5]~11_combout ),
	.datac(ram_rom_data_shift_cntr_reg[2]),
	.datad(\ram_rom_data_shift_cntr_reg[5]~12_combout ),
	.cin(gnd),
	.combout(\ram_rom_data_shift_cntr_reg[2]~9_combout ),
	.cout());
// synopsys translate_off
defparam \ram_rom_data_shift_cntr_reg[2]~9 .lut_mask = 16'hC0EA;
defparam \ram_rom_data_shift_cntr_reg[2]~9 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X47_Y34_N9
dffeas \ram_rom_data_shift_cntr_reg[2] (
	.clk(raw_tck),
	.d(\ram_rom_data_shift_cntr_reg[2]~9_combout ),
	.asdata(vcc),
	.clrn(!ir_in[3]),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(ram_rom_data_shift_cntr_reg[2]),
	.prn(vcc));
// synopsys translate_off
defparam \ram_rom_data_shift_cntr_reg[2] .is_wysiwyg = "true";
defparam \ram_rom_data_shift_cntr_reg[2] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X47_Y34_N26
cycloneive_lcell_comb \ram_rom_data_shift_cntr_reg[5]~10 (
	.dataa(\Add1~10_combout ),
	.datab(\ram_rom_data_shift_cntr_reg[5]~11_combout ),
	.datac(ram_rom_data_shift_cntr_reg[5]),
	.datad(\ram_rom_data_shift_cntr_reg[5]~12_combout ),
	.cin(gnd),
	.combout(\ram_rom_data_shift_cntr_reg[5]~10_combout ),
	.cout());
// synopsys translate_off
defparam \ram_rom_data_shift_cntr_reg[5]~10 .lut_mask = 16'hC0EA;
defparam \ram_rom_data_shift_cntr_reg[5]~10 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X47_Y34_N27
dffeas \ram_rom_data_shift_cntr_reg[5] (
	.clk(raw_tck),
	.d(\ram_rom_data_shift_cntr_reg[5]~10_combout ),
	.asdata(vcc),
	.clrn(!ir_in[3]),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(ram_rom_data_shift_cntr_reg[5]),
	.prn(vcc));
// synopsys translate_off
defparam \ram_rom_data_shift_cntr_reg[5] .is_wysiwyg = "true";
defparam \ram_rom_data_shift_cntr_reg[5] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X47_Y34_N24
cycloneive_lcell_comb \ram_rom_data_shift_cntr_reg[4]~7 (
	.dataa(\Add1~8_combout ),
	.datab(\ram_rom_data_shift_cntr_reg[5]~11_combout ),
	.datac(ram_rom_data_shift_cntr_reg[4]),
	.datad(\ram_rom_data_shift_cntr_reg[5]~12_combout ),
	.cin(gnd),
	.combout(\ram_rom_data_shift_cntr_reg[4]~7_combout ),
	.cout());
// synopsys translate_off
defparam \ram_rom_data_shift_cntr_reg[4]~7 .lut_mask = 16'hC0EA;
defparam \ram_rom_data_shift_cntr_reg[4]~7 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X47_Y34_N25
dffeas \ram_rom_data_shift_cntr_reg[4] (
	.clk(raw_tck),
	.d(\ram_rom_data_shift_cntr_reg[4]~7_combout ),
	.asdata(vcc),
	.clrn(!ir_in[3]),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(ram_rom_data_shift_cntr_reg[4]),
	.prn(vcc));
// synopsys translate_off
defparam \ram_rom_data_shift_cntr_reg[4] .is_wysiwyg = "true";
defparam \ram_rom_data_shift_cntr_reg[4] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X47_Y34_N0
cycloneive_lcell_comb \Equal1~0 (
	.dataa(ram_rom_data_shift_cntr_reg[3]),
	.datab(ram_rom_data_shift_cntr_reg[2]),
	.datac(ram_rom_data_shift_cntr_reg[5]),
	.datad(ram_rom_data_shift_cntr_reg[4]),
	.cin(gnd),
	.combout(\Equal1~0_combout ),
	.cout());
// synopsys translate_off
defparam \Equal1~0 .lut_mask = 16'h0800;
defparam \Equal1~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X47_Y34_N28
cycloneive_lcell_comb \ram_rom_data_shift_cntr_reg[5]~11 (
	.dataa(ram_rom_data_shift_cntr_reg[0]),
	.datab(ram_rom_data_shift_cntr_reg[1]),
	.datac(\ram_rom_data_shift_cntr_reg[5]~4_combout ),
	.datad(\Equal1~0_combout ),
	.cin(gnd),
	.combout(\ram_rom_data_shift_cntr_reg[5]~11_combout ),
	.cout());
// synopsys translate_off
defparam \ram_rom_data_shift_cntr_reg[5]~11 .lut_mask = 16'h070F;
defparam \ram_rom_data_shift_cntr_reg[5]~11 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X47_Y34_N30
cycloneive_lcell_comb \ram_rom_data_shift_cntr_reg[0]~6 (
	.dataa(\Add1~0_combout ),
	.datab(\ram_rom_data_shift_cntr_reg[5]~11_combout ),
	.datac(ram_rom_data_shift_cntr_reg[0]),
	.datad(\ram_rom_data_shift_cntr_reg[5]~12_combout ),
	.cin(gnd),
	.combout(\ram_rom_data_shift_cntr_reg[0]~6_combout ),
	.cout());
// synopsys translate_off
defparam \ram_rom_data_shift_cntr_reg[0]~6 .lut_mask = 16'hC0EA;
defparam \ram_rom_data_shift_cntr_reg[0]~6 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X47_Y34_N31
dffeas \ram_rom_data_shift_cntr_reg[0] (
	.clk(raw_tck),
	.d(\ram_rom_data_shift_cntr_reg[0]~6_combout ),
	.asdata(vcc),
	.clrn(!ir_in[3]),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(ram_rom_data_shift_cntr_reg[0]),
	.prn(vcc));
// synopsys translate_off
defparam \ram_rom_data_shift_cntr_reg[0] .is_wysiwyg = "true";
defparam \ram_rom_data_shift_cntr_reg[0] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X47_Y34_N6
cycloneive_lcell_comb \Equal1~1 (
	.dataa(gnd),
	.datab(gnd),
	.datac(ram_rom_data_shift_cntr_reg[0]),
	.datad(\Equal1~0_combout ),
	.cin(gnd),
	.combout(\Equal1~1_combout ),
	.cout());
// synopsys translate_off
defparam \Equal1~1 .lut_mask = 16'hF000;
defparam \Equal1~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X47_Y34_N4
cycloneive_lcell_comb \ram_rom_data_shift_cntr_reg[1]~5 (
	.dataa(\ram_rom_data_shift_cntr_reg[5]~4_combout ),
	.datab(\Add1~2_combout ),
	.datac(ram_rom_data_shift_cntr_reg[1]),
	.datad(\Equal1~1_combout ),
	.cin(gnd),
	.combout(\ram_rom_data_shift_cntr_reg[1]~5_combout ),
	.cout());
// synopsys translate_off
defparam \ram_rom_data_shift_cntr_reg[1]~5 .lut_mask = 16'h08D8;
defparam \ram_rom_data_shift_cntr_reg[1]~5 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X47_Y34_N5
dffeas \ram_rom_data_shift_cntr_reg[1] (
	.clk(raw_tck),
	.d(\ram_rom_data_shift_cntr_reg[1]~5_combout ),
	.asdata(vcc),
	.clrn(!ir_in[3]),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(ram_rom_data_shift_cntr_reg[1]),
	.prn(vcc));
// synopsys translate_off
defparam \ram_rom_data_shift_cntr_reg[1] .is_wysiwyg = "true";
defparam \ram_rom_data_shift_cntr_reg[1] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X46_Y34_N12
cycloneive_lcell_comb \process_0~2 (
	.dataa(ram_rom_data_shift_cntr_reg[1]),
	.datab(irf_reg_1_1),
	.datac(ir_in[3]),
	.datad(\Equal1~1_combout ),
	.cin(gnd),
	.combout(\process_0~2_combout ),
	.cout());
// synopsys translate_off
defparam \process_0~2 .lut_mask = 16'h070F;
defparam \process_0~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X48_Y35_N6
cycloneive_lcell_comb \ram_rom_data_reg[12]~32 (
	.dataa(\process_0~2_combout ),
	.datab(gnd),
	.datac(\ram_rom_data_shift_cntr_reg[5]~4_combout ),
	.datad(gnd),
	.cin(gnd),
	.combout(\ram_rom_data_reg[12]~32_combout ),
	.cout());
// synopsys translate_off
defparam \ram_rom_data_reg[12]~32 .lut_mask = 16'hF5F5;
defparam \ram_rom_data_reg[12]~32 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X46_Y35_N2
cycloneive_lcell_comb \ram_rom_addr_reg[0]~14 (
	.dataa(gnd),
	.datab(ram_rom_addr_reg_0),
	.datac(gnd),
	.datad(vcc),
	.cin(gnd),
	.combout(\ram_rom_addr_reg[0]~14_combout ),
	.cout(\ram_rom_addr_reg[0]~15 ));
// synopsys translate_off
defparam \ram_rom_addr_reg[0]~14 .lut_mask = 16'h33CC;
defparam \ram_rom_addr_reg[0]~14 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X46_Y35_N4
cycloneive_lcell_comb \ram_rom_addr_reg[1]~16 (
	.dataa(gnd),
	.datab(ram_rom_addr_reg_1),
	.datac(gnd),
	.datad(vcc),
	.cin(\ram_rom_addr_reg[0]~15 ),
	.combout(\ram_rom_addr_reg[1]~16_combout ),
	.cout(\ram_rom_addr_reg[1]~17 ));
// synopsys translate_off
defparam \ram_rom_addr_reg[1]~16 .lut_mask = 16'h3C3F;
defparam \ram_rom_addr_reg[1]~16 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X46_Y35_N6
cycloneive_lcell_comb \ram_rom_addr_reg[2]~18 (
	.dataa(gnd),
	.datab(ram_rom_addr_reg_2),
	.datac(gnd),
	.datad(vcc),
	.cin(\ram_rom_addr_reg[1]~17 ),
	.combout(\ram_rom_addr_reg[2]~18_combout ),
	.cout(\ram_rom_addr_reg[2]~19 ));
// synopsys translate_off
defparam \ram_rom_addr_reg[2]~18 .lut_mask = 16'hC30C;
defparam \ram_rom_addr_reg[2]~18 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X46_Y35_N8
cycloneive_lcell_comb \ram_rom_addr_reg[3]~20 (
	.dataa(gnd),
	.datab(ram_rom_addr_reg_3),
	.datac(gnd),
	.datad(vcc),
	.cin(\ram_rom_addr_reg[2]~19 ),
	.combout(\ram_rom_addr_reg[3]~20_combout ),
	.cout(\ram_rom_addr_reg[3]~21 ));
// synopsys translate_off
defparam \ram_rom_addr_reg[3]~20 .lut_mask = 16'h3C3F;
defparam \ram_rom_addr_reg[3]~20 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X46_Y35_N10
cycloneive_lcell_comb \ram_rom_addr_reg[4]~22 (
	.dataa(gnd),
	.datab(ram_rom_addr_reg_4),
	.datac(gnd),
	.datad(vcc),
	.cin(\ram_rom_addr_reg[3]~21 ),
	.combout(\ram_rom_addr_reg[4]~22_combout ),
	.cout(\ram_rom_addr_reg[4]~23 ));
// synopsys translate_off
defparam \ram_rom_addr_reg[4]~22 .lut_mask = 16'hC30C;
defparam \ram_rom_addr_reg[4]~22 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X46_Y35_N12
cycloneive_lcell_comb \ram_rom_addr_reg[5]~24 (
	.dataa(gnd),
	.datab(ram_rom_addr_reg_5),
	.datac(gnd),
	.datad(vcc),
	.cin(\ram_rom_addr_reg[4]~23 ),
	.combout(\ram_rom_addr_reg[5]~24_combout ),
	.cout(\ram_rom_addr_reg[5]~25 ));
// synopsys translate_off
defparam \ram_rom_addr_reg[5]~24 .lut_mask = 16'h3C3F;
defparam \ram_rom_addr_reg[5]~24 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X46_Y35_N14
cycloneive_lcell_comb \ram_rom_addr_reg[6]~26 (
	.dataa(gnd),
	.datab(ram_rom_addr_reg_6),
	.datac(gnd),
	.datad(vcc),
	.cin(\ram_rom_addr_reg[5]~25 ),
	.combout(\ram_rom_addr_reg[6]~26_combout ),
	.cout(\ram_rom_addr_reg[6]~27 ));
// synopsys translate_off
defparam \ram_rom_addr_reg[6]~26 .lut_mask = 16'hC30C;
defparam \ram_rom_addr_reg[6]~26 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X46_Y35_N16
cycloneive_lcell_comb \ram_rom_addr_reg[7]~28 (
	.dataa(ram_rom_addr_reg_7),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\ram_rom_addr_reg[6]~27 ),
	.combout(\ram_rom_addr_reg[7]~28_combout ),
	.cout(\ram_rom_addr_reg[7]~29 ));
// synopsys translate_off
defparam \ram_rom_addr_reg[7]~28 .lut_mask = 16'h5A5F;
defparam \ram_rom_addr_reg[7]~28 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X46_Y35_N18
cycloneive_lcell_comb \ram_rom_addr_reg[8]~30 (
	.dataa(ram_rom_addr_reg_8),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\ram_rom_addr_reg[7]~29 ),
	.combout(\ram_rom_addr_reg[8]~30_combout ),
	.cout(\ram_rom_addr_reg[8]~31 ));
// synopsys translate_off
defparam \ram_rom_addr_reg[8]~30 .lut_mask = 16'hA50A;
defparam \ram_rom_addr_reg[8]~30 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X46_Y35_N20
cycloneive_lcell_comb \ram_rom_addr_reg[9]~32 (
	.dataa(ram_rom_addr_reg_9),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\ram_rom_addr_reg[8]~31 ),
	.combout(\ram_rom_addr_reg[9]~32_combout ),
	.cout(\ram_rom_addr_reg[9]~33 ));
// synopsys translate_off
defparam \ram_rom_addr_reg[9]~32 .lut_mask = 16'h5A5F;
defparam \ram_rom_addr_reg[9]~32 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X46_Y35_N22
cycloneive_lcell_comb \ram_rom_addr_reg[10]~34 (
	.dataa(ram_rom_addr_reg_10),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\ram_rom_addr_reg[9]~33 ),
	.combout(\ram_rom_addr_reg[10]~34_combout ),
	.cout(\ram_rom_addr_reg[10]~35 ));
// synopsys translate_off
defparam \ram_rom_addr_reg[10]~34 .lut_mask = 16'hA50A;
defparam \ram_rom_addr_reg[10]~34 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X46_Y35_N24
cycloneive_lcell_comb \ram_rom_addr_reg[11]~36 (
	.dataa(ram_rom_addr_reg_11),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\ram_rom_addr_reg[10]~35 ),
	.combout(\ram_rom_addr_reg[11]~36_combout ),
	.cout(\ram_rom_addr_reg[11]~37 ));
// synopsys translate_off
defparam \ram_rom_addr_reg[11]~36 .lut_mask = 16'h5A5F;
defparam \ram_rom_addr_reg[11]~36 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X46_Y35_N26
cycloneive_lcell_comb \ram_rom_addr_reg[12]~38 (
	.dataa(ram_rom_addr_reg_12),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\ram_rom_addr_reg[11]~37 ),
	.combout(\ram_rom_addr_reg[12]~38_combout ),
	.cout(\ram_rom_addr_reg[12]~39 ));
// synopsys translate_off
defparam \ram_rom_addr_reg[12]~38 .lut_mask = 16'hA50A;
defparam \ram_rom_addr_reg[12]~38 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X46_Y35_N28
cycloneive_lcell_comb \ram_rom_addr_reg[13]~40 (
	.dataa(gnd),
	.datab(ram_rom_addr_reg_13),
	.datac(gnd),
	.datad(gnd),
	.cin(\ram_rom_addr_reg[12]~39 ),
	.combout(\ram_rom_addr_reg[13]~40_combout ),
	.cout());
// synopsys translate_off
defparam \ram_rom_addr_reg[13]~40 .lut_mask = 16'h3C3C;
defparam \ram_rom_addr_reg[13]~40 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X46_Y34_N0
cycloneive_lcell_comb \process_0~3 (
	.dataa(node_ena_1),
	.datab(ir_in[3]),
	.datac(virtual_ir_scan_reg),
	.datad(state_4),
	.cin(gnd),
	.combout(\process_0~3_combout ),
	.cout());
// synopsys translate_off
defparam \process_0~3 .lut_mask = 16'h0800;
defparam \process_0~3 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X46_Y34_N22
cycloneive_lcell_comb \ram_rom_addr_reg[5]~42 (
	.dataa(ram_rom_data_shift_cntr_reg[1]),
	.datab(\process_0~3_combout ),
	.datac(irf_reg_1_1),
	.datad(\Equal1~1_combout ),
	.cin(gnd),
	.combout(\ram_rom_addr_reg[5]~42_combout ),
	.cout());
// synopsys translate_off
defparam \ram_rom_addr_reg[5]~42 .lut_mask = 16'hDCCC;
defparam \ram_rom_addr_reg[5]~42 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X46_Y34_N4
cycloneive_lcell_comb \ram_rom_addr_reg[5]~43 (
	.dataa(sdr),
	.datab(state_8),
	.datac(\ram_rom_addr_reg[5]~42_combout ),
	.datad(irf_reg_2_1),
	.cin(gnd),
	.combout(\ram_rom_addr_reg[5]~43_combout ),
	.cout());
// synopsys translate_off
defparam \ram_rom_addr_reg[5]~43 .lut_mask = 16'hF8F0;
defparam \ram_rom_addr_reg[5]~43 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X50_Y29_N18
cycloneive_lcell_comb \ram_rom_data_reg[1]~1 (
	.dataa(address_reg_b_0),
	.datab(ram_block3a33),
	.datac(gnd),
	.datad(ram_block3a1),
	.cin(gnd),
	.combout(\ram_rom_data_reg[1]~1_combout ),
	.cout());
// synopsys translate_off
defparam \ram_rom_data_reg[1]~1 .lut_mask = 16'hDD88;
defparam \ram_rom_data_reg[1]~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X50_Y29_N12
cycloneive_lcell_comb \ram_rom_data_reg[2]~2 (
	.dataa(address_reg_b_0),
	.datab(ram_block3a2),
	.datac(gnd),
	.datad(ram_block3a34),
	.cin(gnd),
	.combout(\ram_rom_data_reg[2]~2_combout ),
	.cout());
// synopsys translate_off
defparam \ram_rom_data_reg[2]~2 .lut_mask = 16'hEE44;
defparam \ram_rom_data_reg[2]~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X50_Y29_N30
cycloneive_lcell_comb \ram_rom_data_reg[3]~3 (
	.dataa(address_reg_b_0),
	.datab(ram_block3a3),
	.datac(gnd),
	.datad(ram_block3a35),
	.cin(gnd),
	.combout(\ram_rom_data_reg[3]~3_combout ),
	.cout());
// synopsys translate_off
defparam \ram_rom_data_reg[3]~3 .lut_mask = 16'hEE44;
defparam \ram_rom_data_reg[3]~3 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X50_Y29_N0
cycloneive_lcell_comb \ram_rom_data_reg[4]~4 (
	.dataa(ram_block3a4),
	.datab(ram_block3a36),
	.datac(gnd),
	.datad(address_reg_b_0),
	.cin(gnd),
	.combout(\ram_rom_data_reg[4]~4_combout ),
	.cout());
// synopsys translate_off
defparam \ram_rom_data_reg[4]~4 .lut_mask = 16'hCCAA;
defparam \ram_rom_data_reg[4]~4 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X50_Y29_N14
cycloneive_lcell_comb \ram_rom_data_reg[5]~5 (
	.dataa(address_reg_b_0),
	.datab(ram_block3a37),
	.datac(gnd),
	.datad(ram_block3a5),
	.cin(gnd),
	.combout(\ram_rom_data_reg[5]~5_combout ),
	.cout());
// synopsys translate_off
defparam \ram_rom_data_reg[5]~5 .lut_mask = 16'hDD88;
defparam \ram_rom_data_reg[5]~5 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X50_Y29_N8
cycloneive_lcell_comb \ram_rom_data_reg[6]~6 (
	.dataa(address_reg_b_0),
	.datab(ram_block3a38),
	.datac(gnd),
	.datad(ram_block3a6),
	.cin(gnd),
	.combout(\ram_rom_data_reg[6]~6_combout ),
	.cout());
// synopsys translate_off
defparam \ram_rom_data_reg[6]~6 .lut_mask = 16'hDD88;
defparam \ram_rom_data_reg[6]~6 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X50_Y29_N22
cycloneive_lcell_comb \ram_rom_data_reg[7]~7 (
	.dataa(address_reg_b_0),
	.datab(ram_block3a39),
	.datac(gnd),
	.datad(ram_block3a7),
	.cin(gnd),
	.combout(\ram_rom_data_reg[7]~7_combout ),
	.cout());
// synopsys translate_off
defparam \ram_rom_data_reg[7]~7 .lut_mask = 16'hDD88;
defparam \ram_rom_data_reg[7]~7 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X50_Y29_N28
cycloneive_lcell_comb \ram_rom_data_reg[8]~8 (
	.dataa(address_reg_b_0),
	.datab(ram_block3a40),
	.datac(gnd),
	.datad(ram_block3a8),
	.cin(gnd),
	.combout(\ram_rom_data_reg[8]~8_combout ),
	.cout());
// synopsys translate_off
defparam \ram_rom_data_reg[8]~8 .lut_mask = 16'hDD88;
defparam \ram_rom_data_reg[8]~8 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X48_Y35_N12
cycloneive_lcell_comb \ram_rom_data_reg[9]~9 (
	.dataa(address_reg_b_0),
	.datab(ram_block3a41),
	.datac(gnd),
	.datad(ram_block3a9),
	.cin(gnd),
	.combout(\ram_rom_data_reg[9]~9_combout ),
	.cout());
// synopsys translate_off
defparam \ram_rom_data_reg[9]~9 .lut_mask = 16'hDD88;
defparam \ram_rom_data_reg[9]~9 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X48_Y35_N30
cycloneive_lcell_comb \ram_rom_data_reg[10]~10 (
	.dataa(address_reg_b_0),
	.datab(ram_block3a10),
	.datac(gnd),
	.datad(ram_block3a42),
	.cin(gnd),
	.combout(\ram_rom_data_reg[10]~10_combout ),
	.cout());
// synopsys translate_off
defparam \ram_rom_data_reg[10]~10 .lut_mask = 16'hEE44;
defparam \ram_rom_data_reg[10]~10 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X48_Y35_N8
cycloneive_lcell_comb \ram_rom_data_reg[11]~11 (
	.dataa(address_reg_b_0),
	.datab(ram_block3a11),
	.datac(gnd),
	.datad(ram_block3a43),
	.cin(gnd),
	.combout(\ram_rom_data_reg[11]~11_combout ),
	.cout());
// synopsys translate_off
defparam \ram_rom_data_reg[11]~11 .lut_mask = 16'hEE44;
defparam \ram_rom_data_reg[11]~11 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X48_Y35_N26
cycloneive_lcell_comb \ram_rom_data_reg[12]~12 (
	.dataa(address_reg_b_0),
	.datab(ram_block3a12),
	.datac(gnd),
	.datad(ram_block3a44),
	.cin(gnd),
	.combout(\ram_rom_data_reg[12]~12_combout ),
	.cout());
// synopsys translate_off
defparam \ram_rom_data_reg[12]~12 .lut_mask = 16'hEE44;
defparam \ram_rom_data_reg[12]~12 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X48_Y35_N16
cycloneive_lcell_comb \ram_rom_data_reg[13]~13 (
	.dataa(address_reg_b_0),
	.datab(ram_block3a13),
	.datac(gnd),
	.datad(ram_block3a45),
	.cin(gnd),
	.combout(\ram_rom_data_reg[13]~13_combout ),
	.cout());
// synopsys translate_off
defparam \ram_rom_data_reg[13]~13 .lut_mask = 16'hEE44;
defparam \ram_rom_data_reg[13]~13 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X48_Y35_N18
cycloneive_lcell_comb \ram_rom_data_reg[14]~14 (
	.dataa(address_reg_b_0),
	.datab(ram_block3a46),
	.datac(gnd),
	.datad(ram_block3a14),
	.cin(gnd),
	.combout(\ram_rom_data_reg[14]~14_combout ),
	.cout());
// synopsys translate_off
defparam \ram_rom_data_reg[14]~14 .lut_mask = 16'hDD88;
defparam \ram_rom_data_reg[14]~14 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X48_Y35_N28
cycloneive_lcell_comb \ram_rom_data_reg[15]~15 (
	.dataa(address_reg_b_0),
	.datab(ram_block3a47),
	.datac(gnd),
	.datad(ram_block3a15),
	.cin(gnd),
	.combout(\ram_rom_data_reg[15]~15_combout ),
	.cout());
// synopsys translate_off
defparam \ram_rom_data_reg[15]~15 .lut_mask = 16'hDD88;
defparam \ram_rom_data_reg[15]~15 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X48_Y35_N14
cycloneive_lcell_comb \ram_rom_data_reg[16]~16 (
	.dataa(address_reg_b_0),
	.datab(ram_block3a48),
	.datac(gnd),
	.datad(ram_block3a16),
	.cin(gnd),
	.combout(\ram_rom_data_reg[16]~16_combout ),
	.cout());
// synopsys translate_off
defparam \ram_rom_data_reg[16]~16 .lut_mask = 16'hDD88;
defparam \ram_rom_data_reg[16]~16 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X48_Y35_N20
cycloneive_lcell_comb \ram_rom_data_reg[17]~17 (
	.dataa(address_reg_b_0),
	.datab(ram_block3a49),
	.datac(gnd),
	.datad(ram_block3a17),
	.cin(gnd),
	.combout(\ram_rom_data_reg[17]~17_combout ),
	.cout());
// synopsys translate_off
defparam \ram_rom_data_reg[17]~17 .lut_mask = 16'hDD88;
defparam \ram_rom_data_reg[17]~17 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X63_Y29_N24
cycloneive_lcell_comb \ram_rom_data_reg[18]~18 (
	.dataa(address_reg_b_0),
	.datab(ram_block3a50),
	.datac(gnd),
	.datad(ram_block3a18),
	.cin(gnd),
	.combout(\ram_rom_data_reg[18]~18_combout ),
	.cout());
// synopsys translate_off
defparam \ram_rom_data_reg[18]~18 .lut_mask = 16'hDD88;
defparam \ram_rom_data_reg[18]~18 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X63_Y29_N30
cycloneive_lcell_comb \ram_rom_data_reg[19]~19 (
	.dataa(ram_block3a19),
	.datab(ram_block3a51),
	.datac(gnd),
	.datad(address_reg_b_0),
	.cin(gnd),
	.combout(\ram_rom_data_reg[19]~19_combout ),
	.cout());
// synopsys translate_off
defparam \ram_rom_data_reg[19]~19 .lut_mask = 16'hCCAA;
defparam \ram_rom_data_reg[19]~19 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X74_Y31_N28
cycloneive_lcell_comb \ram_rom_data_reg[20]~20 (
	.dataa(ram_block3a20),
	.datab(address_reg_b_0),
	.datac(gnd),
	.datad(ram_block3a52),
	.cin(gnd),
	.combout(\ram_rom_data_reg[20]~20_combout ),
	.cout());
// synopsys translate_off
defparam \ram_rom_data_reg[20]~20 .lut_mask = 16'hEE22;
defparam \ram_rom_data_reg[20]~20 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X74_Y31_N26
cycloneive_lcell_comb \ram_rom_data_reg[21]~21 (
	.dataa(ram_block3a53),
	.datab(address_reg_b_0),
	.datac(gnd),
	.datad(ram_block3a21),
	.cin(gnd),
	.combout(\ram_rom_data_reg[21]~21_combout ),
	.cout());
// synopsys translate_off
defparam \ram_rom_data_reg[21]~21 .lut_mask = 16'hBB88;
defparam \ram_rom_data_reg[21]~21 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X74_Y31_N24
cycloneive_lcell_comb \ram_rom_data_reg[22]~22 (
	.dataa(address_reg_b_0),
	.datab(ram_block3a22),
	.datac(gnd),
	.datad(ram_block3a54),
	.cin(gnd),
	.combout(\ram_rom_data_reg[22]~22_combout ),
	.cout());
// synopsys translate_off
defparam \ram_rom_data_reg[22]~22 .lut_mask = 16'hEE44;
defparam \ram_rom_data_reg[22]~22 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X74_Y31_N14
cycloneive_lcell_comb \ram_rom_data_reg[23]~23 (
	.dataa(ram_block3a55),
	.datab(address_reg_b_0),
	.datac(gnd),
	.datad(ram_block3a23),
	.cin(gnd),
	.combout(\ram_rom_data_reg[23]~23_combout ),
	.cout());
// synopsys translate_off
defparam \ram_rom_data_reg[23]~23 .lut_mask = 16'hBB88;
defparam \ram_rom_data_reg[23]~23 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X74_Y31_N0
cycloneive_lcell_comb \ram_rom_data_reg[24]~24 (
	.dataa(address_reg_b_0),
	.datab(ram_block3a56),
	.datac(gnd),
	.datad(ram_block3a24),
	.cin(gnd),
	.combout(\ram_rom_data_reg[24]~24_combout ),
	.cout());
// synopsys translate_off
defparam \ram_rom_data_reg[24]~24 .lut_mask = 16'hDD88;
defparam \ram_rom_data_reg[24]~24 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X74_Y31_N30
cycloneive_lcell_comb \ram_rom_data_reg[25]~25 (
	.dataa(address_reg_b_0),
	.datab(ram_block3a25),
	.datac(gnd),
	.datad(ram_block3a57),
	.cin(gnd),
	.combout(\ram_rom_data_reg[25]~25_combout ),
	.cout());
// synopsys translate_off
defparam \ram_rom_data_reg[25]~25 .lut_mask = 16'hEE44;
defparam \ram_rom_data_reg[25]~25 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X74_Y31_N20
cycloneive_lcell_comb \ram_rom_data_reg[26]~26 (
	.dataa(ram_block3a26),
	.datab(address_reg_b_0),
	.datac(gnd),
	.datad(ram_block3a58),
	.cin(gnd),
	.combout(\ram_rom_data_reg[26]~26_combout ),
	.cout());
// synopsys translate_off
defparam \ram_rom_data_reg[26]~26 .lut_mask = 16'hEE22;
defparam \ram_rom_data_reg[26]~26 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X74_Y31_N10
cycloneive_lcell_comb \ram_rom_data_reg[27]~27 (
	.dataa(ram_block3a59),
	.datab(address_reg_b_0),
	.datac(gnd),
	.datad(ram_block3a27),
	.cin(gnd),
	.combout(\ram_rom_data_reg[27]~27_combout ),
	.cout());
// synopsys translate_off
defparam \ram_rom_data_reg[27]~27 .lut_mask = 16'hBB88;
defparam \ram_rom_data_reg[27]~27 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X74_Y31_N8
cycloneive_lcell_comb \ram_rom_data_reg[28]~28 (
	.dataa(ram_block3a60),
	.datab(ram_block3a28),
	.datac(gnd),
	.datad(address_reg_b_0),
	.cin(gnd),
	.combout(\ram_rom_data_reg[28]~28_combout ),
	.cout());
// synopsys translate_off
defparam \ram_rom_data_reg[28]~28 .lut_mask = 16'hAACC;
defparam \ram_rom_data_reg[28]~28 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X74_Y31_N18
cycloneive_lcell_comb \ram_rom_data_reg[29]~29 (
	.dataa(ram_block3a61),
	.datab(address_reg_b_0),
	.datac(gnd),
	.datad(ram_block3a29),
	.cin(gnd),
	.combout(\ram_rom_data_reg[29]~29_combout ),
	.cout());
// synopsys translate_off
defparam \ram_rom_data_reg[29]~29 .lut_mask = 16'hBB88;
defparam \ram_rom_data_reg[29]~29 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X50_Y29_N26
cycloneive_lcell_comb \ram_rom_data_reg[30]~30 (
	.dataa(address_reg_b_0),
	.datab(ram_block3a30),
	.datac(gnd),
	.datad(ram_block3a62),
	.cin(gnd),
	.combout(\ram_rom_data_reg[30]~30_combout ),
	.cout());
// synopsys translate_off
defparam \ram_rom_data_reg[30]~30 .lut_mask = 16'hEE44;
defparam \ram_rom_data_reg[30]~30 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X50_Y29_N24
cycloneive_lcell_comb \ram_rom_data_reg[31]~31 (
	.dataa(address_reg_b_0),
	.datab(ram_block3a31),
	.datac(gnd),
	.datad(ram_block3a63),
	.cin(gnd),
	.combout(\ram_rom_data_reg[31]~31_combout ),
	.cout());
// synopsys translate_off
defparam \ram_rom_data_reg[31]~31 .lut_mask = 16'hEE44;
defparam \ram_rom_data_reg[31]~31 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X46_Y34_N30
cycloneive_lcell_comb \ir_loaded_address_reg[0]~feeder (
	.dataa(gnd),
	.datab(gnd),
	.datac(ram_rom_addr_reg_0),
	.datad(gnd),
	.cin(gnd),
	.combout(\ir_loaded_address_reg[0]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \ir_loaded_address_reg[0]~feeder .lut_mask = 16'hF0F0;
defparam \ir_loaded_address_reg[0]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X46_Y34_N16
cycloneive_lcell_comb \process_0~0 (
	.dataa(irf_reg_4_1),
	.datab(gnd),
	.datac(ir_in[0]),
	.datad(gnd),
	.cin(gnd),
	.combout(\process_0~0_combout ),
	.cout());
// synopsys translate_off
defparam \process_0~0 .lut_mask = 16'hFAFA;
defparam \process_0~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X46_Y34_N18
cycloneive_lcell_comb \process_0~1 (
	.dataa(node_ena_1),
	.datab(ir_in[3]),
	.datac(virtual_ir_scan_reg),
	.datad(state_5),
	.cin(gnd),
	.combout(\process_0~1_combout ),
	.cout());
// synopsys translate_off
defparam \process_0~1 .lut_mask = 16'h0800;
defparam \process_0~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X46_Y31_N0
cycloneive_lcell_comb \ir_loaded_address_reg[1]~feeder (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(ram_rom_addr_reg_1),
	.cin(gnd),
	.combout(\ir_loaded_address_reg[1]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \ir_loaded_address_reg[1]~feeder .lut_mask = 16'hFF00;
defparam \ir_loaded_address_reg[1]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X46_Y31_N10
cycloneive_lcell_comb \ir_loaded_address_reg[2]~feeder (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(ram_rom_addr_reg_2),
	.cin(gnd),
	.combout(\ir_loaded_address_reg[2]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \ir_loaded_address_reg[2]~feeder .lut_mask = 16'hFF00;
defparam \ir_loaded_address_reg[2]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X46_Y31_N4
cycloneive_lcell_comb \ir_loaded_address_reg[3]~feeder (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(ram_rom_addr_reg_3),
	.cin(gnd),
	.combout(\ir_loaded_address_reg[3]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \ir_loaded_address_reg[3]~feeder .lut_mask = 16'hFF00;
defparam \ir_loaded_address_reg[3]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X46_Y34_N24
cycloneive_lcell_comb \bypass_reg_out~0 (
	.dataa(gnd),
	.datab(altera_internal_jtag),
	.datac(\bypass_reg_out~q ),
	.datad(node_ena_1),
	.cin(gnd),
	.combout(\bypass_reg_out~0_combout ),
	.cout());
// synopsys translate_off
defparam \bypass_reg_out~0 .lut_mask = 16'hCCF0;
defparam \bypass_reg_out~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X46_Y34_N25
dffeas bypass_reg_out(
	.clk(raw_tck),
	.d(\bypass_reg_out~0_combout ),
	.asdata(vcc),
	.clrn(!clr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\bypass_reg_out~q ),
	.prn(vcc));
// synopsys translate_off
defparam bypass_reg_out.is_wysiwyg = "true";
defparam bypass_reg_out.power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X46_Y34_N2
cycloneive_lcell_comb \tdo~0 (
	.dataa(ram_rom_data_reg_0),
	.datab(irf_reg_2_1),
	.datac(irf_reg_1_1),
	.datad(\bypass_reg_out~q ),
	.cin(gnd),
	.combout(\tdo~0_combout ),
	.cout());
// synopsys translate_off
defparam \tdo~0 .lut_mask = 16'hABA8;
defparam \tdo~0 .sum_lutc_input = "datac";
// synopsys translate_on

endmodule

module sld_rom_sr (
	WORD_SR_0,
	sdr,
	altera_internal_jtag,
	state_4,
	virtual_ir_scan_reg,
	state_3,
	state_8,
	TCK,
	devpor,
	devclrn,
	devoe);
output 	WORD_SR_0;
input 	sdr;
input 	altera_internal_jtag;
input 	state_4;
input 	virtual_ir_scan_reg;
input 	state_3;
input 	state_8;
input 	TCK;

// Design Ports Information

input 	devpor;
input 	devclrn;
input 	devoe;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
assign unknown = 1'bx;

wire \WORD_SR~3_combout ;
wire \WORD_SR~7_combout ;
wire \WORD_SR~8_combout ;
wire \word_counter[4]~13_combout ;
wire \WORD_SR~10_combout ;
wire \WORD_SR~11_combout ;
wire \clear_signal~combout ;
wire \word_counter[0]~7_combout ;
wire \word_counter[4]~19_combout ;
wire \word_counter[4]~14_combout ;
wire \word_counter[0]~8 ;
wire \word_counter[1]~10 ;
wire \word_counter[2]~11_combout ;
wire \word_counter[2]~12 ;
wire \word_counter[3]~15_combout ;
wire \word_counter[3]~16 ;
wire \word_counter[4]~17_combout ;
wire \word_counter[1]~9_combout ;
wire \WORD_SR~13_combout ;
wire \WORD_SR~14_combout ;
wire \WORD_SR~15_combout ;
wire \WORD_SR[0]~6_combout ;
wire \WORD_SR~12_combout ;
wire \WORD_SR~9_combout ;
wire \WORD_SR~2_combout ;
wire \WORD_SR~4_combout ;
wire \WORD_SR~5_combout ;
wire [4:0] word_counter;
wire [3:0] WORD_SR;


// Location: LCCOMB_X47_Y32_N22
cycloneive_lcell_comb \WORD_SR~3 (
	.dataa(word_counter[4]),
	.datab(word_counter[0]),
	.datac(word_counter[2]),
	.datad(word_counter[1]),
	.cin(gnd),
	.combout(\WORD_SR~3_combout ),
	.cout());
// synopsys translate_off
defparam \WORD_SR~3 .lut_mask = 16'hBA02;
defparam \WORD_SR~3 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X46_Y32_N24
cycloneive_lcell_comb \WORD_SR~7 (
	.dataa(word_counter[0]),
	.datab(state_4),
	.datac(word_counter[4]),
	.datad(word_counter[1]),
	.cin(gnd),
	.combout(\WORD_SR~7_combout ),
	.cout());
// synopsys translate_off
defparam \WORD_SR~7 .lut_mask = 16'h1101;
defparam \WORD_SR~7 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X46_Y32_N6
cycloneive_lcell_comb \WORD_SR~8 (
	.dataa(gnd),
	.datab(word_counter[2]),
	.datac(word_counter[3]),
	.datad(\WORD_SR~7_combout ),
	.cin(gnd),
	.combout(\WORD_SR~8_combout ),
	.cout());
// synopsys translate_off
defparam \WORD_SR~8 .lut_mask = 16'h0300;
defparam \WORD_SR~8 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X46_Y32_N26
cycloneive_lcell_comb \word_counter[4]~13 (
	.dataa(word_counter[2]),
	.datab(word_counter[4]),
	.datac(word_counter[3]),
	.datad(word_counter[1]),
	.cin(gnd),
	.combout(\word_counter[4]~13_combout ),
	.cout());
// synopsys translate_off
defparam \word_counter[4]~13 .lut_mask = 16'hFFF7;
defparam \word_counter[4]~13 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X47_Y32_N24
cycloneive_lcell_comb \WORD_SR~10 (
	.dataa(word_counter[4]),
	.datab(word_counter[0]),
	.datac(word_counter[2]),
	.datad(word_counter[1]),
	.cin(gnd),
	.combout(\WORD_SR~10_combout ),
	.cout());
// synopsys translate_off
defparam \WORD_SR~10 .lut_mask = 16'hCABA;
defparam \WORD_SR~10 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X47_Y32_N2
cycloneive_lcell_comb \WORD_SR~11 (
	.dataa(gnd),
	.datab(\WORD_SR~10_combout ),
	.datac(word_counter[0]),
	.datad(\WORD_SR~2_combout ),
	.cin(gnd),
	.combout(\WORD_SR~11_combout ),
	.cout());
// synopsys translate_off
defparam \WORD_SR~11 .lut_mask = 16'hC3C0;
defparam \WORD_SR~11 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X46_Y32_N13
dffeas \WORD_SR[0] (
	.clk(TCK),
	.d(\WORD_SR~5_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\WORD_SR[0]~6_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(WORD_SR_0),
	.prn(vcc));
// synopsys translate_off
defparam \WORD_SR[0] .is_wysiwyg = "true";
defparam \WORD_SR[0] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X46_Y32_N28
cycloneive_lcell_comb clear_signal(
	.dataa(state_8),
	.datab(gnd),
	.datac(virtual_ir_scan_reg),
	.datad(gnd),
	.cin(gnd),
	.combout(\clear_signal~combout ),
	.cout());
// synopsys translate_off
defparam clear_signal.lut_mask = 16'hA0A0;
defparam clear_signal.sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X47_Y32_N4
cycloneive_lcell_comb \word_counter[0]~7 (
	.dataa(gnd),
	.datab(word_counter[0]),
	.datac(gnd),
	.datad(vcc),
	.cin(gnd),
	.combout(\word_counter[0]~7_combout ),
	.cout(\word_counter[0]~8 ));
// synopsys translate_off
defparam \word_counter[0]~7 .lut_mask = 16'h33CC;
defparam \word_counter[0]~7 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X46_Y32_N16
cycloneive_lcell_comb \word_counter[4]~19 (
	.dataa(\word_counter[4]~13_combout ),
	.datab(virtual_ir_scan_reg),
	.datac(state_8),
	.datad(word_counter[0]),
	.cin(gnd),
	.combout(\word_counter[4]~19_combout ),
	.cout());
// synopsys translate_off
defparam \word_counter[4]~19 .lut_mask = 16'hC0D5;
defparam \word_counter[4]~19 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X46_Y32_N0
cycloneive_lcell_comb \word_counter[4]~14 (
	.dataa(sdr),
	.datab(\clear_signal~combout ),
	.datac(state_3),
	.datad(state_4),
	.cin(gnd),
	.combout(\word_counter[4]~14_combout ),
	.cout());
// synopsys translate_off
defparam \word_counter[4]~14 .lut_mask = 16'hCCEC;
defparam \word_counter[4]~14 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X47_Y32_N5
dffeas \word_counter[0] (
	.clk(TCK),
	.d(\word_counter[0]~7_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\word_counter[4]~19_combout ),
	.sload(gnd),
	.ena(\word_counter[4]~14_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(word_counter[0]),
	.prn(vcc));
// synopsys translate_off
defparam \word_counter[0] .is_wysiwyg = "true";
defparam \word_counter[0] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X47_Y32_N6
cycloneive_lcell_comb \word_counter[1]~9 (
	.dataa(word_counter[1]),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\word_counter[0]~8 ),
	.combout(\word_counter[1]~9_combout ),
	.cout(\word_counter[1]~10 ));
// synopsys translate_off
defparam \word_counter[1]~9 .lut_mask = 16'h5A5F;
defparam \word_counter[1]~9 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X47_Y32_N8
cycloneive_lcell_comb \word_counter[2]~11 (
	.dataa(gnd),
	.datab(word_counter[2]),
	.datac(gnd),
	.datad(vcc),
	.cin(\word_counter[1]~10 ),
	.combout(\word_counter[2]~11_combout ),
	.cout(\word_counter[2]~12 ));
// synopsys translate_off
defparam \word_counter[2]~11 .lut_mask = 16'hC30C;
defparam \word_counter[2]~11 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: FF_X47_Y32_N9
dffeas \word_counter[2] (
	.clk(TCK),
	.d(\word_counter[2]~11_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\word_counter[4]~19_combout ),
	.sload(gnd),
	.ena(\word_counter[4]~14_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(word_counter[2]),
	.prn(vcc));
// synopsys translate_off
defparam \word_counter[2] .is_wysiwyg = "true";
defparam \word_counter[2] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X47_Y32_N10
cycloneive_lcell_comb \word_counter[3]~15 (
	.dataa(gnd),
	.datab(word_counter[3]),
	.datac(gnd),
	.datad(vcc),
	.cin(\word_counter[2]~12 ),
	.combout(\word_counter[3]~15_combout ),
	.cout(\word_counter[3]~16 ));
// synopsys translate_off
defparam \word_counter[3]~15 .lut_mask = 16'h3C3F;
defparam \word_counter[3]~15 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: FF_X47_Y32_N11
dffeas \word_counter[3] (
	.clk(TCK),
	.d(\word_counter[3]~15_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\word_counter[4]~19_combout ),
	.sload(gnd),
	.ena(\word_counter[4]~14_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(word_counter[3]),
	.prn(vcc));
// synopsys translate_off
defparam \word_counter[3] .is_wysiwyg = "true";
defparam \word_counter[3] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X47_Y32_N12
cycloneive_lcell_comb \word_counter[4]~17 (
	.dataa(word_counter[4]),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.cin(\word_counter[3]~16 ),
	.combout(\word_counter[4]~17_combout ),
	.cout());
// synopsys translate_off
defparam \word_counter[4]~17 .lut_mask = 16'hA5A5;
defparam \word_counter[4]~17 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: FF_X47_Y32_N13
dffeas \word_counter[4] (
	.clk(TCK),
	.d(\word_counter[4]~17_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\word_counter[4]~19_combout ),
	.sload(gnd),
	.ena(\word_counter[4]~14_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(word_counter[4]),
	.prn(vcc));
// synopsys translate_off
defparam \word_counter[4] .is_wysiwyg = "true";
defparam \word_counter[4] .power_up = "low";
// synopsys translate_on

// Location: FF_X47_Y32_N7
dffeas \word_counter[1] (
	.clk(TCK),
	.d(\word_counter[1]~9_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\word_counter[4]~19_combout ),
	.sload(gnd),
	.ena(\word_counter[4]~14_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(word_counter[1]),
	.prn(vcc));
// synopsys translate_off
defparam \word_counter[1] .is_wysiwyg = "true";
defparam \word_counter[1] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X46_Y32_N20
cycloneive_lcell_comb \WORD_SR~13 (
	.dataa(word_counter[2]),
	.datab(word_counter[4]),
	.datac(word_counter[3]),
	.datad(word_counter[1]),
	.cin(gnd),
	.combout(\WORD_SR~13_combout ),
	.cout());
// synopsys translate_off
defparam \WORD_SR~13 .lut_mask = 16'h2000;
defparam \WORD_SR~13 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X46_Y32_N18
cycloneive_lcell_comb \WORD_SR~14 (
	.dataa(word_counter[0]),
	.datab(state_4),
	.datac(altera_internal_jtag),
	.datad(\WORD_SR~13_combout ),
	.cin(gnd),
	.combout(\WORD_SR~14_combout ),
	.cout());
// synopsys translate_off
defparam \WORD_SR~14 .lut_mask = 16'hD1C0;
defparam \WORD_SR~14 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X46_Y32_N30
cycloneive_lcell_comb \WORD_SR~15 (
	.dataa(state_8),
	.datab(gnd),
	.datac(virtual_ir_scan_reg),
	.datad(\WORD_SR~14_combout ),
	.cin(gnd),
	.combout(\WORD_SR~15_combout ),
	.cout());
// synopsys translate_off
defparam \WORD_SR~15 .lut_mask = 16'h5F00;
defparam \WORD_SR~15 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X46_Y32_N22
cycloneive_lcell_comb \WORD_SR[0]~6 (
	.dataa(sdr),
	.datab(\clear_signal~combout ),
	.datac(state_3),
	.datad(state_4),
	.cin(gnd),
	.combout(\WORD_SR[0]~6_combout ),
	.cout());
// synopsys translate_off
defparam \WORD_SR[0]~6 .lut_mask = 16'hEEEC;
defparam \WORD_SR[0]~6 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X46_Y32_N31
dffeas \WORD_SR[3] (
	.clk(TCK),
	.d(\WORD_SR~15_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\WORD_SR[0]~6_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(WORD_SR[3]),
	.prn(vcc));
// synopsys translate_off
defparam \WORD_SR[3] .is_wysiwyg = "true";
defparam \WORD_SR[3] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X46_Y32_N8
cycloneive_lcell_comb \WORD_SR~12 (
	.dataa(\WORD_SR~11_combout ),
	.datab(\clear_signal~combout ),
	.datac(WORD_SR[3]),
	.datad(state_4),
	.cin(gnd),
	.combout(\WORD_SR~12_combout ),
	.cout());
// synopsys translate_off
defparam \WORD_SR~12 .lut_mask = 16'h3022;
defparam \WORD_SR~12 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X46_Y32_N9
dffeas \WORD_SR[2] (
	.clk(TCK),
	.d(\WORD_SR~12_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\WORD_SR[0]~6_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(WORD_SR[2]),
	.prn(vcc));
// synopsys translate_off
defparam \WORD_SR[2] .is_wysiwyg = "true";
defparam \WORD_SR[2] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X46_Y32_N10
cycloneive_lcell_comb \WORD_SR~9 (
	.dataa(\WORD_SR~8_combout ),
	.datab(\clear_signal~combout ),
	.datac(WORD_SR[2]),
	.datad(state_4),
	.cin(gnd),
	.combout(\WORD_SR~9_combout ),
	.cout());
// synopsys translate_off
defparam \WORD_SR~9 .lut_mask = 16'h3222;
defparam \WORD_SR~9 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X46_Y32_N11
dffeas \WORD_SR[1] (
	.clk(TCK),
	.d(\WORD_SR~9_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\WORD_SR[0]~6_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(WORD_SR[1]),
	.prn(vcc));
// synopsys translate_off
defparam \WORD_SR[1] .is_wysiwyg = "true";
defparam \WORD_SR[1] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X47_Y32_N0
cycloneive_lcell_comb \WORD_SR~2 (
	.dataa(word_counter[4]),
	.datab(word_counter[3]),
	.datac(word_counter[2]),
	.datad(word_counter[1]),
	.cin(gnd),
	.combout(\WORD_SR~2_combout ),
	.cout());
// synopsys translate_off
defparam \WORD_SR~2 .lut_mask = 16'h4043;
defparam \WORD_SR~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X47_Y32_N30
cycloneive_lcell_comb \WORD_SR~4 (
	.dataa(\WORD_SR~3_combout ),
	.datab(gnd),
	.datac(word_counter[0]),
	.datad(\WORD_SR~2_combout ),
	.cin(gnd),
	.combout(\WORD_SR~4_combout ),
	.cout());
// synopsys translate_off
defparam \WORD_SR~4 .lut_mask = 16'hAAA0;
defparam \WORD_SR~4 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X46_Y32_N12
cycloneive_lcell_comb \WORD_SR~5 (
	.dataa(WORD_SR[1]),
	.datab(\clear_signal~combout ),
	.datac(\WORD_SR~4_combout ),
	.datad(state_4),
	.cin(gnd),
	.combout(\WORD_SR~5_combout ),
	.cout());
// synopsys translate_off
defparam \WORD_SR~5 .lut_mask = 16'h2230;
defparam \WORD_SR~5 .sum_lutc_input = "datac";
// synopsys translate_on

endmodule
